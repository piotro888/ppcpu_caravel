magic
tech sky130A
magscale 1 2
timestamp 1672497455
<< metal1 >>
rect 246390 700952 246396 701004
rect 246448 700992 246454 701004
rect 332502 700992 332508 701004
rect 246448 700964 332508 700992
rect 246448 700952 246454 700964
rect 332502 700952 332508 700964
rect 332560 700952 332566 701004
rect 246482 700884 246488 700936
rect 246540 700924 246546 700936
rect 348786 700924 348792 700936
rect 246540 700896 348792 700924
rect 246540 700884 246546 700896
rect 348786 700884 348792 700896
rect 348844 700884 348850 700936
rect 243630 700816 243636 700868
rect 243688 700856 243694 700868
rect 364978 700856 364984 700868
rect 243688 700828 364984 700856
rect 243688 700816 243694 700828
rect 364978 700816 364984 700828
rect 365036 700816 365042 700868
rect 240778 700748 240784 700800
rect 240836 700788 240842 700800
rect 397454 700788 397460 700800
rect 240836 700760 397460 700788
rect 240836 700748 240842 700760
rect 397454 700748 397460 700760
rect 397512 700748 397518 700800
rect 253290 700680 253296 700732
rect 253348 700720 253354 700732
rect 429838 700720 429844 700732
rect 253348 700692 429844 700720
rect 253348 700680 253354 700692
rect 429838 700680 429844 700692
rect 429896 700680 429902 700732
rect 218698 700612 218704 700664
rect 218756 700652 218762 700664
rect 413646 700652 413652 700664
rect 218756 700624 413652 700652
rect 218756 700612 218762 700624
rect 413646 700612 413652 700624
rect 413704 700612 413710 700664
rect 105446 700544 105452 700596
rect 105504 700584 105510 700596
rect 142798 700584 142804 700596
rect 105504 700556 142804 700584
rect 105504 700544 105510 700556
rect 142798 700544 142804 700556
rect 142856 700544 142862 700596
rect 249058 700544 249064 700596
rect 249116 700584 249122 700596
rect 462314 700584 462320 700596
rect 249116 700556 462320 700584
rect 249116 700544 249122 700556
rect 462314 700544 462320 700556
rect 462372 700544 462378 700596
rect 89162 700476 89168 700528
rect 89220 700516 89226 700528
rect 151078 700516 151084 700528
rect 89220 700488 151084 700516
rect 89220 700476 89226 700488
rect 151078 700476 151084 700488
rect 151136 700476 151142 700528
rect 233878 700476 233884 700528
rect 233936 700516 233942 700528
rect 478506 700516 478512 700528
rect 233936 700488 478512 700516
rect 233936 700476 233942 700488
rect 478506 700476 478512 700488
rect 478564 700476 478570 700528
rect 72970 700408 72976 700460
rect 73028 700448 73034 700460
rect 148318 700448 148324 700460
rect 73028 700420 148324 700448
rect 73028 700408 73034 700420
rect 148318 700408 148324 700420
rect 148376 700408 148382 700460
rect 243538 700408 243544 700460
rect 243596 700448 243602 700460
rect 494790 700448 494796 700460
rect 243596 700420 494796 700448
rect 243596 700408 243602 700420
rect 494790 700408 494796 700420
rect 494848 700408 494854 700460
rect 24302 700340 24308 700392
rect 24360 700380 24366 700392
rect 138658 700380 138664 700392
rect 24360 700352 138664 700380
rect 24360 700340 24366 700352
rect 138658 700340 138664 700352
rect 138716 700340 138722 700392
rect 240962 700340 240968 700392
rect 241020 700380 241026 700392
rect 527174 700380 527180 700392
rect 241020 700352 527180 700380
rect 241020 700340 241026 700352
rect 527174 700340 527180 700352
rect 527232 700340 527238 700392
rect 40494 700272 40500 700324
rect 40552 700312 40558 700324
rect 157978 700312 157984 700324
rect 40552 700284 157984 700312
rect 40552 700272 40558 700284
rect 157978 700272 157984 700284
rect 158036 700272 158042 700324
rect 202782 700272 202788 700324
rect 202840 700312 202846 700324
rect 218146 700312 218152 700324
rect 202840 700284 218152 700312
rect 202840 700272 202846 700284
rect 218146 700272 218152 700284
rect 218204 700272 218210 700324
rect 232498 700272 232504 700324
rect 232556 700312 232562 700324
rect 543458 700312 543464 700324
rect 232556 700284 543464 700312
rect 232556 700272 232562 700284
rect 543458 700272 543464 700284
rect 543516 700272 543522 700324
rect 253198 700204 253204 700256
rect 253256 700244 253262 700256
rect 300118 700244 300124 700256
rect 253256 700216 300124 700244
rect 253256 700204 253262 700216
rect 300118 700204 300124 700216
rect 300176 700204 300182 700256
rect 251818 700136 251824 700188
rect 251876 700176 251882 700188
rect 283834 700176 283840 700188
rect 251876 700148 283840 700176
rect 251876 700136 251882 700148
rect 283834 700136 283840 700148
rect 283892 700136 283898 700188
rect 238018 700068 238024 700120
rect 238076 700108 238082 700120
rect 267642 700108 267648 700120
rect 238076 700080 267648 700108
rect 238076 700068 238082 700080
rect 267642 700068 267648 700080
rect 267700 700068 267706 700120
rect 239398 696940 239404 696992
rect 239456 696980 239462 696992
rect 580166 696980 580172 696992
rect 239456 696952 580172 696980
rect 239456 696940 239462 696952
rect 580166 696940 580172 696952
rect 580224 696940 580230 696992
rect 3418 683136 3424 683188
rect 3476 683176 3482 683188
rect 158070 683176 158076 683188
rect 3476 683148 158076 683176
rect 3476 683136 3482 683148
rect 158070 683136 158076 683148
rect 158128 683136 158134 683188
rect 221458 683136 221464 683188
rect 221516 683176 221522 683188
rect 580166 683176 580172 683188
rect 221516 683148 580172 683176
rect 221516 683136 221522 683148
rect 580166 683136 580172 683148
rect 580224 683136 580230 683188
rect 3510 670692 3516 670744
rect 3568 670732 3574 670744
rect 141418 670732 141424 670744
rect 3568 670704 141424 670732
rect 3568 670692 3574 670704
rect 141418 670692 141424 670704
rect 141476 670692 141482 670744
rect 3418 656888 3424 656940
rect 3476 656928 3482 656940
rect 144178 656928 144184 656940
rect 3476 656900 144184 656928
rect 3476 656888 3482 656900
rect 144178 656888 144184 656900
rect 144236 656888 144242 656940
rect 234154 644512 234160 644564
rect 234212 644552 234218 644564
rect 251266 644552 251272 644564
rect 234212 644524 251272 644552
rect 234212 644512 234218 644524
rect 251266 644512 251272 644524
rect 251324 644512 251330 644564
rect 233970 644444 233976 644496
rect 234028 644484 234034 644496
rect 251174 644484 251180 644496
rect 234028 644456 251180 644484
rect 234028 644444 234034 644456
rect 251174 644444 251180 644456
rect 251232 644444 251238 644496
rect 234246 643084 234252 643136
rect 234304 643124 234310 643136
rect 251174 643124 251180 643136
rect 234304 643096 251180 643124
rect 234304 643084 234310 643096
rect 251174 643084 251180 643096
rect 251232 643084 251238 643136
rect 231118 641724 231124 641776
rect 231176 641764 231182 641776
rect 251174 641764 251180 641776
rect 231176 641736 251180 641764
rect 231176 641724 231182 641736
rect 251174 641724 251180 641736
rect 251232 641724 251238 641776
rect 239490 640296 239496 640348
rect 239548 640336 239554 640348
rect 251174 640336 251180 640348
rect 239548 640308 251180 640336
rect 239548 640296 239554 640308
rect 251174 640296 251180 640308
rect 251232 640296 251238 640348
rect 224218 638936 224224 638988
rect 224276 638976 224282 638988
rect 251174 638976 251180 638988
rect 224276 638948 251180 638976
rect 224276 638936 224282 638948
rect 251174 638936 251180 638948
rect 251232 638936 251238 638988
rect 228358 637576 228364 637628
rect 228416 637616 228422 637628
rect 251174 637616 251180 637628
rect 228416 637588 251180 637616
rect 228416 637576 228422 637588
rect 251174 637576 251180 637588
rect 251232 637576 251238 637628
rect 244918 634788 244924 634840
rect 244976 634828 244982 634840
rect 251174 634828 251180 634840
rect 244976 634800 251180 634828
rect 244976 634788 244982 634800
rect 251174 634788 251180 634800
rect 251232 634788 251238 634840
rect 225598 633428 225604 633480
rect 225656 633468 225662 633480
rect 251266 633468 251272 633480
rect 225656 633440 251272 633468
rect 225656 633428 225662 633440
rect 251266 633428 251272 633440
rect 251324 633428 251330 633480
rect 228450 632680 228456 632732
rect 228508 632720 228514 632732
rect 251174 632720 251180 632732
rect 228508 632692 251180 632720
rect 228508 632680 228514 632692
rect 251174 632680 251180 632692
rect 251232 632680 251238 632732
rect 3418 632068 3424 632120
rect 3476 632108 3482 632120
rect 158162 632108 158168 632120
rect 3476 632080 158168 632108
rect 3476 632068 3482 632080
rect 158162 632068 158168 632080
rect 158220 632068 158226 632120
rect 220078 632068 220084 632120
rect 220136 632108 220142 632120
rect 251174 632108 251180 632120
rect 220136 632080 251180 632108
rect 220136 632068 220142 632080
rect 251174 632068 251180 632080
rect 251232 632068 251238 632120
rect 232590 630640 232596 630692
rect 232648 630680 232654 630692
rect 251174 630680 251180 630692
rect 232648 630652 251180 630680
rect 232648 630640 232654 630652
rect 251174 630640 251180 630652
rect 251232 630640 251238 630692
rect 222838 629280 222844 629332
rect 222896 629320 222902 629332
rect 251174 629320 251180 629332
rect 222896 629292 251180 629320
rect 222896 629280 222902 629292
rect 251174 629280 251180 629292
rect 251232 629280 251238 629332
rect 231210 627920 231216 627972
rect 231268 627960 231274 627972
rect 251174 627960 251180 627972
rect 231268 627932 251180 627960
rect 231268 627920 231274 627932
rect 251174 627920 251180 627932
rect 251232 627920 251238 627972
rect 231302 626560 231308 626612
rect 231360 626600 231366 626612
rect 251174 626600 251180 626612
rect 231360 626572 251180 626600
rect 231360 626560 231366 626572
rect 251174 626560 251180 626572
rect 251232 626560 251238 626612
rect 245010 625132 245016 625184
rect 245068 625172 245074 625184
rect 251174 625172 251180 625184
rect 245068 625144 251180 625172
rect 245068 625132 245074 625144
rect 251174 625132 251180 625144
rect 251232 625132 251238 625184
rect 236638 623840 236644 623892
rect 236696 623880 236702 623892
rect 251266 623880 251272 623892
rect 236696 623852 251272 623880
rect 236696 623840 236702 623852
rect 251266 623840 251272 623852
rect 251324 623840 251330 623892
rect 228542 623772 228548 623824
rect 228600 623812 228606 623824
rect 251174 623812 251180 623824
rect 228600 623784 251180 623812
rect 228600 623772 228606 623784
rect 251174 623772 251180 623784
rect 251232 623772 251238 623824
rect 222930 622412 222936 622464
rect 222988 622452 222994 622464
rect 251174 622452 251180 622464
rect 222988 622424 251180 622452
rect 222988 622412 222994 622424
rect 251174 622412 251180 622424
rect 251232 622412 251238 622464
rect 242158 620984 242164 621036
rect 242216 621024 242222 621036
rect 251174 621024 251180 621036
rect 242216 620996 251180 621024
rect 242216 620984 242222 620996
rect 251174 620984 251180 620996
rect 251232 620984 251238 621036
rect 226978 619624 226984 619676
rect 227036 619664 227042 619676
rect 251174 619664 251180 619676
rect 227036 619636 251180 619664
rect 227036 619624 227042 619636
rect 251174 619624 251180 619636
rect 251232 619624 251238 619676
rect 3142 618264 3148 618316
rect 3200 618304 3206 618316
rect 146938 618304 146944 618316
rect 3200 618276 146944 618304
rect 3200 618264 3206 618276
rect 146938 618264 146944 618276
rect 146996 618264 147002 618316
rect 224310 618264 224316 618316
rect 224368 618304 224374 618316
rect 251174 618304 251180 618316
rect 224368 618276 251180 618304
rect 224368 618264 224374 618276
rect 251174 618264 251180 618276
rect 251232 618264 251238 618316
rect 221642 616836 221648 616888
rect 221700 616876 221706 616888
rect 251174 616876 251180 616888
rect 221700 616848 251180 616876
rect 221700 616836 221706 616848
rect 251174 616836 251180 616848
rect 251232 616836 251238 616888
rect 574738 616836 574744 616888
rect 574796 616876 574802 616888
rect 580166 616876 580172 616888
rect 574796 616848 580172 616876
rect 574796 616836 574802 616848
rect 580166 616836 580172 616848
rect 580224 616836 580230 616888
rect 239582 615476 239588 615528
rect 239640 615516 239646 615528
rect 251174 615516 251180 615528
rect 239640 615488 251180 615516
rect 239640 615476 239646 615488
rect 251174 615476 251180 615488
rect 251232 615476 251238 615528
rect 235258 614116 235264 614168
rect 235316 614156 235322 614168
rect 251174 614156 251180 614168
rect 235316 614128 251180 614156
rect 235316 614116 235322 614128
rect 251174 614116 251180 614128
rect 251232 614116 251238 614168
rect 246574 612824 246580 612876
rect 246632 612864 246638 612876
rect 251266 612864 251272 612876
rect 246632 612836 251272 612864
rect 246632 612824 246638 612836
rect 251266 612824 251272 612836
rect 251324 612824 251330 612876
rect 221734 612756 221740 612808
rect 221792 612796 221798 612808
rect 251174 612796 251180 612808
rect 221792 612768 251180 612796
rect 221792 612756 221798 612768
rect 251174 612756 251180 612768
rect 251232 612756 251238 612808
rect 238110 611328 238116 611380
rect 238168 611368 238174 611380
rect 251174 611368 251180 611380
rect 238168 611340 251180 611368
rect 238168 611328 238174 611340
rect 251174 611328 251180 611340
rect 251232 611328 251238 611380
rect 229738 609968 229744 610020
rect 229796 610008 229802 610020
rect 251174 610008 251180 610020
rect 229796 609980 251180 610008
rect 229796 609968 229802 609980
rect 251174 609968 251180 609980
rect 251232 609968 251238 610020
rect 229830 608608 229836 608660
rect 229888 608648 229894 608660
rect 251174 608648 251180 608660
rect 229888 608620 251180 608648
rect 229888 608608 229894 608620
rect 251174 608608 251180 608620
rect 251232 608608 251238 608660
rect 221826 607180 221832 607232
rect 221884 607220 221890 607232
rect 251174 607220 251180 607232
rect 221884 607192 251180 607220
rect 221884 607180 221890 607192
rect 251174 607180 251180 607192
rect 251232 607180 251238 607232
rect 3234 605820 3240 605872
rect 3292 605860 3298 605872
rect 135898 605860 135904 605872
rect 3292 605832 135904 605860
rect 3292 605820 3298 605832
rect 135898 605820 135904 605832
rect 135956 605820 135962 605872
rect 238202 604460 238208 604512
rect 238260 604500 238266 604512
rect 251174 604500 251180 604512
rect 238260 604472 251180 604500
rect 238260 604460 238266 604472
rect 251174 604460 251180 604472
rect 251232 604460 251238 604512
rect 227070 603100 227076 603152
rect 227128 603140 227134 603152
rect 251174 603140 251180 603152
rect 227128 603112 251180 603140
rect 227128 603100 227134 603112
rect 251174 603100 251180 603112
rect 251232 603100 251238 603152
rect 249150 601672 249156 601724
rect 249208 601712 249214 601724
rect 251266 601712 251272 601724
rect 249208 601684 251272 601712
rect 249208 601672 249214 601684
rect 251266 601672 251272 601684
rect 251324 601672 251330 601724
rect 235350 600312 235356 600364
rect 235408 600352 235414 600364
rect 251174 600352 251180 600364
rect 235408 600324 251180 600352
rect 235408 600312 235414 600324
rect 251174 600312 251180 600324
rect 251232 600312 251238 600364
rect 232682 598952 232688 599004
rect 232740 598992 232746 599004
rect 251174 598992 251180 599004
rect 232740 598964 251180 598992
rect 232740 598952 232746 598964
rect 251174 598952 251180 598964
rect 251232 598952 251238 599004
rect 247770 597524 247776 597576
rect 247828 597564 247834 597576
rect 251174 597564 251180 597576
rect 247828 597536 251180 597564
rect 247828 597524 247834 597536
rect 251174 597524 251180 597536
rect 251232 597524 251238 597576
rect 247862 594804 247868 594856
rect 247920 594844 247926 594856
rect 251174 594844 251180 594856
rect 247920 594816 251180 594844
rect 247920 594804 247926 594816
rect 251174 594804 251180 594816
rect 251232 594804 251238 594856
rect 223022 593376 223028 593428
rect 223080 593416 223086 593428
rect 251174 593416 251180 593428
rect 223080 593388 251180 593416
rect 223080 593376 223086 593388
rect 251174 593376 251180 593388
rect 251232 593376 251238 593428
rect 243722 592016 243728 592068
rect 243780 592056 243786 592068
rect 251174 592056 251180 592068
rect 243780 592028 251180 592056
rect 243780 592016 243786 592028
rect 251174 592016 251180 592028
rect 251232 592016 251238 592068
rect 111794 590724 111800 590776
rect 111852 590764 111858 590776
rect 119614 590764 119620 590776
rect 111852 590736 119620 590764
rect 111852 590724 111858 590736
rect 119614 590724 119620 590736
rect 119672 590724 119678 590776
rect 246666 590724 246672 590776
rect 246724 590764 246730 590776
rect 251174 590764 251180 590776
rect 246724 590736 251180 590764
rect 246724 590724 246730 590736
rect 251174 590724 251180 590736
rect 251232 590724 251238 590776
rect 111886 590656 111892 590708
rect 111944 590696 111950 590708
rect 140038 590696 140044 590708
rect 111944 590668 140044 590696
rect 111944 590656 111950 590668
rect 140038 590656 140044 590668
rect 140096 590656 140102 590708
rect 220170 590656 220176 590708
rect 220228 590696 220234 590708
rect 251266 590696 251272 590708
rect 220228 590668 251272 590696
rect 220228 590656 220234 590668
rect 251266 590656 251272 590668
rect 251324 590656 251330 590708
rect 111794 589364 111800 589416
rect 111852 589404 111858 589416
rect 123478 589404 123484 589416
rect 111852 589376 123484 589404
rect 111852 589364 111858 589376
rect 123478 589364 123484 589376
rect 123536 589364 123542 589416
rect 111886 589296 111892 589348
rect 111944 589336 111950 589348
rect 142890 589336 142896 589348
rect 111944 589308 142896 589336
rect 111944 589296 111950 589308
rect 142890 589296 142896 589308
rect 142948 589296 142954 589348
rect 241054 589296 241060 589348
rect 241112 589336 241118 589348
rect 251174 589336 251180 589348
rect 241112 589308 251180 589336
rect 241112 589296 241118 589308
rect 251174 589296 251180 589308
rect 251232 589296 251238 589348
rect 111794 587868 111800 587920
rect 111852 587908 111858 587920
rect 123570 587908 123576 587920
rect 111852 587880 123576 587908
rect 111852 587868 111858 587880
rect 123570 587868 123576 587880
rect 123628 587868 123634 587920
rect 229922 587868 229928 587920
rect 229980 587908 229986 587920
rect 251174 587908 251180 587920
rect 229980 587880 251180 587908
rect 229980 587868 229986 587880
rect 251174 587868 251180 587880
rect 251232 587868 251238 587920
rect 111794 586508 111800 586560
rect 111852 586548 111858 586560
rect 123754 586548 123760 586560
rect 111852 586520 123760 586548
rect 111852 586508 111858 586520
rect 123754 586508 123760 586520
rect 123812 586508 123818 586560
rect 112254 585760 112260 585812
rect 112312 585800 112318 585812
rect 123662 585800 123668 585812
rect 112312 585772 123668 585800
rect 112312 585760 112318 585772
rect 123662 585760 123668 585772
rect 123720 585760 123726 585812
rect 111794 585352 111800 585404
rect 111852 585392 111858 585404
rect 113818 585392 113824 585404
rect 111852 585364 113824 585392
rect 111852 585352 111858 585364
rect 113818 585352 113824 585364
rect 113876 585352 113882 585404
rect 245102 585148 245108 585200
rect 245160 585188 245166 585200
rect 251174 585188 251180 585200
rect 245160 585160 251180 585188
rect 245160 585148 245166 585160
rect 251174 585148 251180 585160
rect 251232 585148 251238 585200
rect 111978 584400 111984 584452
rect 112036 584440 112042 584452
rect 120718 584440 120724 584452
rect 112036 584412 120724 584440
rect 112036 584400 112042 584412
rect 120718 584400 120724 584412
rect 120776 584400 120782 584452
rect 111886 583856 111892 583908
rect 111944 583896 111950 583908
rect 113910 583896 113916 583908
rect 111944 583868 113916 583896
rect 111944 583856 111950 583868
rect 113910 583856 113916 583868
rect 113968 583856 113974 583908
rect 111794 583720 111800 583772
rect 111852 583760 111858 583772
rect 117958 583760 117964 583772
rect 111852 583732 117964 583760
rect 111852 583720 111858 583732
rect 117958 583720 117964 583732
rect 118016 583720 118022 583772
rect 232774 583720 232780 583772
rect 232832 583760 232838 583772
rect 251174 583760 251180 583772
rect 232832 583732 251180 583760
rect 232832 583720 232838 583732
rect 251174 583720 251180 583732
rect 251232 583720 251238 583772
rect 111794 582360 111800 582412
rect 111852 582400 111858 582412
rect 115198 582400 115204 582412
rect 111852 582372 115204 582400
rect 111852 582360 111858 582372
rect 115198 582360 115204 582372
rect 115256 582360 115262 582412
rect 230014 582360 230020 582412
rect 230072 582400 230078 582412
rect 251174 582400 251180 582412
rect 230072 582372 251180 582400
rect 230072 582360 230078 582372
rect 251174 582360 251180 582372
rect 251232 582360 251238 582412
rect 111886 581612 111892 581664
rect 111944 581652 111950 581664
rect 138750 581652 138756 581664
rect 111944 581624 138756 581652
rect 111944 581612 111950 581624
rect 138750 581612 138756 581624
rect 138808 581612 138814 581664
rect 111794 581000 111800 581052
rect 111852 581040 111858 581052
rect 122098 581040 122104 581052
rect 111852 581012 122104 581040
rect 111852 581000 111858 581012
rect 122098 581000 122104 581012
rect 122156 581000 122162 581052
rect 220262 581000 220268 581052
rect 220320 581040 220326 581052
rect 251174 581040 251180 581052
rect 220320 581012 251180 581040
rect 220320 581000 220326 581012
rect 251174 581000 251180 581012
rect 251232 581000 251238 581052
rect 111978 580252 111984 580304
rect 112036 580292 112042 580304
rect 122190 580292 122196 580304
rect 112036 580264 122196 580292
rect 112036 580252 112042 580264
rect 122190 580252 122196 580264
rect 122248 580252 122254 580304
rect 111886 579708 111892 579760
rect 111944 579748 111950 579760
rect 116762 579748 116768 579760
rect 111944 579720 116768 579748
rect 111944 579708 111950 579720
rect 116762 579708 116768 579720
rect 116820 579708 116826 579760
rect 249334 579708 249340 579760
rect 249392 579748 249398 579760
rect 251266 579748 251272 579760
rect 249392 579720 251272 579748
rect 249392 579708 249398 579720
rect 251266 579708 251272 579720
rect 251324 579708 251330 579760
rect 3326 579640 3332 579692
rect 3384 579680 3390 579692
rect 29638 579680 29644 579692
rect 3384 579652 29644 579680
rect 3384 579640 3390 579652
rect 29638 579640 29644 579652
rect 29696 579640 29702 579692
rect 111794 579640 111800 579692
rect 111852 579680 111858 579692
rect 134518 579680 134524 579692
rect 111852 579652 134524 579680
rect 111852 579640 111858 579652
rect 134518 579640 134524 579652
rect 134576 579640 134582 579692
rect 242250 579640 242256 579692
rect 242308 579680 242314 579692
rect 251174 579680 251180 579692
rect 242308 579652 251180 579680
rect 242308 579640 242314 579652
rect 251174 579640 251180 579652
rect 251232 579640 251238 579692
rect 111794 578280 111800 578332
rect 111852 578320 111858 578332
rect 130378 578320 130384 578332
rect 111852 578292 130384 578320
rect 111852 578280 111858 578292
rect 130378 578280 130384 578292
rect 130436 578280 130442 578332
rect 111886 578212 111892 578264
rect 111944 578252 111950 578264
rect 133138 578252 133144 578264
rect 111944 578224 133144 578252
rect 111944 578212 111950 578224
rect 133138 578212 133144 578224
rect 133196 578212 133202 578264
rect 227162 578212 227168 578264
rect 227220 578252 227226 578264
rect 251174 578252 251180 578264
rect 227220 578224 251180 578252
rect 227220 578212 227226 578224
rect 251174 578212 251180 578224
rect 251232 578212 251238 578264
rect 249426 576988 249432 577040
rect 249484 577028 249490 577040
rect 251266 577028 251272 577040
rect 249484 577000 251272 577028
rect 249484 576988 249490 577000
rect 251266 576988 251272 577000
rect 251324 576988 251330 577040
rect 111794 576852 111800 576904
rect 111852 576892 111858 576904
rect 152550 576892 152556 576904
rect 111852 576864 152556 576892
rect 111852 576852 111858 576864
rect 152550 576852 152556 576864
rect 152608 576852 152614 576904
rect 111886 575560 111892 575612
rect 111944 575600 111950 575612
rect 132034 575600 132040 575612
rect 111944 575572 132040 575600
rect 111944 575560 111950 575572
rect 132034 575560 132040 575572
rect 132092 575560 132098 575612
rect 111794 575492 111800 575544
rect 111852 575532 111858 575544
rect 141510 575532 141516 575544
rect 111852 575504 141516 575532
rect 111852 575492 111858 575504
rect 141510 575492 141516 575504
rect 141568 575492 141574 575544
rect 239674 575492 239680 575544
rect 239732 575532 239738 575544
rect 251174 575532 251180 575544
rect 239732 575504 251180 575532
rect 239732 575492 239738 575504
rect 251174 575492 251180 575504
rect 251232 575492 251238 575544
rect 111886 574336 111892 574388
rect 111944 574376 111950 574388
rect 114002 574376 114008 574388
rect 111944 574348 114008 574376
rect 111944 574336 111950 574348
rect 114002 574336 114008 574348
rect 114060 574336 114066 574388
rect 111794 574064 111800 574116
rect 111852 574104 111858 574116
rect 152642 574104 152648 574116
rect 111852 574076 152648 574104
rect 111852 574064 111858 574076
rect 152642 574064 152648 574076
rect 152700 574064 152706 574116
rect 231394 574064 231400 574116
rect 231452 574104 231458 574116
rect 251174 574104 251180 574116
rect 231452 574076 251180 574104
rect 231452 574064 231458 574076
rect 251174 574064 251180 574076
rect 251232 574064 251238 574116
rect 111794 572772 111800 572824
rect 111852 572812 111858 572824
rect 134610 572812 134616 572824
rect 111852 572784 134616 572812
rect 111852 572772 111858 572784
rect 134610 572772 134616 572784
rect 134668 572772 134674 572824
rect 111886 572704 111892 572756
rect 111944 572744 111950 572756
rect 142982 572744 142988 572756
rect 111944 572716 142988 572744
rect 111944 572704 111950 572716
rect 142982 572704 142988 572716
rect 143040 572704 143046 572756
rect 227254 572704 227260 572756
rect 227312 572744 227318 572756
rect 251174 572744 251180 572756
rect 227312 572716 251180 572744
rect 227312 572704 227318 572716
rect 251174 572704 251180 572716
rect 251232 572704 251238 572756
rect 111794 571412 111800 571464
rect 111852 571452 111858 571464
rect 130470 571452 130476 571464
rect 111852 571424 130476 571452
rect 111852 571412 111858 571424
rect 130470 571412 130476 571424
rect 130528 571412 130534 571464
rect 111886 571344 111892 571396
rect 111944 571384 111950 571396
rect 133230 571384 133236 571396
rect 111944 571356 133236 571384
rect 111944 571344 111950 571356
rect 133230 571344 133236 571356
rect 133288 571344 133294 571396
rect 220354 571344 220360 571396
rect 220412 571384 220418 571396
rect 251174 571384 251180 571396
rect 220412 571356 251180 571384
rect 220412 571344 220418 571356
rect 251174 571344 251180 571356
rect 251232 571344 251238 571396
rect 111794 569984 111800 570036
rect 111852 570024 111858 570036
rect 122282 570024 122288 570036
rect 111852 569996 122288 570024
rect 111852 569984 111858 569996
rect 122282 569984 122288 569996
rect 122340 569984 122346 570036
rect 111978 569916 111984 569968
rect 112036 569956 112042 569968
rect 127618 569956 127624 569968
rect 112036 569928 127624 569956
rect 112036 569916 112042 569928
rect 127618 569916 127624 569928
rect 127676 569916 127682 569968
rect 238294 569916 238300 569968
rect 238352 569956 238358 569968
rect 251174 569956 251180 569968
rect 238352 569928 251180 569956
rect 238352 569916 238358 569928
rect 251174 569916 251180 569928
rect 251232 569916 251238 569968
rect 111886 568624 111892 568676
rect 111944 568664 111950 568676
rect 137278 568664 137284 568676
rect 111944 568636 137284 568664
rect 111944 568624 111950 568636
rect 137278 568624 137284 568636
rect 137336 568624 137342 568676
rect 234338 568624 234344 568676
rect 234396 568664 234402 568676
rect 251266 568664 251272 568676
rect 234396 568636 251272 568664
rect 234396 568624 234402 568636
rect 251266 568624 251272 568636
rect 251324 568624 251330 568676
rect 111794 568556 111800 568608
rect 111852 568596 111858 568608
rect 152734 568596 152740 568608
rect 111852 568568 152740 568596
rect 111852 568556 111858 568568
rect 152734 568556 152740 568568
rect 152792 568556 152798 568608
rect 225690 568556 225696 568608
rect 225748 568596 225754 568608
rect 251174 568596 251180 568608
rect 225748 568568 251180 568596
rect 225748 568556 225754 568568
rect 251174 568556 251180 568568
rect 251232 568556 251238 568608
rect 111794 567196 111800 567248
rect 111852 567236 111858 567248
rect 141602 567236 141608 567248
rect 111852 567208 141608 567236
rect 111852 567196 111858 567208
rect 141602 567196 141608 567208
rect 141660 567196 141666 567248
rect 220446 567196 220452 567248
rect 220504 567236 220510 567248
rect 251174 567236 251180 567248
rect 220504 567208 251180 567236
rect 220504 567196 220510 567208
rect 251174 567196 251180 567208
rect 251232 567196 251238 567248
rect 111794 565904 111800 565956
rect 111852 565944 111858 565956
rect 116578 565944 116584 565956
rect 111852 565916 116584 565944
rect 111852 565904 111858 565916
rect 116578 565904 116584 565916
rect 116636 565904 116642 565956
rect 3418 565836 3424 565888
rect 3476 565876 3482 565888
rect 29730 565876 29736 565888
rect 3476 565848 29736 565876
rect 3476 565836 3482 565848
rect 29730 565836 29736 565848
rect 29788 565836 29794 565888
rect 111886 565836 111892 565888
rect 111944 565876 111950 565888
rect 134702 565876 134708 565888
rect 111944 565848 134708 565876
rect 111944 565836 111950 565848
rect 134702 565836 134708 565848
rect 134760 565836 134766 565888
rect 236730 565836 236736 565888
rect 236788 565876 236794 565888
rect 251174 565876 251180 565888
rect 236788 565848 251180 565876
rect 236788 565836 236794 565848
rect 251174 565836 251180 565848
rect 251232 565836 251238 565888
rect 111794 564476 111800 564528
rect 111852 564516 111858 564528
rect 127710 564516 127716 564528
rect 111852 564488 127716 564516
rect 111852 564476 111858 564488
rect 127710 564476 127716 564488
rect 127768 564476 127774 564528
rect 111886 564408 111892 564460
rect 111944 564448 111950 564460
rect 130562 564448 130568 564460
rect 111944 564420 130568 564448
rect 111944 564408 111950 564420
rect 130562 564408 130568 564420
rect 130620 564408 130626 564460
rect 234430 564408 234436 564460
rect 234488 564448 234494 564460
rect 251174 564448 251180 564460
rect 234488 564420 251180 564448
rect 234488 564408 234494 564420
rect 251174 564408 251180 564420
rect 251232 564408 251238 564460
rect 112438 563660 112444 563712
rect 112496 563700 112502 563712
rect 122374 563700 122380 563712
rect 112496 563672 122380 563700
rect 112496 563660 112502 563672
rect 122374 563660 122380 563672
rect 122432 563660 122438 563712
rect 111794 563048 111800 563100
rect 111852 563088 111858 563100
rect 140130 563088 140136 563100
rect 111852 563060 140136 563088
rect 111852 563048 111858 563060
rect 140130 563048 140136 563060
rect 140188 563048 140194 563100
rect 242342 563048 242348 563100
rect 242400 563088 242406 563100
rect 251174 563088 251180 563100
rect 242400 563060 251180 563088
rect 242400 563048 242406 563060
rect 251174 563048 251180 563060
rect 251232 563048 251238 563100
rect 111978 562300 111984 562352
rect 112036 562340 112042 562352
rect 144270 562340 144276 562352
rect 112036 562312 144276 562340
rect 112036 562300 112042 562312
rect 144270 562300 144276 562312
rect 144328 562300 144334 562352
rect 111794 561688 111800 561740
rect 111852 561728 111858 561740
rect 115290 561728 115296 561740
rect 111852 561700 115296 561728
rect 111852 561688 111858 561700
rect 115290 561688 115296 561700
rect 115348 561688 115354 561740
rect 243814 561688 243820 561740
rect 243872 561728 243878 561740
rect 251174 561728 251180 561740
rect 243872 561700 251180 561728
rect 243872 561688 243878 561700
rect 251174 561688 251180 561700
rect 251232 561688 251238 561740
rect 111794 560260 111800 560312
rect 111852 560300 111858 560312
rect 140222 560300 140228 560312
rect 111852 560272 140228 560300
rect 111852 560260 111858 560272
rect 140222 560260 140228 560272
rect 140280 560260 140286 560312
rect 236822 560260 236828 560312
rect 236880 560300 236886 560312
rect 251174 560300 251180 560312
rect 236880 560272 251180 560300
rect 236880 560260 236886 560272
rect 251174 560260 251180 560272
rect 251232 560260 251238 560312
rect 111794 558968 111800 559020
rect 111852 559008 111858 559020
rect 115382 559008 115388 559020
rect 111852 558980 115388 559008
rect 111852 558968 111858 558980
rect 115382 558968 115388 558980
rect 115440 558968 115446 559020
rect 111886 558900 111892 558952
rect 111944 558940 111950 558952
rect 118050 558940 118056 558952
rect 111944 558912 118056 558940
rect 111944 558900 111950 558912
rect 118050 558900 118056 558912
rect 118108 558900 118114 558952
rect 234522 558900 234528 558952
rect 234580 558940 234586 558952
rect 251174 558940 251180 558952
rect 234580 558912 251180 558940
rect 234580 558900 234586 558912
rect 251174 558900 251180 558912
rect 251232 558900 251238 558952
rect 111794 557608 111800 557660
rect 111852 557648 111858 557660
rect 127802 557648 127808 557660
rect 111852 557620 127808 557648
rect 111852 557608 111858 557620
rect 127802 557608 127808 557620
rect 127860 557608 127866 557660
rect 245194 557608 245200 557660
rect 245252 557648 245258 557660
rect 251174 557648 251180 557660
rect 245252 557620 251180 557648
rect 245252 557608 245258 557620
rect 251174 557608 251180 557620
rect 251232 557608 251238 557660
rect 111886 557540 111892 557592
rect 111944 557580 111950 557592
rect 130654 557580 130660 557592
rect 111944 557552 130660 557580
rect 111944 557540 111950 557552
rect 130654 557540 130660 557552
rect 130712 557540 130718 557592
rect 223114 557540 223120 557592
rect 223172 557580 223178 557592
rect 251266 557580 251272 557592
rect 223172 557552 251272 557580
rect 223172 557540 223178 557552
rect 251266 557540 251272 557552
rect 251324 557540 251330 557592
rect 112622 556792 112628 556844
rect 112680 556832 112686 556844
rect 148410 556832 148416 556844
rect 112680 556804 148416 556832
rect 112680 556792 112686 556804
rect 148410 556792 148416 556804
rect 148468 556792 148474 556844
rect 111794 556180 111800 556232
rect 111852 556220 111858 556232
rect 147030 556220 147036 556232
rect 111852 556192 147036 556220
rect 111852 556180 111858 556192
rect 147030 556180 147036 556192
rect 147088 556180 147094 556232
rect 246758 556180 246764 556232
rect 246816 556220 246822 556232
rect 251174 556220 251180 556232
rect 246816 556192 251180 556220
rect 246816 556180 246822 556192
rect 251174 556180 251180 556192
rect 251232 556180 251238 556232
rect 111794 554888 111800 554940
rect 111852 554928 111858 554940
rect 115474 554928 115480 554940
rect 111852 554900 115480 554928
rect 111852 554888 111858 554900
rect 115474 554888 115480 554900
rect 115532 554888 115538 554940
rect 111886 554752 111892 554804
rect 111944 554792 111950 554804
rect 151170 554792 151176 554804
rect 111944 554764 151176 554792
rect 111944 554752 111950 554764
rect 151170 554752 151176 554764
rect 151228 554752 151234 554804
rect 236914 554752 236920 554804
rect 236972 554792 236978 554804
rect 251174 554792 251180 554804
rect 236972 554764 251180 554792
rect 236972 554752 236978 554764
rect 251174 554752 251180 554764
rect 251232 554752 251238 554804
rect 111978 554004 111984 554056
rect 112036 554044 112042 554056
rect 119338 554044 119344 554056
rect 112036 554016 119344 554044
rect 112036 554004 112042 554016
rect 119338 554004 119344 554016
rect 119396 554004 119402 554056
rect 111794 553392 111800 553444
rect 111852 553432 111858 553444
rect 138842 553432 138848 553444
rect 111852 553404 138848 553432
rect 111852 553392 111858 553404
rect 138842 553392 138848 553404
rect 138900 553392 138906 553444
rect 232866 553392 232872 553444
rect 232924 553432 232930 553444
rect 251174 553432 251180 553444
rect 232924 553404 251180 553432
rect 232924 553392 232930 553404
rect 251174 553392 251180 553404
rect 251232 553392 251238 553444
rect 112530 552644 112536 552696
rect 112588 552684 112594 552696
rect 113082 552684 113088 552696
rect 112588 552656 113088 552684
rect 112588 552644 112594 552656
rect 113082 552644 113088 552656
rect 113140 552644 113146 552696
rect 111886 552100 111892 552152
rect 111944 552140 111950 552152
rect 126238 552140 126244 552152
rect 111944 552112 126244 552140
rect 111944 552100 111950 552112
rect 126238 552100 126244 552112
rect 126296 552100 126302 552152
rect 111794 552032 111800 552084
rect 111852 552072 111858 552084
rect 149698 552072 149704 552084
rect 111852 552044 149704 552072
rect 111852 552032 111858 552044
rect 149698 552032 149704 552044
rect 149756 552032 149762 552084
rect 221918 552032 221924 552084
rect 221976 552072 221982 552084
rect 251174 552072 251180 552084
rect 221976 552044 251180 552072
rect 221976 552032 221982 552044
rect 251174 552032 251180 552044
rect 251232 552032 251238 552084
rect 111794 550672 111800 550724
rect 111852 550712 111858 550724
rect 116670 550712 116676 550724
rect 111852 550684 116676 550712
rect 111852 550672 111858 550684
rect 116670 550672 116676 550684
rect 116728 550672 116734 550724
rect 111886 550604 111892 550656
rect 111944 550644 111950 550656
rect 130746 550644 130752 550656
rect 111944 550616 130752 550644
rect 111944 550604 111950 550616
rect 130746 550604 130752 550616
rect 130804 550604 130810 550656
rect 220538 550604 220544 550656
rect 220596 550644 220602 550656
rect 251174 550644 251180 550656
rect 220596 550616 251180 550644
rect 220596 550604 220602 550616
rect 251174 550604 251180 550616
rect 251232 550604 251238 550656
rect 111794 549312 111800 549364
rect 111852 549352 111858 549364
rect 119430 549352 119436 549364
rect 111852 549324 119436 549352
rect 111852 549312 111858 549324
rect 119430 549312 119436 549324
rect 119488 549312 119494 549364
rect 111886 549244 111892 549296
rect 111944 549284 111950 549296
rect 153838 549284 153844 549296
rect 111944 549256 153844 549284
rect 111944 549244 111950 549256
rect 153838 549244 153844 549256
rect 153896 549244 153902 549296
rect 247954 549244 247960 549296
rect 248012 549284 248018 549296
rect 251174 549284 251180 549296
rect 248012 549256 251180 549284
rect 248012 549244 248018 549256
rect 251174 549244 251180 549256
rect 251232 549244 251238 549296
rect 112070 548496 112076 548548
rect 112128 548536 112134 548548
rect 143074 548536 143080 548548
rect 112128 548508 143080 548536
rect 112128 548496 112134 548508
rect 143074 548496 143080 548508
rect 143132 548496 143138 548548
rect 111794 548088 111800 548140
rect 111852 548128 111858 548140
rect 115566 548128 115572 548140
rect 111852 548100 115572 548128
rect 111852 548088 111858 548100
rect 115566 548088 115572 548100
rect 115624 548088 115630 548140
rect 235442 547952 235448 548004
rect 235500 547992 235506 548004
rect 251266 547992 251272 548004
rect 235500 547964 251272 547992
rect 235500 547952 235506 547964
rect 251266 547952 251272 547964
rect 251324 547952 251330 548004
rect 111886 547884 111892 547936
rect 111944 547924 111950 547936
rect 126514 547924 126520 547936
rect 111944 547896 126520 547924
rect 111944 547884 111950 547896
rect 126514 547884 126520 547896
rect 126572 547884 126578 547936
rect 232958 547884 232964 547936
rect 233016 547924 233022 547936
rect 251174 547924 251180 547936
rect 233016 547896 251180 547924
rect 233016 547884 233022 547896
rect 251174 547884 251180 547896
rect 251232 547884 251238 547936
rect 111794 546456 111800 546508
rect 111852 546496 111858 546508
rect 152826 546496 152832 546508
rect 111852 546468 152832 546496
rect 111852 546456 111858 546468
rect 152826 546456 152832 546468
rect 152884 546456 152890 546508
rect 231486 546456 231492 546508
rect 231544 546496 231550 546508
rect 251174 546496 251180 546508
rect 231544 546468 251180 546496
rect 231544 546456 231550 546468
rect 251174 546456 251180 546468
rect 251232 546456 251238 546508
rect 111886 545164 111892 545216
rect 111944 545204 111950 545216
rect 118142 545204 118148 545216
rect 111944 545176 118148 545204
rect 111944 545164 111950 545176
rect 118142 545164 118148 545176
rect 118200 545164 118206 545216
rect 111794 545096 111800 545148
rect 111852 545136 111858 545148
rect 131758 545136 131764 545148
rect 111852 545108 131764 545136
rect 111852 545096 111858 545108
rect 131758 545096 131764 545108
rect 131816 545096 131822 545148
rect 227346 545096 227352 545148
rect 227404 545136 227410 545148
rect 251174 545136 251180 545148
rect 227404 545108 251180 545136
rect 227404 545096 227410 545108
rect 251174 545096 251180 545108
rect 251232 545096 251238 545148
rect 111794 543736 111800 543788
rect 111852 543776 111858 543788
rect 144362 543776 144368 543788
rect 111852 543748 144368 543776
rect 111852 543736 111858 543748
rect 144362 543736 144368 543748
rect 144420 543736 144426 543788
rect 227438 543736 227444 543788
rect 227496 543776 227502 543788
rect 251174 543776 251180 543788
rect 227496 543748 251180 543776
rect 227496 543736 227502 543748
rect 251174 543736 251180 543748
rect 251232 543736 251238 543788
rect 116762 542988 116768 543040
rect 116820 543028 116826 543040
rect 155218 543028 155224 543040
rect 116820 543000 155224 543028
rect 116820 542988 116826 543000
rect 155218 542988 155224 543000
rect 155276 542988 155282 543040
rect 111886 542444 111892 542496
rect 111944 542484 111950 542496
rect 116854 542484 116860 542496
rect 111944 542456 116860 542484
rect 111944 542444 111950 542456
rect 116854 542444 116860 542456
rect 116912 542444 116918 542496
rect 111794 542376 111800 542428
rect 111852 542416 111858 542428
rect 119522 542416 119528 542428
rect 111852 542388 119528 542416
rect 111852 542376 111858 542388
rect 119522 542376 119528 542388
rect 119580 542376 119586 542428
rect 113082 541628 113088 541680
rect 113140 541668 113146 541680
rect 149790 541668 149796 541680
rect 113140 541640 149796 541668
rect 113140 541628 113146 541640
rect 149790 541628 149796 541640
rect 149848 541628 149854 541680
rect 111794 540948 111800 541000
rect 111852 540988 111858 541000
rect 116762 540988 116768 541000
rect 111852 540960 116768 540988
rect 111852 540948 111858 540960
rect 116762 540948 116768 540960
rect 116820 540948 116826 541000
rect 249518 540948 249524 541000
rect 249576 540988 249582 541000
rect 251174 540988 251180 541000
rect 249576 540960 251180 540988
rect 249576 540948 249582 540960
rect 251174 540948 251180 540960
rect 251232 540948 251238 541000
rect 111794 539588 111800 539640
rect 111852 539628 111858 539640
rect 137370 539628 137376 539640
rect 111852 539600 137376 539628
rect 111852 539588 111858 539600
rect 137370 539588 137376 539600
rect 137428 539588 137434 539640
rect 235534 539588 235540 539640
rect 235592 539628 235598 539640
rect 251174 539628 251180 539640
rect 235592 539600 251180 539628
rect 235592 539588 235598 539600
rect 251174 539588 251180 539600
rect 251232 539588 251238 539640
rect 111794 538296 111800 538348
rect 111852 538336 111858 538348
rect 127894 538336 127900 538348
rect 111852 538308 127900 538336
rect 111852 538296 111858 538308
rect 127894 538296 127900 538308
rect 127952 538296 127958 538348
rect 111886 538228 111892 538280
rect 111944 538268 111950 538280
rect 151262 538268 151268 538280
rect 111944 538240 151268 538268
rect 111944 538228 111950 538240
rect 151262 538228 151268 538240
rect 151320 538228 151326 538280
rect 235626 538228 235632 538280
rect 235684 538268 235690 538280
rect 251174 538268 251180 538280
rect 235684 538240 251180 538268
rect 235684 538228 235690 538240
rect 251174 538228 251180 538240
rect 251232 538228 251238 538280
rect 111794 536868 111800 536920
rect 111852 536908 111858 536920
rect 128998 536908 129004 536920
rect 111852 536880 129004 536908
rect 111852 536868 111858 536880
rect 128998 536868 129004 536880
rect 129056 536868 129062 536920
rect 111886 536800 111892 536852
rect 111944 536840 111950 536852
rect 131850 536840 131856 536852
rect 111944 536812 131856 536840
rect 111944 536800 111950 536812
rect 131850 536800 131856 536812
rect 131908 536800 131914 536852
rect 235718 536800 235724 536852
rect 235776 536840 235782 536852
rect 251174 536840 251180 536852
rect 235776 536812 251180 536840
rect 235776 536800 235782 536812
rect 251174 536800 251180 536812
rect 251232 536800 251238 536852
rect 111886 535508 111892 535560
rect 111944 535548 111950 535560
rect 148502 535548 148508 535560
rect 111944 535520 148508 535548
rect 111944 535508 111950 535520
rect 148502 535508 148508 535520
rect 148560 535508 148566 535560
rect 111794 535440 111800 535492
rect 111852 535480 111858 535492
rect 151354 535480 151360 535492
rect 111852 535452 151360 535480
rect 111852 535440 111858 535452
rect 151354 535440 151360 535452
rect 151412 535440 151418 535492
rect 220630 535440 220636 535492
rect 220688 535480 220694 535492
rect 251174 535480 251180 535492
rect 220688 535452 251180 535480
rect 220688 535440 220694 535452
rect 251174 535440 251180 535452
rect 251232 535440 251238 535492
rect 113082 534692 113088 534744
rect 113140 534732 113146 534744
rect 145558 534732 145564 534744
rect 113140 534704 145564 534732
rect 113140 534692 113146 534704
rect 145558 534692 145564 534704
rect 145616 534692 145622 534744
rect 111794 534080 111800 534132
rect 111852 534120 111858 534132
rect 143166 534120 143172 534132
rect 111852 534092 143172 534120
rect 111852 534080 111858 534092
rect 143166 534080 143172 534092
rect 143224 534080 143230 534132
rect 235810 534080 235816 534132
rect 235868 534120 235874 534132
rect 251174 534120 251180 534132
rect 235868 534092 251180 534120
rect 235868 534080 235874 534092
rect 251174 534080 251180 534092
rect 251232 534080 251238 534132
rect 111886 533740 111892 533792
rect 111944 533780 111950 533792
rect 116946 533780 116952 533792
rect 111944 533752 116952 533780
rect 111944 533740 111950 533752
rect 116946 533740 116952 533752
rect 117004 533740 117010 533792
rect 113082 532720 113088 532772
rect 113140 532760 113146 532772
rect 147122 532760 147128 532772
rect 113140 532732 147128 532760
rect 113140 532720 113146 532732
rect 147122 532720 147128 532732
rect 147180 532720 147186 532772
rect 113082 531360 113088 531412
rect 113140 531400 113146 531412
rect 138934 531400 138940 531412
rect 113140 531372 138940 531400
rect 113140 531360 113146 531372
rect 138934 531360 138940 531372
rect 138992 531360 138998 531412
rect 112254 531292 112260 531344
rect 112312 531332 112318 531344
rect 148594 531332 148600 531344
rect 112312 531304 148600 531332
rect 112312 531292 112318 531304
rect 148594 531292 148600 531304
rect 148652 531292 148658 531344
rect 112254 531156 112260 531208
rect 112312 531196 112318 531208
rect 112622 531196 112628 531208
rect 112312 531168 112628 531196
rect 112312 531156 112318 531168
rect 112622 531156 112628 531168
rect 112680 531156 112686 531208
rect 112438 530000 112444 530052
rect 112496 530000 112502 530052
rect 113082 530000 113088 530052
rect 113140 530040 113146 530052
rect 131942 530040 131948 530052
rect 113140 530012 131948 530040
rect 113140 530000 113146 530012
rect 131942 530000 131948 530012
rect 132000 530000 132006 530052
rect 112456 529848 112484 530000
rect 112622 529932 112628 529984
rect 112680 529972 112686 529984
rect 153930 529972 153936 529984
rect 112680 529944 153936 529972
rect 112680 529932 112686 529944
rect 153930 529932 153936 529944
rect 153988 529932 153994 529984
rect 112438 529796 112444 529848
rect 112496 529796 112502 529848
rect 249242 529320 249248 529372
rect 249300 529360 249306 529372
rect 580626 529360 580632 529372
rect 249300 529332 580632 529360
rect 249300 529320 249306 529332
rect 580626 529320 580632 529332
rect 580684 529320 580690 529372
rect 247678 529252 247684 529304
rect 247736 529292 247742 529304
rect 580166 529292 580172 529304
rect 247736 529264 580172 529292
rect 247736 529252 247742 529264
rect 580166 529252 580172 529264
rect 580224 529252 580230 529304
rect 112254 529184 112260 529236
rect 112312 529224 112318 529236
rect 123846 529224 123852 529236
rect 112312 529196 123852 529224
rect 112312 529184 112318 529196
rect 123846 529184 123852 529196
rect 123904 529184 123910 529236
rect 132034 529184 132040 529236
rect 132092 529224 132098 529236
rect 155310 529224 155316 529236
rect 132092 529196 155316 529224
rect 132092 529184 132098 529196
rect 155310 529184 155316 529196
rect 155368 529184 155374 529236
rect 240870 529184 240876 529236
rect 240928 529224 240934 529236
rect 580534 529224 580540 529236
rect 240928 529196 580540 529224
rect 240928 529184 240934 529196
rect 580534 529184 580540 529196
rect 580592 529184 580598 529236
rect 112346 528572 112352 528624
rect 112404 528612 112410 528624
rect 124858 528612 124864 528624
rect 112404 528584 124864 528612
rect 112404 528572 112410 528584
rect 124858 528572 124864 528584
rect 124916 528572 124922 528624
rect 111794 527212 111800 527264
rect 111852 527252 111858 527264
rect 114094 527252 114100 527264
rect 111852 527224 114100 527252
rect 111852 527212 111858 527224
rect 114094 527212 114100 527224
rect 114152 527212 114158 527264
rect 2958 527144 2964 527196
rect 3016 527184 3022 527196
rect 29822 527184 29828 527196
rect 3016 527156 29828 527184
rect 3016 527144 3022 527156
rect 29822 527144 29828 527156
rect 29880 527144 29886 527196
rect 112346 525852 112352 525904
rect 112404 525892 112410 525904
rect 139026 525892 139032 525904
rect 112404 525864 139032 525892
rect 112404 525852 112410 525864
rect 139026 525852 139032 525864
rect 139084 525852 139090 525904
rect 113082 525784 113088 525836
rect 113140 525824 113146 525836
rect 144454 525824 144460 525836
rect 113140 525796 144460 525824
rect 113140 525784 113146 525796
rect 144454 525784 144460 525796
rect 144512 525784 144518 525836
rect 112254 525716 112260 525768
rect 112312 525756 112318 525768
rect 117038 525756 117044 525768
rect 112312 525728 117044 525756
rect 112312 525716 112318 525728
rect 117038 525716 117044 525728
rect 117096 525716 117102 525768
rect 112070 524424 112076 524476
rect 112128 524464 112134 524476
rect 147214 524464 147220 524476
rect 112128 524436 147220 524464
rect 112128 524424 112134 524436
rect 147214 524424 147220 524436
rect 147272 524424 147278 524476
rect 221550 524424 221556 524476
rect 221608 524464 221614 524476
rect 580166 524464 580172 524476
rect 221608 524436 580172 524464
rect 221608 524424 221614 524436
rect 580166 524424 580172 524436
rect 580224 524424 580230 524476
rect 111886 523064 111892 523116
rect 111944 523104 111950 523116
rect 132034 523104 132040 523116
rect 111944 523076 132040 523104
rect 111944 523064 111950 523076
rect 132034 523064 132040 523076
rect 132092 523064 132098 523116
rect 111794 522996 111800 523048
rect 111852 523036 111858 523048
rect 143258 523036 143264 523048
rect 111852 523008 143264 523036
rect 111852 522996 111858 523008
rect 143258 522996 143264 523008
rect 143316 522996 143322 523048
rect 111886 521704 111892 521756
rect 111944 521744 111950 521756
rect 118234 521744 118240 521756
rect 111944 521716 118240 521744
rect 111944 521704 111950 521716
rect 118234 521704 118240 521716
rect 118292 521704 118298 521756
rect 111794 521636 111800 521688
rect 111852 521676 111858 521688
rect 126330 521676 126336 521688
rect 111852 521648 126336 521676
rect 111852 521636 111858 521648
rect 126330 521636 126336 521648
rect 126388 521636 126394 521688
rect 112898 521160 112904 521212
rect 112956 521200 112962 521212
rect 113174 521200 113180 521212
rect 112956 521172 113180 521200
rect 112956 521160 112962 521172
rect 113174 521160 113180 521172
rect 113232 521160 113238 521212
rect 113082 520888 113088 520940
rect 113140 520928 113146 520940
rect 149882 520928 149888 520940
rect 113140 520900 149888 520928
rect 113140 520888 113146 520900
rect 149882 520888 149888 520900
rect 149940 520888 149946 520940
rect 111794 520344 111800 520396
rect 111852 520384 111858 520396
rect 120810 520384 120816 520396
rect 111852 520356 120816 520384
rect 111852 520344 111858 520356
rect 120810 520344 120816 520356
rect 120868 520344 120874 520396
rect 111886 520276 111892 520328
rect 111944 520316 111950 520328
rect 124950 520316 124956 520328
rect 111944 520288 124956 520316
rect 111944 520276 111950 520288
rect 124950 520276 124956 520288
rect 125008 520276 125014 520328
rect 111794 519596 111800 519648
rect 111852 519636 111858 519648
rect 118326 519636 118332 519648
rect 111852 519608 118332 519636
rect 111852 519596 111858 519608
rect 118326 519596 118332 519608
rect 118384 519596 118390 519648
rect 112806 519528 112812 519580
rect 112864 519568 112870 519580
rect 145742 519568 145748 519580
rect 112864 519540 145748 519568
rect 112864 519528 112870 519540
rect 145742 519528 145748 519540
rect 145800 519528 145806 519580
rect 112346 518168 112352 518220
rect 112404 518208 112410 518220
rect 154022 518208 154028 518220
rect 112404 518180 154028 518208
rect 112404 518168 112410 518180
rect 154022 518168 154028 518180
rect 154080 518168 154086 518220
rect 111794 517488 111800 517540
rect 111852 517528 111858 517540
rect 144546 517528 144552 517540
rect 111852 517500 144552 517528
rect 111852 517488 111858 517500
rect 144546 517488 144552 517500
rect 144604 517488 144610 517540
rect 111886 516196 111892 516248
rect 111944 516236 111950 516248
rect 119706 516236 119712 516248
rect 111944 516208 119712 516236
rect 111944 516196 111950 516208
rect 119706 516196 119712 516208
rect 119764 516196 119770 516248
rect 111794 516128 111800 516180
rect 111852 516168 111858 516180
rect 140314 516168 140320 516180
rect 111852 516140 140320 516168
rect 111852 516128 111858 516140
rect 140314 516128 140320 516140
rect 140372 516128 140378 516180
rect 113082 515380 113088 515432
rect 113140 515420 113146 515432
rect 130838 515420 130844 515432
rect 113140 515392 130844 515420
rect 113140 515380 113146 515392
rect 130838 515380 130844 515392
rect 130896 515380 130902 515432
rect 111794 514836 111800 514888
rect 111852 514876 111858 514888
rect 114186 514876 114192 514888
rect 111852 514848 114192 514876
rect 111852 514836 111858 514848
rect 114186 514836 114192 514848
rect 114244 514836 114250 514888
rect 3510 514768 3516 514820
rect 3568 514808 3574 514820
rect 29914 514808 29920 514820
rect 3568 514780 29920 514808
rect 3568 514768 3574 514780
rect 29914 514768 29920 514780
rect 29972 514768 29978 514820
rect 111886 514768 111892 514820
rect 111944 514808 111950 514820
rect 120902 514808 120908 514820
rect 111944 514780 120908 514808
rect 111944 514768 111950 514780
rect 120902 514768 120908 514780
rect 120960 514768 120966 514820
rect 111794 513408 111800 513460
rect 111852 513448 111858 513460
rect 125042 513448 125048 513460
rect 111852 513420 125048 513448
rect 111852 513408 111858 513420
rect 125042 513408 125048 513420
rect 125100 513408 125106 513460
rect 111886 513340 111892 513392
rect 111944 513380 111950 513392
rect 145650 513380 145656 513392
rect 111944 513352 145656 513380
rect 111944 513340 111950 513352
rect 145650 513340 145656 513352
rect 145708 513340 145714 513392
rect 112254 512592 112260 512644
rect 112312 512632 112318 512644
rect 147306 512632 147312 512644
rect 112312 512604 147312 512632
rect 112312 512592 112318 512604
rect 147306 512592 147312 512604
rect 147364 512592 147370 512644
rect 111794 511980 111800 512032
rect 111852 512020 111858 512032
rect 139118 512020 139124 512032
rect 111852 511992 139124 512020
rect 111852 511980 111858 511992
rect 139118 511980 139124 511992
rect 139176 511980 139182 512032
rect 111886 510688 111892 510740
rect 111944 510728 111950 510740
rect 117130 510728 117136 510740
rect 111944 510700 117136 510728
rect 111944 510688 111950 510700
rect 117130 510688 117136 510700
rect 117188 510688 117194 510740
rect 111794 510620 111800 510672
rect 111852 510660 111858 510672
rect 141694 510660 141700 510672
rect 111852 510632 141700 510660
rect 111852 510620 111858 510632
rect 141694 510620 141700 510632
rect 141752 510620 141758 510672
rect 234062 510620 234068 510672
rect 234120 510660 234126 510672
rect 580166 510660 580172 510672
rect 234120 510632 580172 510660
rect 234120 510620 234126 510632
rect 580166 510620 580172 510632
rect 580224 510620 580230 510672
rect 111978 509872 111984 509924
rect 112036 509912 112042 509924
rect 120994 509912 121000 509924
rect 112036 509884 121000 509912
rect 112036 509872 112042 509884
rect 120994 509872 121000 509884
rect 121052 509872 121058 509924
rect 111794 509260 111800 509312
rect 111852 509300 111858 509312
rect 143350 509300 143356 509312
rect 111852 509272 143356 509300
rect 111852 509260 111858 509272
rect 143350 509260 143356 509272
rect 143408 509260 143414 509312
rect 112990 508512 112996 508564
rect 113048 508552 113054 508564
rect 122650 508552 122656 508564
rect 113048 508524 122656 508552
rect 113048 508512 113054 508524
rect 122650 508512 122656 508524
rect 122708 508512 122714 508564
rect 111886 507900 111892 507952
rect 111944 507940 111950 507952
rect 126606 507940 126612 507952
rect 111944 507912 126612 507940
rect 111944 507900 111950 507912
rect 126606 507900 126612 507912
rect 126664 507900 126670 507952
rect 111794 507832 111800 507884
rect 111852 507872 111858 507884
rect 141786 507872 141792 507884
rect 111852 507844 141792 507872
rect 111852 507832 111858 507844
rect 141786 507832 141792 507844
rect 141844 507832 141850 507884
rect 111794 506472 111800 506524
rect 111852 506512 111858 506524
rect 129090 506512 129096 506524
rect 111852 506484 129096 506512
rect 111852 506472 111858 506484
rect 129090 506472 129096 506484
rect 129148 506472 129154 506524
rect 111886 505724 111892 505776
rect 111944 505764 111950 505776
rect 147398 505764 147404 505776
rect 111944 505736 147404 505764
rect 111944 505724 111950 505736
rect 147398 505724 147404 505736
rect 147456 505724 147462 505776
rect 111794 505112 111800 505164
rect 111852 505152 111858 505164
rect 126422 505152 126428 505164
rect 111852 505124 126428 505152
rect 111852 505112 111858 505124
rect 126422 505112 126428 505124
rect 126480 505112 126486 505164
rect 126514 504364 126520 504416
rect 126572 504404 126578 504416
rect 155494 504404 155500 504416
rect 126572 504376 155500 504404
rect 126572 504364 126578 504376
rect 155494 504364 155500 504376
rect 155552 504364 155558 504416
rect 111794 503888 111800 503940
rect 111852 503928 111858 503940
rect 114278 503928 114284 503940
rect 111852 503900 114284 503928
rect 111852 503888 111858 503900
rect 114278 503888 114284 503900
rect 114336 503888 114342 503940
rect 111886 503684 111892 503736
rect 111944 503724 111950 503736
rect 121086 503724 121092 503736
rect 111944 503696 121092 503724
rect 111944 503684 111950 503696
rect 121086 503684 121092 503696
rect 121144 503684 121150 503736
rect 111794 502392 111800 502444
rect 111852 502432 111858 502444
rect 140406 502432 140412 502444
rect 111852 502404 140412 502432
rect 111852 502392 111858 502404
rect 140406 502392 140412 502404
rect 140464 502392 140470 502444
rect 111886 502324 111892 502376
rect 111944 502364 111950 502376
rect 140498 502364 140504 502376
rect 111944 502336 140504 502364
rect 111944 502324 111950 502336
rect 140498 502324 140504 502336
rect 140556 502324 140562 502376
rect 111794 500964 111800 501016
rect 111852 501004 111858 501016
rect 148686 501004 148692 501016
rect 111852 500976 148692 501004
rect 111852 500964 111858 500976
rect 148686 500964 148692 500976
rect 148744 500964 148750 501016
rect 111794 499672 111800 499724
rect 111852 499712 111858 499724
rect 115658 499712 115664 499724
rect 111852 499684 115664 499712
rect 111852 499672 111858 499684
rect 115658 499672 115664 499684
rect 115716 499672 115722 499724
rect 111978 499536 111984 499588
rect 112036 499576 112042 499588
rect 133322 499576 133328 499588
rect 112036 499548 133328 499576
rect 112036 499536 112042 499548
rect 133322 499536 133328 499548
rect 133380 499536 133386 499588
rect 111886 498788 111892 498840
rect 111944 498828 111950 498840
rect 141878 498828 141884 498840
rect 111944 498800 141884 498828
rect 111944 498788 111950 498800
rect 141878 498788 141884 498800
rect 141936 498788 141942 498840
rect 111794 498176 111800 498228
rect 111852 498216 111858 498228
rect 127986 498216 127992 498228
rect 111852 498188 127992 498216
rect 111852 498176 111858 498188
rect 127986 498176 127992 498188
rect 128044 498176 128050 498228
rect 126606 497428 126612 497480
rect 126664 497468 126670 497480
rect 155402 497468 155408 497480
rect 126664 497440 155408 497468
rect 126664 497428 126670 497440
rect 155402 497428 155408 497440
rect 155460 497428 155466 497480
rect 233050 497428 233056 497480
rect 233108 497468 233114 497480
rect 252186 497468 252192 497480
rect 233108 497440 252192 497468
rect 233108 497428 233114 497440
rect 252186 497428 252192 497440
rect 252244 497428 252250 497480
rect 111794 496884 111800 496936
rect 111852 496924 111858 496936
rect 119798 496924 119804 496936
rect 111852 496896 119804 496924
rect 111852 496884 111858 496896
rect 119798 496884 119804 496896
rect 119856 496884 119862 496936
rect 111886 496816 111892 496868
rect 111944 496856 111950 496868
rect 126790 496856 126796 496868
rect 111944 496828 126796 496856
rect 111944 496816 111950 496828
rect 126790 496816 126796 496828
rect 126848 496816 126854 496868
rect 111978 496068 111984 496120
rect 112036 496108 112042 496120
rect 135990 496108 135996 496120
rect 112036 496080 135996 496108
rect 112036 496068 112042 496080
rect 135990 496068 135996 496080
rect 136048 496068 136054 496120
rect 111794 495728 111800 495780
rect 111852 495768 111858 495780
rect 115750 495768 115756 495780
rect 111852 495740 115756 495768
rect 111852 495728 111858 495740
rect 115750 495728 115756 495740
rect 115808 495728 115814 495780
rect 111886 495456 111892 495508
rect 111944 495496 111950 495508
rect 121178 495496 121184 495508
rect 111944 495468 121184 495496
rect 111944 495456 111950 495468
rect 121178 495456 121184 495468
rect 121236 495456 121242 495508
rect 225782 495456 225788 495508
rect 225840 495496 225846 495508
rect 251174 495496 251180 495508
rect 225840 495468 251180 495496
rect 225840 495456 225846 495468
rect 251174 495456 251180 495468
rect 251232 495456 251238 495508
rect 111794 495048 111800 495100
rect 111852 495088 111858 495100
rect 114370 495088 114376 495100
rect 111852 495060 114376 495088
rect 111852 495048 111858 495060
rect 114370 495048 114376 495060
rect 114428 495048 114434 495100
rect 111794 494028 111800 494080
rect 111852 494068 111858 494080
rect 148778 494068 148784 494080
rect 111852 494040 148784 494068
rect 111852 494028 111858 494040
rect 148778 494028 148784 494040
rect 148836 494028 148842 494080
rect 225874 494028 225880 494080
rect 225932 494068 225938 494080
rect 251174 494068 251180 494080
rect 225932 494040 251180 494068
rect 225932 494028 225938 494040
rect 251174 494028 251180 494040
rect 251232 494028 251238 494080
rect 111794 492668 111800 492720
rect 111852 492708 111858 492720
rect 151446 492708 151452 492720
rect 111852 492680 151452 492708
rect 111852 492668 111858 492680
rect 151446 492668 151452 492680
rect 151504 492668 151510 492720
rect 243906 492668 243912 492720
rect 243964 492708 243970 492720
rect 251174 492708 251180 492720
rect 243964 492680 251180 492708
rect 243964 492668 243970 492680
rect 251174 492668 251180 492680
rect 251232 492668 251238 492720
rect 111794 491376 111800 491428
rect 111852 491416 111858 491428
rect 122466 491416 122472 491428
rect 111852 491388 122472 491416
rect 111852 491376 111858 491388
rect 122466 491376 122472 491388
rect 122524 491376 122530 491428
rect 111886 491308 111892 491360
rect 111944 491348 111950 491360
rect 126698 491348 126704 491360
rect 111944 491320 126704 491348
rect 111944 491308 111950 491320
rect 126698 491308 126704 491320
rect 126756 491308 126762 491360
rect 225966 491308 225972 491360
rect 226024 491348 226030 491360
rect 251174 491348 251180 491360
rect 226024 491320 251180 491348
rect 226024 491308 226030 491320
rect 251174 491308 251180 491320
rect 251232 491308 251238 491360
rect 111794 489948 111800 490000
rect 111852 489988 111858 490000
rect 128078 489988 128084 490000
rect 111852 489960 128084 489988
rect 111852 489948 111858 489960
rect 128078 489948 128084 489960
rect 128136 489948 128142 490000
rect 111886 489880 111892 489932
rect 111944 489920 111950 489932
rect 129182 489920 129188 489932
rect 111944 489892 129188 489920
rect 111944 489880 111950 489892
rect 129182 489880 129188 489892
rect 129240 489880 129246 489932
rect 224402 489880 224408 489932
rect 224460 489920 224466 489932
rect 251174 489920 251180 489932
rect 224460 489892 251180 489920
rect 224460 489880 224466 489892
rect 251174 489880 251180 489892
rect 251232 489880 251238 489932
rect 111886 488588 111892 488640
rect 111944 488628 111950 488640
rect 126514 488628 126520 488640
rect 111944 488600 126520 488628
rect 111944 488588 111950 488600
rect 126514 488588 126520 488600
rect 126572 488588 126578 488640
rect 111794 488520 111800 488572
rect 111852 488560 111858 488572
rect 137462 488560 137468 488572
rect 111852 488532 137468 488560
rect 111852 488520 111858 488532
rect 137462 488520 137468 488532
rect 137520 488520 137526 488572
rect 241146 488520 241152 488572
rect 241204 488560 241210 488572
rect 251174 488560 251180 488572
rect 241204 488532 251180 488560
rect 241204 488520 241210 488532
rect 251174 488520 251180 488532
rect 251232 488520 251238 488572
rect 111794 487228 111800 487280
rect 111852 487268 111858 487280
rect 118418 487268 118424 487280
rect 111852 487240 118424 487268
rect 111852 487228 111858 487240
rect 118418 487228 118424 487240
rect 118476 487228 118482 487280
rect 111886 487160 111892 487212
rect 111944 487200 111950 487212
rect 144638 487200 144644 487212
rect 111944 487172 144644 487200
rect 111944 487160 111950 487172
rect 144638 487160 144644 487172
rect 144696 487160 144702 487212
rect 238386 487160 238392 487212
rect 238444 487200 238450 487212
rect 251174 487200 251180 487212
rect 238444 487172 251180 487200
rect 238444 487160 238450 487172
rect 251174 487160 251180 487172
rect 251232 487160 251238 487212
rect 111886 485868 111892 485920
rect 111944 485908 111950 485920
rect 137554 485908 137560 485920
rect 111944 485880 137560 485908
rect 111944 485868 111950 485880
rect 137554 485868 137560 485880
rect 137612 485868 137618 485920
rect 111794 485800 111800 485852
rect 111852 485840 111858 485852
rect 151538 485840 151544 485852
rect 111852 485812 151544 485840
rect 111852 485800 111858 485812
rect 151538 485800 151544 485812
rect 151596 485800 151602 485852
rect 246850 485800 246856 485852
rect 246908 485840 246914 485852
rect 251174 485840 251180 485852
rect 246908 485812 251180 485840
rect 246908 485800 246914 485812
rect 251174 485800 251180 485812
rect 251232 485800 251238 485852
rect 113082 485052 113088 485104
rect 113140 485092 113146 485104
rect 140590 485092 140596 485104
rect 113140 485064 140596 485092
rect 113140 485052 113146 485064
rect 140590 485052 140596 485064
rect 140648 485052 140654 485104
rect 111794 484372 111800 484424
rect 111852 484412 111858 484424
rect 134794 484412 134800 484424
rect 111852 484384 134800 484412
rect 111852 484372 111858 484384
rect 134794 484372 134800 484384
rect 134852 484372 134858 484424
rect 224494 484372 224500 484424
rect 224552 484412 224558 484424
rect 251174 484412 251180 484424
rect 224552 484384 251180 484412
rect 224552 484372 224558 484384
rect 251174 484372 251180 484384
rect 251232 484372 251238 484424
rect 111794 483080 111800 483132
rect 111852 483120 111858 483132
rect 123938 483120 123944 483132
rect 111852 483092 123944 483120
rect 111852 483080 111858 483092
rect 123938 483080 123944 483092
rect 123996 483080 124002 483132
rect 111886 483012 111892 483064
rect 111944 483052 111950 483064
rect 133414 483052 133420 483064
rect 111944 483024 133420 483052
rect 111944 483012 111950 483024
rect 133414 483012 133420 483024
rect 133472 483012 133478 483064
rect 224586 483012 224592 483064
rect 224644 483052 224650 483064
rect 251174 483052 251180 483064
rect 224644 483024 251180 483052
rect 224644 483012 224650 483024
rect 251174 483012 251180 483024
rect 251232 483012 251238 483064
rect 111794 481720 111800 481772
rect 111852 481760 111858 481772
rect 128170 481760 128176 481772
rect 111852 481732 128176 481760
rect 111852 481720 111858 481732
rect 128170 481720 128176 481732
rect 128228 481720 128234 481772
rect 111886 481652 111892 481704
rect 111944 481692 111950 481704
rect 129274 481692 129280 481704
rect 111944 481664 129280 481692
rect 111944 481652 111950 481664
rect 129274 481652 129280 481664
rect 129332 481652 129338 481704
rect 224770 481652 224776 481704
rect 224828 481692 224834 481704
rect 251174 481692 251180 481704
rect 224828 481664 251180 481692
rect 224828 481652 224834 481664
rect 251174 481652 251180 481664
rect 251232 481652 251238 481704
rect 126698 480904 126704 480956
rect 126756 480944 126762 480956
rect 155586 480944 155592 480956
rect 126756 480916 155592 480944
rect 126756 480904 126762 480916
rect 155586 480904 155592 480916
rect 155644 480904 155650 480956
rect 111794 480292 111800 480344
rect 111852 480332 111858 480344
rect 124030 480332 124036 480344
rect 111852 480304 124036 480332
rect 111852 480292 111858 480304
rect 124030 480292 124036 480304
rect 124088 480292 124094 480344
rect 111886 480224 111892 480276
rect 111944 480264 111950 480276
rect 126606 480264 126612 480276
rect 111944 480236 126612 480264
rect 111944 480224 111950 480236
rect 126606 480224 126612 480236
rect 126664 480224 126670 480276
rect 224678 480224 224684 480276
rect 224736 480264 224742 480276
rect 251174 480264 251180 480276
rect 224736 480236 251180 480264
rect 224736 480224 224742 480236
rect 251174 480224 251180 480236
rect 251232 480224 251238 480276
rect 239766 479476 239772 479528
rect 239824 479516 239830 479528
rect 252370 479516 252376 479528
rect 239824 479488 252376 479516
rect 239824 479476 239830 479488
rect 252370 479476 252376 479488
rect 252428 479476 252434 479528
rect 111794 478932 111800 478984
rect 111852 478972 111858 478984
rect 118510 478972 118516 478984
rect 111852 478944 118516 478972
rect 111852 478932 111858 478944
rect 118510 478932 118516 478944
rect 118568 478932 118574 478984
rect 111886 478864 111892 478916
rect 111944 478904 111950 478916
rect 145834 478904 145840 478916
rect 111944 478876 145840 478904
rect 111944 478864 111950 478876
rect 145834 478864 145840 478876
rect 145892 478864 145898 478916
rect 249610 478864 249616 478916
rect 249668 478904 249674 478916
rect 251174 478904 251180 478916
rect 249668 478876 251180 478904
rect 249668 478864 249674 478876
rect 251174 478864 251180 478876
rect 251232 478864 251238 478916
rect 111794 477640 111800 477692
rect 111852 477680 111858 477692
rect 114462 477680 114468 477692
rect 111852 477652 114468 477680
rect 111852 477640 111858 477652
rect 114462 477640 114468 477652
rect 114520 477640 114526 477692
rect 111886 477504 111892 477556
rect 111944 477544 111950 477556
rect 143442 477544 143448 477556
rect 111944 477516 143448 477544
rect 111944 477504 111950 477516
rect 143442 477504 143448 477516
rect 143500 477504 143506 477556
rect 223298 477504 223304 477556
rect 223356 477544 223362 477556
rect 251174 477544 251180 477556
rect 223356 477516 251180 477544
rect 223356 477504 223362 477516
rect 251174 477504 251180 477516
rect 251232 477504 251238 477556
rect 112346 476756 112352 476808
rect 112404 476796 112410 476808
rect 125226 476796 125232 476808
rect 112404 476768 125232 476796
rect 112404 476756 112410 476768
rect 125226 476756 125232 476768
rect 125284 476756 125290 476808
rect 111794 476076 111800 476128
rect 111852 476116 111858 476128
rect 136082 476116 136088 476128
rect 111852 476088 136088 476116
rect 111852 476076 111858 476088
rect 136082 476076 136088 476088
rect 136140 476076 136146 476128
rect 223206 476076 223212 476128
rect 223264 476116 223270 476128
rect 251174 476116 251180 476128
rect 223264 476088 251180 476116
rect 223264 476076 223270 476088
rect 251174 476076 251180 476088
rect 251232 476076 251238 476128
rect 111794 474784 111800 474836
rect 111852 474824 111858 474836
rect 132126 474824 132132 474836
rect 111852 474796 132132 474824
rect 111852 474784 111858 474796
rect 132126 474784 132132 474796
rect 132184 474784 132190 474836
rect 111886 474716 111892 474768
rect 111944 474756 111950 474768
rect 133506 474756 133512 474768
rect 111944 474728 133512 474756
rect 111944 474716 111950 474728
rect 133506 474716 133512 474728
rect 133564 474716 133570 474768
rect 227530 474716 227536 474768
rect 227588 474756 227594 474768
rect 251174 474756 251180 474768
rect 227588 474728 251180 474756
rect 227588 474716 227594 474728
rect 251174 474716 251180 474728
rect 251232 474716 251238 474768
rect 111794 474036 111800 474088
rect 111852 474076 111858 474088
rect 115842 474076 115848 474088
rect 111852 474048 115848 474076
rect 111852 474036 111858 474048
rect 115842 474036 115848 474048
rect 115900 474036 115906 474088
rect 111794 473424 111800 473476
rect 111852 473464 111858 473476
rect 128262 473464 128268 473476
rect 111852 473436 128268 473464
rect 111852 473424 111858 473436
rect 128262 473424 128268 473436
rect 128320 473424 128326 473476
rect 111886 473356 111892 473408
rect 111944 473396 111950 473408
rect 129366 473396 129372 473408
rect 111944 473368 129372 473396
rect 111944 473356 111950 473368
rect 129366 473356 129372 473368
rect 129424 473356 129430 473408
rect 242434 473356 242440 473408
rect 242492 473396 242498 473408
rect 251174 473396 251180 473408
rect 242492 473368 251180 473396
rect 242492 473356 242498 473368
rect 251174 473356 251180 473368
rect 251232 473356 251238 473408
rect 111794 472064 111800 472116
rect 111852 472104 111858 472116
rect 122558 472104 122564 472116
rect 111852 472076 122564 472104
rect 111852 472064 111858 472076
rect 122558 472064 122564 472076
rect 122616 472064 122622 472116
rect 111886 471996 111892 472048
rect 111944 472036 111950 472048
rect 126698 472036 126704 472048
rect 111944 472008 126704 472036
rect 111944 471996 111950 472008
rect 126698 471996 126704 472008
rect 126756 471996 126762 472048
rect 224862 471996 224868 472048
rect 224920 472036 224926 472048
rect 251174 472036 251180 472048
rect 224920 472008 251180 472036
rect 224920 471996 224926 472008
rect 251174 471996 251180 472008
rect 251232 471996 251238 472048
rect 111886 470636 111892 470688
rect 111944 470676 111950 470688
rect 141970 470676 141976 470688
rect 111944 470648 141976 470676
rect 111944 470636 111950 470648
rect 141970 470636 141976 470648
rect 142028 470636 142034 470688
rect 111794 470568 111800 470620
rect 111852 470608 111858 470620
rect 147490 470608 147496 470620
rect 111852 470580 147496 470608
rect 111852 470568 111858 470580
rect 147490 470568 147496 470580
rect 147548 470568 147554 470620
rect 230106 470568 230112 470620
rect 230164 470608 230170 470620
rect 251174 470608 251180 470620
rect 230164 470580 251180 470608
rect 230164 470568 230170 470580
rect 251174 470568 251180 470580
rect 251232 470568 251238 470620
rect 111794 469344 111800 469396
rect 111852 469384 111858 469396
rect 115106 469384 115112 469396
rect 111852 469356 115112 469384
rect 111852 469344 111858 469356
rect 115106 469344 115112 469356
rect 115164 469344 115170 469396
rect 245286 469276 245292 469328
rect 245344 469316 245350 469328
rect 251174 469316 251180 469328
rect 245344 469288 251180 469316
rect 245344 469276 245350 469288
rect 251174 469276 251180 469288
rect 251232 469276 251238 469328
rect 111794 469208 111800 469260
rect 111852 469248 111858 469260
rect 154114 469248 154120 469260
rect 111852 469220 154120 469248
rect 111852 469208 111858 469220
rect 154114 469208 154120 469220
rect 154172 469208 154178 469260
rect 227622 469208 227628 469260
rect 227680 469248 227686 469260
rect 251266 469248 251272 469260
rect 227680 469220 251272 469248
rect 227680 469208 227686 469220
rect 251266 469208 251272 469220
rect 251324 469208 251330 469260
rect 111794 467916 111800 467968
rect 111852 467956 111858 467968
rect 117222 467956 117228 467968
rect 111852 467928 117228 467956
rect 111852 467916 111858 467928
rect 117222 467916 117228 467928
rect 117280 467916 117286 467968
rect 111886 467848 111892 467900
rect 111944 467888 111950 467900
rect 152918 467888 152924 467900
rect 111944 467860 152924 467888
rect 111944 467848 111950 467860
rect 152918 467848 152924 467860
rect 152976 467848 152982 467900
rect 111794 466488 111800 466540
rect 111852 466528 111858 466540
rect 132218 466528 132224 466540
rect 111852 466500 132224 466528
rect 111852 466488 111858 466500
rect 132218 466488 132224 466500
rect 132276 466488 132282 466540
rect 111886 466420 111892 466472
rect 111944 466460 111950 466472
rect 137646 466460 137652 466472
rect 111944 466432 137652 466460
rect 111944 466420 111950 466432
rect 137646 466420 137652 466432
rect 137704 466420 137710 466472
rect 230198 466420 230204 466472
rect 230256 466460 230262 466472
rect 251174 466460 251180 466472
rect 230256 466432 251180 466460
rect 230256 466420 230262 466432
rect 251174 466420 251180 466432
rect 251232 466420 251238 466472
rect 111886 465128 111892 465180
rect 111944 465168 111950 465180
rect 125134 465168 125140 465180
rect 111944 465140 125140 465168
rect 111944 465128 111950 465140
rect 125134 465128 125140 465140
rect 125192 465128 125198 465180
rect 111794 465060 111800 465112
rect 111852 465100 111858 465112
rect 151630 465100 151636 465112
rect 111852 465072 151636 465100
rect 111852 465060 111858 465072
rect 151630 465060 151636 465072
rect 151688 465060 151694 465112
rect 249702 465060 249708 465112
rect 249760 465100 249766 465112
rect 251634 465100 251640 465112
rect 249760 465072 251640 465100
rect 249760 465060 249766 465072
rect 251634 465060 251640 465072
rect 251692 465060 251698 465112
rect 111794 463768 111800 463820
rect 111852 463808 111858 463820
rect 126882 463808 126888 463820
rect 111852 463780 126888 463808
rect 111852 463768 111858 463780
rect 126882 463768 126888 463780
rect 126940 463768 126946 463820
rect 111886 463700 111892 463752
rect 111944 463740 111950 463752
rect 149974 463740 149980 463752
rect 111944 463712 149980 463740
rect 111944 463700 111950 463712
rect 149974 463700 149980 463712
rect 150032 463700 150038 463752
rect 244090 463700 244096 463752
rect 244148 463740 244154 463752
rect 251174 463740 251180 463752
rect 244148 463712 251180 463740
rect 244148 463700 244154 463712
rect 251174 463700 251180 463712
rect 251232 463700 251238 463752
rect 111794 462408 111800 462460
rect 111852 462448 111858 462460
rect 119890 462448 119896 462460
rect 111852 462420 119896 462448
rect 111852 462408 111858 462420
rect 119890 462408 119896 462420
rect 119948 462408 119954 462460
rect 111886 462340 111892 462392
rect 111944 462380 111950 462392
rect 153010 462380 153016 462392
rect 111944 462352 153016 462380
rect 111944 462340 111950 462352
rect 153010 462340 153016 462352
rect 153068 462340 153074 462392
rect 243998 462340 244004 462392
rect 244056 462380 244062 462392
rect 251174 462380 251180 462392
rect 244056 462352 251180 462380
rect 244056 462340 244062 462352
rect 251174 462340 251180 462352
rect 251232 462340 251238 462392
rect 111794 460980 111800 461032
rect 111852 461020 111858 461032
rect 137738 461020 137744 461032
rect 111852 460992 137744 461020
rect 111852 460980 111858 460992
rect 137738 460980 137744 460992
rect 137796 460980 137802 461032
rect 111886 460912 111892 460964
rect 111944 460952 111950 460964
rect 144730 460952 144736 460964
rect 111944 460924 144736 460952
rect 111944 460912 111950 460924
rect 144730 460912 144736 460924
rect 144788 460912 144794 460964
rect 237006 460164 237012 460216
rect 237064 460204 237070 460216
rect 252094 460204 252100 460216
rect 237064 460176 252100 460204
rect 237064 460164 237070 460176
rect 252094 460164 252100 460176
rect 252152 460164 252158 460216
rect 111794 459552 111800 459604
rect 111852 459592 111858 459604
rect 150066 459592 150072 459604
rect 111852 459564 150072 459592
rect 111852 459552 111858 459564
rect 150066 459552 150072 459564
rect 150124 459552 150130 459604
rect 226058 459552 226064 459604
rect 226116 459592 226122 459604
rect 251174 459592 251180 459604
rect 226116 459564 251180 459592
rect 226116 459552 226122 459564
rect 251174 459552 251180 459564
rect 251232 459552 251238 459604
rect 111794 458260 111800 458312
rect 111852 458300 111858 458312
rect 130930 458300 130936 458312
rect 111852 458272 130936 458300
rect 111852 458260 111858 458272
rect 130930 458260 130936 458272
rect 130988 458260 130994 458312
rect 111886 458192 111892 458244
rect 111944 458232 111950 458244
rect 133598 458232 133604 458244
rect 111944 458204 133604 458232
rect 111944 458192 111950 458204
rect 133598 458192 133604 458204
rect 133656 458192 133662 458244
rect 248046 458192 248052 458244
rect 248104 458232 248110 458244
rect 251174 458232 251180 458244
rect 248104 458204 251180 458232
rect 248104 458192 248110 458204
rect 251174 458192 251180 458204
rect 251232 458192 251238 458244
rect 111794 456764 111800 456816
rect 111852 456804 111858 456816
rect 132310 456804 132316 456816
rect 111852 456776 132316 456804
rect 111852 456764 111858 456776
rect 132310 456764 132316 456776
rect 132368 456764 132374 456816
rect 238478 456764 238484 456816
rect 238536 456804 238542 456816
rect 251174 456804 251180 456816
rect 238536 456776 251180 456804
rect 238536 456764 238542 456776
rect 251174 456764 251180 456776
rect 251232 456764 251238 456816
rect 573358 456764 573364 456816
rect 573416 456804 573422 456816
rect 580166 456804 580172 456816
rect 573416 456776 580172 456804
rect 573416 456764 573422 456776
rect 580166 456764 580172 456776
rect 580224 456764 580230 456816
rect 111886 455472 111892 455524
rect 111944 455512 111950 455524
rect 132402 455512 132408 455524
rect 111944 455484 132408 455512
rect 111944 455472 111950 455484
rect 132402 455472 132408 455484
rect 132460 455472 132466 455524
rect 111794 455404 111800 455456
rect 111852 455444 111858 455456
rect 139210 455444 139216 455456
rect 111852 455416 139216 455444
rect 111852 455404 111858 455416
rect 139210 455404 139216 455416
rect 139268 455404 139274 455456
rect 239858 455404 239864 455456
rect 239916 455444 239922 455456
rect 251174 455444 251180 455456
rect 239916 455416 251180 455444
rect 239916 455404 239922 455416
rect 251174 455404 251180 455416
rect 251232 455404 251238 455456
rect 111794 454520 111800 454572
rect 111852 454560 111858 454572
rect 115014 454560 115020 454572
rect 111852 454532 115020 454560
rect 111852 454520 111858 454532
rect 115014 454520 115020 454532
rect 115072 454520 115078 454572
rect 111794 454044 111800 454096
rect 111852 454084 111858 454096
rect 142062 454084 142068 454096
rect 111852 454056 142068 454084
rect 111852 454044 111858 454056
rect 142062 454044 142068 454056
rect 142120 454044 142126 454096
rect 223390 454044 223396 454096
rect 223448 454084 223454 454096
rect 251174 454084 251180 454096
rect 223448 454056 251180 454084
rect 223448 454044 223454 454056
rect 251174 454044 251180 454056
rect 251232 454044 251238 454096
rect 111794 452684 111800 452736
rect 111852 452724 111858 452736
rect 116394 452724 116400 452736
rect 111852 452696 116400 452724
rect 111852 452684 111858 452696
rect 116394 452684 116400 452696
rect 116452 452684 116458 452736
rect 111886 452616 111892 452668
rect 111944 452656 111950 452668
rect 122742 452656 122748 452668
rect 111944 452628 122748 452656
rect 111944 452616 111950 452628
rect 122742 452616 122748 452628
rect 122800 452616 122806 452668
rect 111886 451324 111892 451376
rect 111944 451364 111950 451376
rect 124122 451364 124128 451376
rect 111944 451336 124128 451364
rect 111944 451324 111950 451336
rect 124122 451324 124128 451336
rect 124180 451324 124186 451376
rect 111794 451256 111800 451308
rect 111852 451296 111858 451308
rect 148870 451296 148876 451308
rect 111852 451268 148876 451296
rect 111852 451256 111858 451268
rect 148870 451256 148876 451268
rect 148928 451256 148934 451308
rect 241238 451256 241244 451308
rect 241296 451296 241302 451308
rect 251174 451296 251180 451308
rect 241296 451268 251180 451296
rect 241296 451256 241302 451268
rect 251174 451256 251180 451268
rect 251232 451256 251238 451308
rect 119614 450508 119620 450560
rect 119672 450548 119678 450560
rect 155678 450548 155684 450560
rect 119672 450520 155684 450548
rect 119672 450508 119678 450520
rect 155678 450508 155684 450520
rect 155736 450508 155742 450560
rect 111794 449964 111800 450016
rect 111852 450004 111858 450016
rect 119246 450004 119252 450016
rect 111852 449976 119252 450004
rect 111852 449964 111858 449976
rect 119246 449964 119252 449976
rect 119304 449964 119310 450016
rect 111886 449896 111892 449948
rect 111944 449936 111950 449948
rect 119982 449936 119988 449948
rect 111944 449908 119988 449936
rect 111944 449896 111950 449908
rect 119982 449896 119988 449908
rect 120040 449896 120046 449948
rect 226886 449896 226892 449948
rect 226944 449936 226950 449948
rect 251174 449936 251180 449948
rect 226944 449908 251180 449936
rect 226944 449896 226950 449908
rect 251174 449896 251180 449908
rect 251232 449896 251238 449948
rect 111794 448604 111800 448656
rect 111852 448644 111858 448656
rect 116486 448644 116492 448656
rect 111852 448616 116492 448644
rect 111852 448604 111858 448616
rect 116486 448604 116492 448616
rect 116544 448604 116550 448656
rect 111886 448536 111892 448588
rect 111944 448576 111950 448588
rect 145926 448576 145932 448588
rect 111944 448548 145932 448576
rect 111944 448536 111950 448548
rect 145926 448536 145932 448548
rect 145984 448536 145990 448588
rect 223482 448536 223488 448588
rect 223540 448576 223546 448588
rect 251174 448576 251180 448588
rect 223540 448548 251180 448576
rect 223540 448536 223546 448548
rect 251174 448536 251180 448548
rect 251232 448536 251238 448588
rect 111794 447108 111800 447160
rect 111852 447148 111858 447160
rect 140682 447148 140688 447160
rect 111852 447120 140688 447148
rect 111852 447108 111858 447120
rect 140682 447108 140688 447120
rect 140740 447108 140746 447160
rect 231578 447108 231584 447160
rect 231636 447148 231642 447160
rect 251174 447148 251180 447160
rect 231636 447120 251180 447148
rect 231636 447108 231642 447120
rect 251174 447108 251180 447120
rect 251232 447108 251238 447160
rect 251726 446428 251732 446480
rect 251784 446468 251790 446480
rect 252278 446468 252284 446480
rect 251784 446440 252284 446468
rect 251784 446428 251790 446440
rect 252278 446428 252284 446440
rect 252336 446428 252342 446480
rect 251726 446292 251732 446344
rect 251784 446332 251790 446344
rect 252462 446332 252468 446344
rect 251784 446304 252468 446332
rect 251784 446292 251790 446304
rect 252462 446292 252468 446304
rect 252520 446292 252526 446344
rect 226794 445748 226800 445800
rect 226852 445788 226858 445800
rect 251174 445788 251180 445800
rect 226852 445760 251180 445788
rect 226852 445748 226858 445760
rect 251174 445748 251180 445760
rect 251232 445748 251238 445800
rect 242526 444388 242532 444440
rect 242584 444428 242590 444440
rect 251174 444428 251180 444440
rect 242584 444400 251180 444428
rect 242584 444388 242590 444400
rect 251174 444388 251180 444400
rect 251232 444388 251238 444440
rect 231670 441600 231676 441652
rect 231728 441640 231734 441652
rect 251174 441640 251180 441652
rect 231728 441612 251180 441640
rect 231728 441600 231734 441612
rect 251174 441600 251180 441612
rect 251232 441600 251238 441652
rect 228634 440240 228640 440292
rect 228692 440280 228698 440292
rect 251174 440280 251180 440292
rect 228692 440252 251180 440280
rect 228692 440240 228698 440252
rect 251174 440240 251180 440252
rect 251232 440240 251238 440292
rect 230290 439492 230296 439544
rect 230348 439532 230354 439544
rect 251726 439532 251732 439544
rect 230348 439504 251732 439532
rect 230348 439492 230354 439504
rect 251726 439492 251732 439504
rect 251784 439492 251790 439544
rect 222010 438880 222016 438932
rect 222068 438920 222074 438932
rect 251174 438920 251180 438932
rect 222068 438892 251180 438920
rect 222068 438880 222074 438892
rect 251174 438880 251180 438892
rect 251232 438880 251238 438932
rect 246206 437452 246212 437504
rect 246264 437492 246270 437504
rect 251174 437492 251180 437504
rect 246264 437464 251180 437492
rect 246264 437452 246270 437464
rect 251174 437452 251180 437464
rect 251232 437452 251238 437504
rect 246942 436160 246948 436212
rect 247000 436200 247006 436212
rect 251174 436200 251180 436212
rect 247000 436172 251180 436200
rect 247000 436160 247006 436172
rect 251174 436160 251180 436172
rect 251232 436160 251238 436212
rect 231762 436092 231768 436144
rect 231820 436132 231826 436144
rect 251266 436132 251272 436144
rect 231820 436104 251272 436132
rect 231820 436092 231826 436104
rect 251266 436092 251272 436104
rect 251324 436092 251330 436144
rect 226150 434732 226156 434784
rect 226208 434772 226214 434784
rect 251174 434772 251180 434784
rect 226208 434744 251180 434772
rect 226208 434732 226214 434744
rect 251174 434732 251180 434744
rect 251232 434732 251238 434784
rect 238570 433304 238576 433356
rect 238628 433344 238634 433356
rect 251174 433344 251180 433356
rect 238628 433316 251180 433344
rect 238628 433304 238634 433316
rect 251174 433304 251180 433316
rect 251232 433304 251238 433356
rect 224126 431944 224132 431996
rect 224184 431984 224190 431996
rect 251174 431984 251180 431996
rect 224184 431956 251180 431984
rect 224184 431944 224190 431956
rect 251174 431944 251180 431956
rect 251232 431944 251238 431996
rect 228726 430584 228732 430636
rect 228784 430624 228790 430636
rect 251174 430624 251180 430636
rect 228784 430596 251180 430624
rect 228784 430584 228790 430596
rect 251174 430584 251180 430596
rect 251232 430584 251238 430636
rect 158438 429836 158444 429888
rect 158496 429876 158502 429888
rect 169754 429876 169760 429888
rect 158496 429848 169760 429876
rect 158496 429836 158502 429848
rect 169754 429836 169760 429848
rect 169812 429836 169818 429888
rect 245378 429156 245384 429208
rect 245436 429196 245442 429208
rect 251174 429196 251180 429208
rect 245436 429168 251180 429196
rect 245436 429156 245442 429168
rect 251174 429156 251180 429168
rect 251232 429156 251238 429208
rect 239950 427796 239956 427848
rect 240008 427836 240014 427848
rect 251174 427836 251180 427848
rect 240008 427808 251180 427836
rect 240008 427796 240014 427808
rect 251174 427796 251180 427808
rect 251232 427796 251238 427848
rect 245470 426504 245476 426556
rect 245528 426544 245534 426556
rect 251266 426544 251272 426556
rect 245528 426516 251272 426544
rect 245528 426504 245534 426516
rect 251266 426504 251272 426516
rect 251324 426504 251330 426556
rect 228818 426436 228824 426488
rect 228876 426476 228882 426488
rect 251174 426476 251180 426488
rect 228876 426448 251180 426476
rect 228876 426436 228882 426448
rect 251174 426436 251180 426448
rect 251232 426436 251238 426488
rect 222746 425076 222752 425128
rect 222804 425116 222810 425128
rect 251174 425116 251180 425128
rect 222804 425088 251180 425116
rect 222804 425076 222810 425088
rect 251174 425076 251180 425088
rect 251232 425076 251238 425128
rect 248966 423648 248972 423700
rect 249024 423688 249030 423700
rect 251174 423688 251180 423700
rect 249024 423660 251180 423688
rect 249024 423648 249030 423660
rect 251174 423648 251180 423660
rect 251232 423648 251238 423700
rect 3326 422288 3332 422340
rect 3384 422328 3390 422340
rect 156598 422328 156604 422340
rect 3384 422300 156604 422328
rect 3384 422288 3390 422300
rect 156598 422288 156604 422300
rect 156656 422288 156662 422340
rect 228910 420928 228916 420980
rect 228968 420968 228974 420980
rect 251174 420968 251180 420980
rect 228968 420940 251180 420968
rect 228968 420928 228974 420940
rect 251174 420928 251180 420940
rect 251232 420928 251238 420980
rect 226242 419500 226248 419552
rect 226300 419540 226306 419552
rect 251174 419540 251180 419552
rect 226300 419512 251180 419540
rect 226300 419500 226306 419512
rect 251174 419500 251180 419512
rect 251232 419500 251238 419552
rect 242618 418140 242624 418192
rect 242676 418180 242682 418192
rect 251174 418180 251180 418192
rect 242676 418152 251180 418180
rect 242676 418140 242682 418152
rect 251174 418140 251180 418152
rect 251232 418140 251238 418192
rect 244182 416780 244188 416832
rect 244240 416820 244246 416832
rect 251174 416820 251180 416832
rect 244240 416792 251180 416820
rect 244240 416780 244246 416792
rect 251174 416780 251180 416792
rect 251232 416780 251238 416832
rect 229002 415488 229008 415540
rect 229060 415528 229066 415540
rect 251266 415528 251272 415540
rect 229060 415500 251272 415528
rect 229060 415488 229066 415500
rect 251266 415488 251272 415500
rect 251324 415488 251330 415540
rect 224034 415420 224040 415472
rect 224092 415460 224098 415472
rect 251174 415460 251180 415472
rect 224092 415432 251180 415460
rect 224092 415420 224098 415432
rect 251174 415420 251180 415432
rect 251232 415420 251238 415472
rect 245562 413992 245568 414044
rect 245620 414032 245626 414044
rect 251174 414032 251180 414044
rect 245620 414004 251180 414032
rect 245620 413992 245626 414004
rect 251174 413992 251180 414004
rect 251232 413992 251238 414044
rect 219710 413924 219716 413976
rect 219768 413964 219774 413976
rect 234246 413964 234252 413976
rect 219768 413936 234252 413964
rect 219768 413924 219774 413936
rect 234246 413924 234252 413936
rect 234304 413924 234310 413976
rect 219986 413856 219992 413908
rect 220044 413896 220050 413908
rect 233970 413896 233976 413908
rect 220044 413868 233976 413896
rect 220044 413856 220050 413868
rect 233970 413856 233976 413868
rect 234028 413856 234034 413908
rect 220722 413788 220728 413840
rect 220780 413828 220786 413840
rect 234154 413828 234160 413840
rect 220780 413800 234160 413828
rect 220780 413788 220786 413800
rect 234154 413788 234160 413800
rect 234212 413788 234218 413840
rect 219802 413720 219808 413772
rect 219860 413760 219866 413772
rect 231118 413760 231124 413772
rect 219860 413732 231124 413760
rect 219860 413720 219866 413732
rect 231118 413720 231124 413732
rect 231176 413720 231182 413772
rect 248138 412632 248144 412684
rect 248196 412672 248202 412684
rect 251174 412672 251180 412684
rect 248196 412644 251180 412672
rect 248196 412632 248202 412644
rect 251174 412632 251180 412644
rect 251232 412632 251238 412684
rect 220722 412564 220728 412616
rect 220780 412604 220786 412616
rect 239490 412604 239496 412616
rect 220780 412576 239496 412604
rect 220780 412564 220786 412576
rect 239490 412564 239496 412576
rect 239548 412564 239554 412616
rect 219894 412088 219900 412140
rect 219952 412128 219958 412140
rect 228358 412128 228364 412140
rect 219952 412100 228364 412128
rect 219952 412088 219958 412100
rect 228358 412088 228364 412100
rect 228416 412088 228422 412140
rect 220078 411884 220084 411936
rect 220136 411924 220142 411936
rect 224218 411924 224224 411936
rect 220136 411896 224224 411924
rect 220136 411884 220142 411896
rect 224218 411884 224224 411896
rect 224276 411884 224282 411936
rect 223942 411272 223948 411324
rect 224000 411312 224006 411324
rect 251174 411312 251180 411324
rect 224000 411284 251180 411312
rect 224000 411272 224006 411284
rect 251174 411272 251180 411284
rect 251232 411272 251238 411324
rect 220722 411204 220728 411256
rect 220780 411244 220786 411256
rect 250438 411244 250444 411256
rect 220780 411216 250444 411244
rect 220780 411204 220786 411216
rect 250438 411204 250444 411216
rect 250496 411204 250502 411256
rect 219802 411136 219808 411188
rect 219860 411176 219866 411188
rect 244918 411176 244924 411188
rect 219860 411148 244924 411176
rect 219860 411136 219866 411148
rect 244918 411136 244924 411148
rect 244976 411136 244982 411188
rect 220078 410932 220084 410984
rect 220136 410972 220142 410984
rect 225598 410972 225604 410984
rect 220136 410944 225604 410972
rect 220136 410932 220142 410944
rect 225598 410932 225604 410944
rect 225656 410932 225662 410984
rect 3326 409844 3332 409896
rect 3384 409884 3390 409896
rect 152458 409884 152464 409896
rect 3384 409856 152464 409884
rect 3384 409844 3390 409856
rect 152458 409844 152464 409856
rect 152516 409844 152522 409896
rect 233970 409844 233976 409896
rect 234028 409884 234034 409896
rect 251174 409884 251180 409896
rect 234028 409856 251180 409884
rect 234028 409844 234034 409856
rect 251174 409844 251180 409856
rect 251232 409844 251238 409896
rect 220078 409776 220084 409828
rect 220136 409816 220142 409828
rect 232590 409816 232596 409828
rect 220136 409788 232596 409816
rect 220136 409776 220142 409788
rect 232590 409776 232596 409788
rect 232648 409776 232654 409828
rect 220722 409708 220728 409760
rect 220780 409748 220786 409760
rect 228450 409748 228456 409760
rect 220780 409720 228456 409748
rect 220780 409708 220786 409720
rect 228450 409708 228456 409720
rect 228508 409708 228514 409760
rect 219894 409640 219900 409692
rect 219952 409680 219958 409692
rect 222838 409680 222844 409692
rect 219952 409652 222844 409680
rect 219952 409640 219958 409652
rect 222838 409640 222844 409652
rect 222896 409640 222902 409692
rect 123754 409096 123760 409148
rect 123812 409136 123818 409148
rect 154666 409136 154672 409148
rect 123812 409108 154672 409136
rect 123812 409096 123818 409108
rect 154666 409096 154672 409108
rect 154724 409096 154730 409148
rect 234154 408484 234160 408536
rect 234212 408524 234218 408536
rect 251174 408524 251180 408536
rect 234212 408496 251180 408524
rect 234212 408484 234218 408496
rect 251174 408484 251180 408496
rect 251232 408484 251238 408536
rect 140038 408416 140044 408468
rect 140096 408456 140102 408468
rect 154942 408456 154948 408468
rect 140096 408428 154948 408456
rect 140096 408416 140102 408428
rect 154942 408416 154948 408428
rect 155000 408416 155006 408468
rect 220078 408416 220084 408468
rect 220136 408456 220142 408468
rect 245010 408456 245016 408468
rect 220136 408428 245016 408456
rect 220136 408416 220142 408428
rect 245010 408416 245016 408428
rect 245068 408416 245074 408468
rect 219894 408348 219900 408400
rect 219952 408388 219958 408400
rect 231302 408388 231308 408400
rect 219952 408360 231308 408388
rect 219952 408348 219958 408360
rect 231302 408348 231308 408360
rect 231360 408348 231366 408400
rect 220722 408280 220728 408332
rect 220780 408320 220786 408332
rect 231210 408320 231216 408332
rect 220780 408292 231216 408320
rect 220780 408280 220786 408292
rect 231210 408280 231216 408292
rect 231268 408280 231274 408332
rect 117958 407736 117964 407788
rect 118016 407776 118022 407788
rect 155770 407776 155776 407788
rect 118016 407748 155776 407776
rect 118016 407736 118022 407748
rect 155770 407736 155776 407748
rect 155828 407736 155834 407788
rect 231026 407124 231032 407176
rect 231084 407164 231090 407176
rect 251174 407164 251180 407176
rect 231084 407136 251180 407164
rect 231084 407124 231090 407136
rect 251174 407124 251180 407136
rect 251232 407124 251238 407176
rect 123570 407056 123576 407108
rect 123628 407096 123634 407108
rect 154850 407096 154856 407108
rect 123628 407068 154856 407096
rect 123628 407056 123634 407068
rect 154850 407056 154856 407068
rect 154908 407056 154914 407108
rect 220078 407056 220084 407108
rect 220136 407096 220142 407108
rect 242158 407096 242164 407108
rect 220136 407068 242164 407096
rect 220136 407056 220142 407068
rect 242158 407056 242164 407068
rect 242216 407056 242222 407108
rect 123662 406988 123668 407040
rect 123720 407028 123726 407040
rect 154758 407028 154764 407040
rect 123720 407000 154764 407028
rect 123720 406988 123726 407000
rect 154758 406988 154764 407000
rect 154816 406988 154822 407040
rect 220722 406988 220728 407040
rect 220780 407028 220786 407040
rect 236638 407028 236644 407040
rect 220780 407000 236644 407028
rect 220780 406988 220786 407000
rect 236638 406988 236644 407000
rect 236696 406988 236702 407040
rect 123478 406920 123484 406972
rect 123536 406960 123542 406972
rect 154942 406960 154948 406972
rect 123536 406932 154948 406960
rect 123536 406920 123542 406932
rect 154942 406920 154948 406932
rect 155000 406920 155006 406972
rect 142890 406852 142896 406904
rect 142948 406892 142954 406904
rect 154574 406892 154580 406904
rect 142948 406864 154580 406892
rect 142948 406852 142954 406864
rect 154574 406852 154580 406864
rect 154632 406852 154638 406904
rect 220722 406648 220728 406700
rect 220780 406688 220786 406700
rect 228542 406688 228548 406700
rect 220780 406660 228548 406688
rect 220780 406648 220786 406660
rect 228542 406648 228548 406660
rect 228600 406648 228606 406700
rect 219894 406376 219900 406428
rect 219952 406416 219958 406428
rect 222930 406416 222936 406428
rect 219952 406388 222936 406416
rect 219952 406376 219958 406388
rect 222930 406376 222936 406388
rect 222988 406376 222994 406428
rect 113818 405628 113824 405680
rect 113876 405668 113882 405680
rect 154758 405668 154764 405680
rect 113876 405640 154764 405668
rect 113876 405628 113882 405640
rect 154758 405628 154764 405640
rect 154816 405628 154822 405680
rect 220078 405628 220084 405680
rect 220136 405668 220142 405680
rect 221642 405668 221648 405680
rect 220136 405640 221648 405668
rect 220136 405628 220142 405640
rect 221642 405628 221648 405640
rect 221700 405628 221706 405680
rect 113910 405560 113916 405612
rect 113968 405600 113974 405612
rect 154850 405600 154856 405612
rect 113968 405572 154856 405600
rect 113968 405560 113974 405572
rect 154850 405560 154856 405572
rect 154908 405560 154914 405612
rect 155034 405560 155040 405612
rect 155092 405600 155098 405612
rect 155310 405600 155316 405612
rect 155092 405572 155316 405600
rect 155092 405560 155098 405572
rect 155310 405560 155316 405572
rect 155368 405560 155374 405612
rect 120718 405492 120724 405544
rect 120776 405532 120782 405544
rect 154942 405532 154948 405544
rect 120776 405504 154948 405532
rect 120776 405492 120782 405504
rect 154942 405492 154948 405504
rect 155000 405492 155006 405544
rect 123846 405424 123852 405476
rect 123904 405464 123910 405476
rect 154574 405464 154580 405476
rect 123904 405436 154580 405464
rect 123904 405424 123910 405436
rect 154574 405424 154580 405436
rect 154632 405424 154638 405476
rect 220722 405356 220728 405408
rect 220780 405396 220786 405408
rect 226978 405396 226984 405408
rect 220780 405368 226984 405396
rect 220780 405356 220786 405368
rect 226978 405356 226984 405368
rect 227036 405356 227042 405408
rect 219894 405288 219900 405340
rect 219952 405328 219958 405340
rect 224310 405328 224316 405340
rect 219952 405300 224316 405328
rect 219952 405288 219958 405300
rect 224310 405288 224316 405300
rect 224368 405288 224374 405340
rect 222102 404336 222108 404388
rect 222160 404376 222166 404388
rect 251174 404376 251180 404388
rect 222160 404348 251180 404376
rect 222160 404336 222166 404348
rect 251174 404336 251180 404348
rect 251232 404336 251238 404388
rect 115198 404268 115204 404320
rect 115256 404308 115262 404320
rect 154666 404308 154672 404320
rect 115256 404280 154672 404308
rect 115256 404268 115262 404280
rect 154666 404268 154672 404280
rect 154724 404268 154730 404320
rect 219986 404268 219992 404320
rect 220044 404308 220050 404320
rect 246574 404308 246580 404320
rect 220044 404280 246580 404308
rect 220044 404268 220050 404280
rect 246574 404268 246580 404280
rect 246632 404268 246638 404320
rect 122098 404200 122104 404252
rect 122156 404240 122162 404252
rect 154942 404240 154948 404252
rect 122156 404212 154948 404240
rect 122156 404200 122162 404212
rect 154942 404200 154948 404212
rect 155000 404200 155006 404252
rect 220722 404200 220728 404252
rect 220780 404240 220786 404252
rect 239582 404240 239588 404252
rect 220780 404212 239588 404240
rect 220780 404200 220786 404212
rect 239582 404200 239588 404212
rect 239640 404200 239646 404252
rect 122190 404132 122196 404184
rect 122248 404172 122254 404184
rect 154850 404172 154856 404184
rect 122248 404144 154856 404172
rect 122248 404132 122254 404144
rect 154850 404132 154856 404144
rect 154908 404132 154914 404184
rect 220078 404132 220084 404184
rect 220136 404172 220142 404184
rect 235258 404172 235264 404184
rect 220136 404144 235264 404172
rect 220136 404132 220142 404144
rect 235258 404132 235264 404144
rect 235316 404132 235322 404184
rect 138750 404064 138756 404116
rect 138808 404104 138814 404116
rect 154758 404104 154764 404116
rect 138808 404076 154764 404104
rect 138808 404064 138814 404076
rect 154758 404064 154764 404076
rect 154816 404064 154822 404116
rect 219710 402908 219716 402960
rect 219768 402948 219774 402960
rect 238110 402948 238116 402960
rect 219768 402920 238116 402948
rect 219768 402908 219774 402920
rect 238110 402908 238116 402920
rect 238168 402908 238174 402960
rect 130378 402840 130384 402892
rect 130436 402880 130442 402892
rect 154758 402880 154764 402892
rect 130436 402852 154764 402880
rect 130436 402840 130442 402852
rect 154758 402840 154764 402852
rect 154816 402840 154822 402892
rect 220170 402840 220176 402892
rect 220228 402880 220234 402892
rect 229830 402880 229836 402892
rect 220228 402852 229836 402880
rect 220228 402840 220234 402852
rect 229830 402840 229836 402852
rect 229888 402840 229894 402892
rect 133138 402772 133144 402824
rect 133196 402812 133202 402824
rect 154850 402812 154856 402824
rect 133196 402784 154856 402812
rect 133196 402772 133202 402784
rect 154850 402772 154856 402784
rect 154908 402772 154914 402824
rect 220722 402772 220728 402824
rect 220780 402812 220786 402824
rect 229738 402812 229744 402824
rect 220780 402784 229744 402812
rect 220780 402772 220786 402784
rect 229738 402772 229744 402784
rect 229796 402772 229802 402824
rect 134518 402704 134524 402756
rect 134576 402744 134582 402756
rect 154666 402744 154672 402756
rect 134576 402716 154672 402744
rect 134576 402704 134582 402716
rect 154666 402704 154672 402716
rect 154724 402704 154730 402756
rect 219802 402704 219808 402756
rect 219860 402744 219866 402756
rect 221734 402744 221740 402756
rect 219860 402716 221740 402744
rect 219860 402704 219866 402716
rect 221734 402704 221740 402716
rect 221792 402704 221798 402756
rect 122374 402636 122380 402688
rect 122432 402676 122438 402688
rect 154942 402676 154948 402688
rect 122432 402648 154948 402676
rect 122432 402636 122438 402648
rect 154942 402636 154948 402648
rect 155000 402636 155006 402688
rect 152550 402432 152556 402484
rect 152608 402472 152614 402484
rect 155218 402472 155224 402484
rect 152608 402444 155224 402472
rect 152608 402432 152614 402444
rect 155218 402432 155224 402444
rect 155276 402432 155282 402484
rect 231210 401616 231216 401668
rect 231268 401656 231274 401668
rect 251174 401656 251180 401668
rect 231268 401628 251180 401656
rect 231268 401616 231274 401628
rect 251174 401616 251180 401628
rect 251232 401616 251238 401668
rect 152642 401548 152648 401600
rect 152700 401588 152706 401600
rect 155218 401588 155224 401600
rect 152700 401560 155224 401588
rect 152700 401548 152706 401560
rect 155218 401548 155224 401560
rect 155276 401548 155282 401600
rect 220722 401548 220728 401600
rect 220780 401588 220786 401600
rect 250530 401588 250536 401600
rect 220780 401560 250536 401588
rect 220780 401548 220786 401560
rect 250530 401548 250536 401560
rect 250588 401548 250594 401600
rect 141510 401480 141516 401532
rect 141568 401520 141574 401532
rect 154850 401520 154856 401532
rect 141568 401492 154856 401520
rect 141568 401480 141574 401492
rect 154850 401480 154856 401492
rect 154908 401480 154914 401532
rect 220170 401480 220176 401532
rect 220228 401520 220234 401532
rect 238202 401520 238208 401532
rect 220228 401492 238208 401520
rect 220228 401480 220234 401492
rect 238202 401480 238208 401492
rect 238260 401480 238266 401532
rect 142982 401412 142988 401464
rect 143040 401452 143046 401464
rect 155034 401452 155040 401464
rect 143040 401424 155040 401452
rect 143040 401412 143046 401424
rect 155034 401412 155040 401424
rect 155092 401412 155098 401464
rect 114002 401344 114008 401396
rect 114060 401384 114066 401396
rect 154942 401384 154948 401396
rect 114060 401356 154948 401384
rect 114060 401344 114066 401356
rect 154942 401344 154948 401356
rect 155000 401344 155006 401396
rect 220078 401276 220084 401328
rect 220136 401316 220142 401328
rect 221826 401316 221832 401328
rect 220136 401288 221832 401316
rect 220136 401276 220142 401288
rect 221826 401276 221832 401288
rect 221884 401276 221890 401328
rect 122282 400868 122288 400920
rect 122340 400908 122346 400920
rect 155126 400908 155132 400920
rect 122340 400880 155132 400908
rect 122340 400868 122346 400880
rect 155126 400868 155132 400880
rect 155184 400868 155190 400920
rect 229738 400868 229744 400920
rect 229796 400908 229802 400920
rect 251634 400908 251640 400920
rect 229796 400880 251640 400908
rect 229796 400868 229802 400880
rect 251634 400868 251640 400880
rect 251692 400868 251698 400920
rect 251542 400800 251548 400852
rect 251600 400840 251606 400852
rect 251910 400840 251916 400852
rect 251600 400812 251916 400840
rect 251600 400800 251606 400812
rect 251910 400800 251916 400812
rect 251968 400800 251974 400852
rect 127618 400120 127624 400172
rect 127676 400160 127682 400172
rect 154758 400160 154764 400172
rect 127676 400132 154764 400160
rect 127676 400120 127682 400132
rect 154758 400120 154764 400132
rect 154816 400120 154822 400172
rect 220722 400120 220728 400172
rect 220780 400160 220786 400172
rect 251542 400160 251548 400172
rect 220780 400132 251548 400160
rect 220780 400120 220786 400132
rect 251542 400120 251548 400132
rect 251600 400120 251606 400172
rect 130470 400052 130476 400104
rect 130528 400092 130534 400104
rect 155034 400092 155040 400104
rect 130528 400064 155040 400092
rect 130528 400052 130534 400064
rect 155034 400052 155040 400064
rect 155092 400052 155098 400104
rect 220078 400052 220084 400104
rect 220136 400092 220142 400104
rect 249150 400092 249156 400104
rect 220136 400064 249156 400092
rect 220136 400052 220142 400064
rect 249150 400052 249156 400064
rect 249208 400052 249214 400104
rect 133230 399984 133236 400036
rect 133288 400024 133294 400036
rect 154850 400024 154856 400036
rect 133288 399996 154856 400024
rect 133288 399984 133294 399996
rect 154850 399984 154856 399996
rect 154908 399984 154914 400036
rect 220170 399984 220176 400036
rect 220228 400024 220234 400036
rect 235350 400024 235356 400036
rect 220228 399996 235356 400024
rect 220228 399984 220234 399996
rect 235350 399984 235356 399996
rect 235408 399984 235414 400036
rect 134610 399916 134616 399968
rect 134668 399956 134674 399968
rect 154942 399956 154948 399968
rect 134668 399928 154948 399956
rect 134668 399916 134674 399928
rect 154942 399916 154948 399928
rect 155000 399916 155006 399968
rect 219986 399916 219992 399968
rect 220044 399956 220050 399968
rect 227070 399956 227076 399968
rect 220044 399928 227076 399956
rect 220044 399916 220050 399928
rect 227070 399916 227076 399928
rect 227128 399916 227134 399968
rect 226978 398828 226984 398880
rect 227036 398868 227042 398880
rect 251174 398868 251180 398880
rect 227036 398840 251180 398868
rect 227036 398828 227042 398840
rect 251174 398828 251180 398840
rect 251232 398828 251238 398880
rect 152734 398760 152740 398812
rect 152792 398800 152798 398812
rect 154574 398800 154580 398812
rect 152792 398772 154580 398800
rect 152792 398760 152798 398772
rect 154574 398760 154580 398772
rect 154632 398760 154638 398812
rect 220078 398760 220084 398812
rect 220136 398800 220142 398812
rect 247770 398800 247776 398812
rect 220136 398772 247776 398800
rect 220136 398760 220142 398772
rect 247770 398760 247776 398772
rect 247828 398760 247834 398812
rect 141602 398692 141608 398744
rect 141660 398732 141666 398744
rect 154666 398732 154672 398744
rect 141660 398704 154672 398732
rect 141660 398692 141666 398704
rect 154666 398692 154672 398704
rect 154724 398692 154730 398744
rect 220170 398692 220176 398744
rect 220228 398732 220234 398744
rect 237006 398732 237012 398744
rect 220228 398704 237012 398732
rect 220228 398692 220234 398704
rect 237006 398692 237012 398704
rect 237064 398692 237070 398744
rect 144270 398624 144276 398676
rect 144328 398664 144334 398676
rect 154850 398664 154856 398676
rect 144328 398636 154856 398664
rect 144328 398624 144334 398636
rect 154850 398624 154856 398636
rect 154908 398624 154914 398676
rect 220722 398624 220728 398676
rect 220780 398664 220786 398676
rect 232682 398664 232688 398676
rect 220780 398636 232688 398664
rect 220780 398624 220786 398636
rect 232682 398624 232688 398636
rect 232740 398624 232746 398676
rect 149790 398556 149796 398608
rect 149848 398596 149854 398608
rect 155034 398596 155040 398608
rect 149848 398568 155040 398596
rect 149848 398556 149854 398568
rect 155034 398556 155040 398568
rect 155092 398556 155098 398608
rect 137278 398488 137284 398540
rect 137336 398528 137342 398540
rect 154942 398528 154948 398540
rect 137336 398500 154948 398528
rect 137336 398488 137342 398500
rect 154942 398488 154948 398500
rect 155000 398488 155006 398540
rect 127710 398080 127716 398132
rect 127768 398120 127774 398132
rect 154758 398120 154764 398132
rect 127768 398092 154764 398120
rect 127768 398080 127774 398092
rect 154758 398080 154764 398092
rect 154816 398080 154822 398132
rect 251726 398080 251732 398132
rect 251784 398120 251790 398132
rect 252462 398120 252468 398132
rect 251784 398092 252468 398120
rect 251784 398080 251790 398092
rect 252462 398080 252468 398092
rect 252520 398080 252526 398132
rect 3326 397468 3332 397520
rect 3384 397508 3390 397520
rect 134518 397508 134524 397520
rect 3384 397480 134524 397508
rect 3384 397468 3390 397480
rect 134518 397468 134524 397480
rect 134576 397468 134582 397520
rect 222838 397468 222844 397520
rect 222896 397508 222902 397520
rect 251174 397508 251180 397520
rect 222896 397480 251180 397508
rect 222896 397468 222902 397480
rect 251174 397468 251180 397480
rect 251232 397468 251238 397520
rect 116578 397400 116584 397452
rect 116636 397440 116642 397452
rect 155034 397440 155040 397452
rect 116636 397412 155040 397440
rect 116636 397400 116642 397412
rect 155034 397400 155040 397412
rect 155092 397400 155098 397452
rect 220722 397400 220728 397452
rect 220780 397440 220786 397452
rect 247862 397440 247868 397452
rect 220780 397412 247868 397440
rect 220780 397400 220786 397412
rect 247862 397400 247868 397412
rect 247920 397400 247926 397452
rect 122650 397332 122656 397384
rect 122708 397372 122714 397384
rect 155126 397372 155132 397384
rect 122708 397344 155132 397372
rect 122708 397332 122714 397344
rect 155126 397332 155132 397344
rect 155184 397332 155190 397384
rect 220170 397332 220176 397384
rect 220228 397372 220234 397384
rect 243722 397372 243728 397384
rect 220228 397344 243728 397372
rect 220228 397332 220234 397344
rect 243722 397332 243728 397344
rect 243780 397332 243786 397384
rect 130562 397264 130568 397316
rect 130620 397304 130626 397316
rect 154850 397304 154856 397316
rect 130620 397276 154856 397304
rect 130620 397264 130626 397276
rect 154850 397264 154856 397276
rect 154908 397264 154914 397316
rect 134702 397196 134708 397248
rect 134760 397236 134766 397248
rect 154942 397236 154948 397248
rect 134760 397208 154948 397236
rect 134760 397196 134766 397208
rect 154942 397196 154948 397208
rect 155000 397196 155006 397248
rect 220722 396856 220728 396908
rect 220780 396896 220786 396908
rect 223022 396896 223028 396908
rect 220780 396868 223028 396896
rect 220780 396856 220786 396868
rect 223022 396856 223028 396868
rect 223080 396856 223086 396908
rect 247770 396040 247776 396092
rect 247828 396080 247834 396092
rect 251174 396080 251180 396092
rect 247828 396052 251180 396080
rect 247828 396040 247834 396052
rect 251174 396040 251180 396052
rect 251232 396040 251238 396092
rect 112438 395972 112444 396024
rect 112496 396012 112502 396024
rect 154758 396012 154764 396024
rect 112496 395984 154764 396012
rect 112496 395972 112502 395984
rect 154758 395972 154764 395984
rect 154816 395972 154822 396024
rect 155218 395972 155224 396024
rect 155276 396012 155282 396024
rect 155494 396012 155500 396024
rect 155276 395984 155500 396012
rect 155276 395972 155282 395984
rect 155494 395972 155500 395984
rect 155552 395972 155558 396024
rect 220078 395972 220084 396024
rect 220136 396012 220142 396024
rect 246666 396012 246672 396024
rect 220136 395984 246672 396012
rect 220136 395972 220142 395984
rect 246666 395972 246672 395984
rect 246724 395972 246730 396024
rect 115290 395904 115296 395956
rect 115348 395944 115354 395956
rect 154850 395944 154856 395956
rect 115348 395916 154856 395944
rect 115348 395904 115354 395916
rect 154850 395904 154856 395916
rect 154908 395904 154914 395956
rect 220170 395904 220176 395956
rect 220228 395944 220234 395956
rect 241054 395944 241060 395956
rect 220228 395916 241060 395944
rect 220228 395904 220234 395916
rect 241054 395904 241060 395916
rect 241112 395904 241118 395956
rect 140130 395836 140136 395888
rect 140188 395876 140194 395888
rect 154942 395876 154948 395888
rect 140188 395848 154948 395876
rect 140188 395836 140194 395848
rect 154942 395836 154948 395848
rect 155000 395836 155006 395888
rect 220722 395836 220728 395888
rect 220780 395876 220786 395888
rect 229922 395876 229928 395888
rect 220780 395848 229928 395876
rect 220780 395836 220786 395848
rect 229922 395836 229928 395848
rect 229980 395836 229986 395888
rect 140222 395768 140228 395820
rect 140280 395808 140286 395820
rect 155034 395808 155040 395820
rect 140280 395780 155040 395808
rect 140280 395768 140286 395780
rect 155034 395768 155040 395780
rect 155092 395768 155098 395820
rect 148410 395700 148416 395752
rect 148468 395740 148474 395752
rect 154666 395740 154672 395752
rect 148468 395712 154672 395740
rect 148468 395700 148474 395712
rect 154666 395700 154672 395712
rect 154724 395700 154730 395752
rect 127802 395292 127808 395344
rect 127860 395332 127866 395344
rect 154942 395332 154948 395344
rect 127860 395304 154948 395332
rect 127860 395292 127866 395304
rect 154942 395292 154948 395304
rect 155000 395292 155006 395344
rect 221734 394680 221740 394732
rect 221792 394720 221798 394732
rect 251174 394720 251180 394732
rect 221792 394692 251180 394720
rect 221792 394680 221798 394692
rect 251174 394680 251180 394692
rect 251232 394680 251238 394732
rect 115382 394612 115388 394664
rect 115440 394652 115446 394664
rect 154574 394652 154580 394664
rect 115440 394624 154580 394652
rect 115440 394612 115446 394624
rect 154574 394612 154580 394624
rect 154632 394612 154638 394664
rect 220722 394612 220728 394664
rect 220780 394652 220786 394664
rect 250622 394652 250628 394664
rect 220780 394624 250628 394652
rect 220780 394612 220786 394624
rect 250622 394612 250628 394624
rect 250680 394612 250686 394664
rect 118050 394544 118056 394596
rect 118108 394584 118114 394596
rect 154666 394584 154672 394596
rect 118108 394556 154672 394584
rect 118108 394544 118114 394556
rect 154666 394544 154672 394556
rect 154724 394544 154730 394596
rect 219986 394544 219992 394596
rect 220044 394584 220050 394596
rect 245102 394584 245108 394596
rect 220044 394556 245108 394584
rect 220044 394544 220050 394556
rect 245102 394544 245108 394556
rect 245160 394544 245166 394596
rect 130654 394476 130660 394528
rect 130712 394516 130718 394528
rect 154758 394516 154764 394528
rect 130712 394488 154764 394516
rect 130712 394476 130718 394488
rect 154758 394476 154764 394488
rect 154816 394476 154822 394528
rect 220170 394476 220176 394528
rect 220228 394516 220234 394528
rect 232774 394516 232780 394528
rect 220228 394488 232780 394516
rect 220228 394476 220234 394488
rect 232774 394476 232780 394488
rect 232832 394476 232838 394528
rect 147030 394408 147036 394460
rect 147088 394448 147094 394460
rect 154850 394448 154856 394460
rect 147088 394420 154856 394448
rect 147088 394408 147094 394420
rect 154850 394408 154856 394420
rect 154908 394408 154914 394460
rect 128998 393932 129004 393984
rect 129056 393972 129062 393984
rect 155126 393972 155132 393984
rect 129056 393944 155132 393972
rect 129056 393932 129062 393944
rect 155126 393932 155132 393944
rect 155184 393932 155190 393984
rect 250438 393864 250444 393916
rect 250496 393904 250502 393916
rect 251910 393904 251916 393916
rect 250496 393876 251916 393904
rect 250496 393864 250502 393876
rect 251910 393864 251916 393876
rect 251968 393864 251974 393916
rect 221642 393320 221648 393372
rect 221700 393360 221706 393372
rect 251174 393360 251180 393372
rect 221700 393332 251180 393360
rect 221700 393320 221706 393332
rect 251174 393320 251180 393332
rect 251232 393320 251238 393372
rect 151170 393252 151176 393304
rect 151228 393292 151234 393304
rect 155034 393292 155040 393304
rect 151228 393264 155040 393292
rect 151228 393252 151234 393264
rect 155034 393252 155040 393264
rect 155092 393252 155098 393304
rect 220170 393252 220176 393304
rect 220228 393292 220234 393304
rect 242250 393292 242256 393304
rect 220228 393264 242256 393292
rect 220228 393252 220234 393264
rect 242250 393252 242256 393264
rect 242308 393252 242314 393304
rect 119338 393184 119344 393236
rect 119396 393224 119402 393236
rect 154942 393224 154948 393236
rect 119396 393196 154948 393224
rect 119396 393184 119402 393196
rect 154942 393184 154948 393196
rect 155000 393184 155006 393236
rect 220722 393184 220728 393236
rect 220780 393224 220786 393236
rect 230014 393224 230020 393236
rect 220780 393196 230020 393224
rect 220780 393184 220786 393196
rect 230014 393184 230020 393196
rect 230072 393184 230078 393236
rect 138842 393116 138848 393168
rect 138900 393156 138906 393168
rect 154758 393156 154764 393168
rect 138900 393128 154764 393156
rect 138900 393116 138906 393128
rect 154758 393116 154764 393128
rect 154816 393116 154822 393168
rect 143074 393048 143080 393100
rect 143132 393088 143138 393100
rect 154850 393088 154856 393100
rect 143132 393060 154856 393088
rect 143132 393048 143138 393060
rect 154850 393048 154856 393060
rect 154908 393048 154914 393100
rect 115474 392980 115480 393032
rect 115532 393020 115538 393032
rect 154942 393020 154948 393032
rect 115532 392992 154948 393020
rect 115532 392980 115538 392992
rect 154942 392980 154948 392992
rect 155000 392980 155006 393032
rect 220170 391960 220176 392012
rect 220228 392000 220234 392012
rect 220446 392000 220452 392012
rect 220228 391972 220452 392000
rect 220228 391960 220234 391972
rect 220446 391960 220452 391972
rect 220504 391960 220510 392012
rect 236638 391960 236644 392012
rect 236696 392000 236702 392012
rect 251174 392000 251180 392012
rect 236696 391972 251180 392000
rect 236696 391960 236702 391972
rect 251174 391960 251180 391972
rect 251232 391960 251238 392012
rect 220262 391892 220268 391944
rect 220320 391932 220326 391944
rect 249426 391932 249432 391944
rect 220320 391904 249432 391932
rect 220320 391892 220326 391904
rect 249426 391892 249432 391904
rect 249484 391892 249490 391944
rect 126238 391824 126244 391876
rect 126296 391864 126302 391876
rect 154942 391864 154948 391876
rect 126296 391836 154948 391864
rect 126296 391824 126302 391836
rect 154942 391824 154948 391836
rect 155000 391824 155006 391876
rect 220722 391824 220728 391876
rect 220780 391864 220786 391876
rect 249334 391864 249340 391876
rect 220780 391836 249340 391864
rect 220780 391824 220786 391836
rect 249334 391824 249340 391836
rect 249392 391824 249398 391876
rect 130746 391756 130752 391808
rect 130804 391796 130810 391808
rect 154758 391796 154764 391808
rect 130804 391768 154764 391796
rect 130804 391756 130810 391768
rect 154758 391756 154764 391768
rect 154816 391756 154822 391808
rect 220446 391756 220452 391808
rect 220504 391796 220510 391808
rect 239674 391796 239680 391808
rect 220504 391768 239680 391796
rect 220504 391756 220510 391768
rect 239674 391756 239680 391768
rect 239732 391756 239738 391808
rect 149698 391688 149704 391740
rect 149756 391728 149762 391740
rect 154666 391728 154672 391740
rect 149756 391700 154672 391728
rect 149756 391688 149762 391700
rect 154666 391688 154672 391700
rect 154724 391688 154730 391740
rect 116670 391620 116676 391672
rect 116728 391660 116734 391672
rect 154942 391660 154948 391672
rect 116728 391632 154948 391660
rect 116728 391620 116734 391632
rect 154942 391620 154948 391632
rect 155000 391620 155006 391672
rect 220722 391484 220728 391536
rect 220780 391524 220786 391536
rect 227162 391524 227168 391536
rect 220780 391496 227168 391524
rect 220780 391484 220786 391496
rect 227162 391484 227168 391496
rect 227220 391484 227226 391536
rect 219986 390532 219992 390584
rect 220044 390572 220050 390584
rect 251174 390572 251180 390584
rect 220044 390544 251180 390572
rect 220044 390532 220050 390544
rect 251174 390532 251180 390544
rect 251232 390532 251238 390584
rect 152826 390464 152832 390516
rect 152884 390504 152890 390516
rect 154574 390504 154580 390516
rect 152884 390476 154580 390504
rect 152884 390464 152890 390476
rect 154574 390464 154580 390476
rect 154632 390464 154638 390516
rect 220722 390464 220728 390516
rect 220780 390504 220786 390516
rect 231394 390504 231400 390516
rect 220780 390476 231400 390504
rect 220780 390464 220786 390476
rect 231394 390464 231400 390476
rect 231452 390464 231458 390516
rect 118142 390396 118148 390448
rect 118200 390436 118206 390448
rect 155034 390436 155040 390448
rect 118200 390408 155040 390436
rect 118200 390396 118206 390408
rect 155034 390396 155040 390408
rect 155092 390396 155098 390448
rect 119430 390328 119436 390380
rect 119488 390368 119494 390380
rect 154942 390368 154948 390380
rect 119488 390340 154948 390368
rect 119488 390328 119494 390340
rect 154942 390328 154948 390340
rect 155000 390328 155006 390380
rect 219894 390328 219900 390380
rect 219952 390368 219958 390380
rect 227254 390368 227260 390380
rect 219952 390340 227260 390368
rect 219952 390328 219958 390340
rect 227254 390328 227260 390340
rect 227312 390328 227318 390380
rect 145742 390260 145748 390312
rect 145800 390300 145806 390312
rect 154850 390300 154856 390312
rect 145800 390272 154856 390300
rect 145800 390260 145806 390272
rect 154850 390260 154856 390272
rect 154908 390260 154914 390312
rect 115566 390192 115572 390244
rect 115624 390232 115630 390244
rect 154942 390232 154948 390244
rect 115624 390204 154948 390232
rect 115624 390192 115630 390204
rect 154942 390192 154948 390204
rect 155000 390192 155006 390244
rect 119522 389784 119528 389836
rect 119580 389824 119586 389836
rect 155218 389824 155224 389836
rect 119580 389796 155224 389824
rect 119580 389784 119586 389796
rect 155218 389784 155224 389796
rect 155276 389784 155282 389836
rect 219894 389172 219900 389224
rect 219952 389212 219958 389224
rect 251174 389212 251180 389224
rect 219952 389184 251180 389212
rect 219952 389172 219958 389184
rect 251174 389172 251180 389184
rect 251232 389172 251238 389224
rect 116854 389104 116860 389156
rect 116912 389144 116918 389156
rect 154850 389144 154856 389156
rect 116912 389116 154856 389144
rect 116912 389104 116918 389116
rect 154850 389104 154856 389116
rect 154908 389104 154914 389156
rect 220722 389104 220728 389156
rect 220780 389144 220786 389156
rect 238294 389144 238300 389156
rect 220780 389116 238300 389144
rect 220780 389104 220786 389116
rect 238294 389104 238300 389116
rect 238352 389104 238358 389156
rect 130838 389036 130844 389088
rect 130896 389076 130902 389088
rect 154758 389076 154764 389088
rect 130896 389048 154764 389076
rect 130896 389036 130902 389048
rect 154758 389036 154764 389048
rect 154816 389036 154822 389088
rect 220446 389036 220452 389088
rect 220504 389076 220510 389088
rect 234338 389076 234344 389088
rect 220504 389048 234344 389076
rect 220504 389036 220510 389048
rect 234338 389036 234344 389048
rect 234396 389036 234402 389088
rect 131758 388968 131764 389020
rect 131816 389008 131822 389020
rect 154666 389008 154672 389020
rect 131816 388980 154672 389008
rect 131816 388968 131822 388980
rect 154666 388968 154672 388980
rect 154724 388968 154730 389020
rect 220078 388968 220084 389020
rect 220136 389008 220142 389020
rect 225690 389008 225696 389020
rect 220136 388980 225696 389008
rect 220136 388968 220142 388980
rect 225690 388968 225696 388980
rect 225748 388968 225754 389020
rect 144362 388900 144368 388952
rect 144420 388940 144426 388952
rect 154942 388940 154948 388952
rect 144420 388912 154948 388940
rect 144420 388900 144426 388912
rect 154942 388900 154948 388912
rect 155000 388900 155006 388952
rect 251634 388424 251640 388476
rect 251692 388464 251698 388476
rect 251910 388464 251916 388476
rect 251692 388436 251916 388464
rect 251692 388424 251698 388436
rect 251910 388424 251916 388436
rect 251968 388424 251974 388476
rect 249150 387812 249156 387864
rect 249208 387852 249214 387864
rect 251450 387852 251456 387864
rect 249208 387824 251456 387852
rect 249208 387812 249214 387824
rect 251450 387812 251456 387824
rect 251508 387812 251514 387864
rect 151262 387744 151268 387796
rect 151320 387784 151326 387796
rect 155126 387784 155132 387796
rect 151320 387756 155132 387784
rect 151320 387744 151326 387756
rect 155126 387744 155132 387756
rect 155184 387744 155190 387796
rect 220446 387744 220452 387796
rect 220504 387784 220510 387796
rect 242342 387784 242348 387796
rect 220504 387756 242348 387784
rect 220504 387744 220510 387756
rect 242342 387744 242348 387756
rect 242400 387744 242406 387796
rect 116762 387676 116768 387728
rect 116820 387716 116826 387728
rect 154942 387716 154948 387728
rect 116820 387688 154948 387716
rect 116820 387676 116826 387688
rect 154942 387676 154948 387688
rect 155000 387676 155006 387728
rect 220722 387676 220728 387728
rect 220780 387716 220786 387728
rect 236730 387716 236736 387728
rect 220780 387688 236736 387716
rect 220780 387676 220786 387688
rect 236730 387676 236736 387688
rect 236788 387676 236794 387728
rect 137370 387608 137376 387660
rect 137428 387648 137434 387660
rect 154758 387648 154764 387660
rect 137428 387620 154764 387648
rect 137428 387608 137434 387620
rect 154758 387608 154764 387620
rect 154816 387608 154822 387660
rect 220262 387608 220268 387660
rect 220320 387648 220326 387660
rect 234430 387648 234436 387660
rect 220320 387620 234436 387648
rect 220320 387608 220326 387620
rect 234430 387608 234436 387620
rect 234488 387608 234494 387660
rect 145558 387540 145564 387592
rect 145616 387580 145622 387592
rect 154850 387580 154856 387592
rect 145616 387552 154856 387580
rect 145616 387540 145622 387552
rect 154850 387540 154856 387552
rect 154908 387540 154914 387592
rect 112530 387472 112536 387524
rect 112588 387512 112594 387524
rect 155034 387512 155040 387524
rect 112588 387484 155040 387512
rect 112588 387472 112594 387484
rect 155034 387472 155040 387484
rect 155092 387472 155098 387524
rect 147214 387064 147220 387116
rect 147272 387104 147278 387116
rect 155494 387104 155500 387116
rect 147272 387076 155500 387104
rect 147272 387064 147278 387076
rect 155494 387064 155500 387076
rect 155552 387064 155558 387116
rect 151354 386316 151360 386368
rect 151412 386356 151418 386368
rect 155034 386356 155040 386368
rect 151412 386328 155040 386356
rect 151412 386316 151418 386328
rect 155034 386316 155040 386328
rect 155092 386316 155098 386368
rect 220722 386316 220728 386368
rect 220780 386356 220786 386368
rect 243814 386356 243820 386368
rect 220780 386328 243820 386356
rect 220780 386316 220786 386328
rect 243814 386316 243820 386328
rect 243872 386316 243878 386368
rect 131850 386248 131856 386300
rect 131908 386288 131914 386300
rect 154666 386288 154672 386300
rect 131908 386260 154672 386288
rect 131908 386248 131914 386260
rect 154666 386248 154672 386260
rect 154724 386248 154730 386300
rect 220170 386248 220176 386300
rect 220228 386288 220234 386300
rect 236822 386288 236828 386300
rect 220228 386260 236828 386288
rect 220228 386248 220234 386260
rect 236822 386248 236828 386260
rect 236880 386248 236886 386300
rect 148502 386180 148508 386232
rect 148560 386220 148566 386232
rect 154850 386220 154856 386232
rect 148560 386192 154856 386220
rect 148560 386180 148566 386192
rect 154850 386180 154856 386192
rect 154908 386180 154914 386232
rect 220446 386180 220452 386232
rect 220504 386220 220510 386232
rect 234522 386220 234528 386232
rect 220504 386192 234528 386220
rect 220504 386180 220510 386192
rect 234522 386180 234528 386192
rect 234580 386180 234586 386232
rect 127894 386112 127900 386164
rect 127952 386152 127958 386164
rect 154942 386152 154948 386164
rect 127952 386124 154948 386152
rect 127952 386112 127958 386124
rect 154942 386112 154948 386124
rect 155000 386112 155006 386164
rect 126790 385636 126796 385688
rect 126848 385676 126854 385688
rect 155218 385676 155224 385688
rect 126848 385648 155224 385676
rect 126848 385636 126854 385648
rect 155218 385636 155224 385648
rect 155276 385636 155282 385688
rect 112622 384956 112628 385008
rect 112680 384996 112686 385008
rect 155126 384996 155132 385008
rect 112680 384968 155132 384996
rect 112680 384956 112686 384968
rect 155126 384956 155132 384968
rect 155184 384956 155190 385008
rect 220262 384956 220268 385008
rect 220320 384996 220326 385008
rect 246758 384996 246764 385008
rect 220320 384968 246764 384996
rect 220320 384956 220326 384968
rect 246758 384956 246764 384968
rect 246816 384956 246822 385008
rect 116946 384888 116952 384940
rect 117004 384928 117010 384940
rect 155034 384928 155040 384940
rect 117004 384900 155040 384928
rect 117004 384888 117010 384900
rect 155034 384888 155040 384900
rect 155092 384888 155098 384940
rect 220722 384888 220728 384940
rect 220780 384928 220786 384940
rect 245194 384928 245200 384940
rect 220780 384900 245200 384928
rect 220780 384888 220786 384900
rect 245194 384888 245200 384900
rect 245252 384888 245258 384940
rect 143166 384820 143172 384872
rect 143224 384860 143230 384872
rect 154942 384860 154948 384872
rect 143224 384832 154948 384860
rect 143224 384820 143230 384832
rect 154942 384820 154948 384832
rect 155000 384820 155006 384872
rect 220446 384820 220452 384872
rect 220504 384860 220510 384872
rect 236914 384860 236920 384872
rect 220504 384832 236920 384860
rect 220504 384820 220510 384832
rect 236914 384820 236920 384832
rect 236972 384820 236978 384872
rect 147122 384752 147128 384804
rect 147180 384792 147186 384804
rect 154850 384792 154856 384804
rect 147180 384764 154856 384792
rect 147180 384752 147186 384764
rect 154850 384752 154856 384764
rect 154908 384752 154914 384804
rect 220354 384752 220360 384804
rect 220412 384792 220418 384804
rect 223114 384792 223120 384804
rect 220412 384764 223120 384792
rect 220412 384752 220418 384764
rect 223114 384752 223120 384764
rect 223172 384752 223178 384804
rect 148594 384684 148600 384736
rect 148652 384724 148658 384736
rect 154666 384724 154672 384736
rect 148652 384696 154672 384724
rect 148652 384684 148658 384696
rect 154666 384684 154672 384696
rect 154724 384684 154730 384736
rect 227070 383664 227076 383716
rect 227128 383704 227134 383716
rect 251174 383704 251180 383716
rect 227128 383676 251180 383704
rect 227128 383664 227134 383676
rect 251174 383664 251180 383676
rect 251232 383664 251238 383716
rect 220078 383596 220084 383648
rect 220136 383636 220142 383648
rect 232866 383636 232872 383648
rect 220136 383608 232872 383636
rect 220136 383596 220142 383608
rect 232866 383596 232872 383608
rect 232924 383596 232930 383648
rect 131942 383528 131948 383580
rect 132000 383568 132006 383580
rect 154850 383568 154856 383580
rect 132000 383540 154856 383568
rect 132000 383528 132006 383540
rect 154850 383528 154856 383540
rect 154908 383528 154914 383580
rect 138934 383460 138940 383512
rect 138992 383500 138998 383512
rect 154942 383500 154948 383512
rect 138992 383472 154948 383500
rect 138992 383460 138998 383472
rect 154942 383460 154948 383472
rect 155000 383460 155006 383512
rect 149882 383392 149888 383444
rect 149940 383432 149946 383444
rect 154666 383432 154672 383444
rect 149940 383404 154672 383432
rect 149940 383392 149946 383404
rect 154666 383392 154672 383404
rect 154724 383392 154730 383444
rect 124858 383324 124864 383376
rect 124916 383364 124922 383376
rect 154942 383364 154948 383376
rect 124916 383336 154948 383364
rect 124916 383324 124922 383336
rect 154942 383324 154948 383336
rect 155000 383324 155006 383376
rect 220446 383256 220452 383308
rect 220504 383296 220510 383308
rect 221918 383296 221924 383308
rect 220504 383268 221924 383296
rect 220504 383256 220510 383268
rect 221918 383256 221924 383268
rect 221976 383256 221982 383308
rect 234246 382236 234252 382288
rect 234304 382276 234310 382288
rect 251174 382276 251180 382288
rect 234304 382248 251180 382276
rect 234304 382236 234310 382248
rect 251174 382236 251180 382248
rect 251232 382236 251238 382288
rect 114094 382168 114100 382220
rect 114152 382208 114158 382220
rect 154942 382208 154948 382220
rect 114152 382180 154948 382208
rect 114152 382168 114158 382180
rect 154942 382168 154948 382180
rect 155000 382168 155006 382220
rect 220722 382168 220728 382220
rect 220780 382208 220786 382220
rect 247954 382208 247960 382220
rect 220780 382180 247960 382208
rect 220780 382168 220786 382180
rect 247954 382168 247960 382180
rect 248012 382168 248018 382220
rect 117038 382100 117044 382152
rect 117096 382140 117102 382152
rect 154574 382140 154580 382152
rect 117096 382112 154580 382140
rect 117096 382100 117102 382112
rect 154574 382100 154580 382112
rect 154632 382100 154638 382152
rect 220630 382100 220636 382152
rect 220688 382140 220694 382152
rect 235442 382140 235448 382152
rect 220688 382112 235448 382140
rect 220688 382100 220694 382112
rect 235442 382100 235448 382112
rect 235500 382100 235506 382152
rect 139026 382032 139032 382084
rect 139084 382072 139090 382084
rect 154850 382072 154856 382084
rect 139084 382044 154856 382072
rect 139084 382032 139090 382044
rect 154850 382032 154856 382044
rect 154908 382032 154914 382084
rect 220538 382032 220544 382084
rect 220596 382072 220602 382084
rect 232958 382072 232964 382084
rect 220596 382044 232964 382072
rect 220596 382032 220602 382044
rect 232958 382032 232964 382044
rect 233016 382032 233022 382084
rect 144454 381964 144460 382016
rect 144512 382004 144518 382016
rect 154942 382004 154948 382016
rect 144512 381976 154948 382004
rect 144512 381964 144518 381976
rect 154942 381964 154948 381976
rect 155000 381964 155006 382016
rect 112714 380808 112720 380860
rect 112772 380848 112778 380860
rect 154942 380848 154948 380860
rect 112772 380820 154948 380848
rect 112772 380808 112778 380820
rect 154942 380808 154948 380820
rect 155000 380808 155006 380860
rect 220630 380808 220636 380860
rect 220688 380848 220694 380860
rect 250714 380848 250720 380860
rect 220688 380820 250720 380848
rect 220688 380808 220694 380820
rect 250714 380808 250720 380820
rect 250772 380808 250778 380860
rect 118234 380740 118240 380792
rect 118292 380780 118298 380792
rect 154758 380780 154764 380792
rect 118292 380752 154764 380780
rect 118292 380740 118298 380752
rect 154758 380740 154764 380752
rect 154816 380740 154822 380792
rect 220722 380740 220728 380792
rect 220780 380780 220786 380792
rect 231486 380780 231492 380792
rect 220780 380752 231492 380780
rect 220780 380740 220786 380752
rect 231486 380740 231492 380752
rect 231544 380740 231550 380792
rect 126330 380672 126336 380724
rect 126388 380712 126394 380724
rect 155034 380712 155040 380724
rect 126388 380684 155040 380712
rect 126388 380672 126394 380684
rect 155034 380672 155040 380684
rect 155092 380672 155098 380724
rect 219710 380672 219716 380724
rect 219768 380712 219774 380724
rect 227438 380712 227444 380724
rect 219768 380684 227444 380712
rect 219768 380672 219774 380684
rect 227438 380672 227444 380684
rect 227496 380672 227502 380724
rect 132034 380604 132040 380656
rect 132092 380644 132098 380656
rect 154850 380644 154856 380656
rect 132092 380616 154856 380644
rect 132092 380604 132098 380616
rect 154850 380604 154856 380616
rect 154908 380604 154914 380656
rect 143258 380536 143264 380588
rect 143316 380576 143322 380588
rect 154942 380576 154948 380588
rect 143316 380548 154948 380576
rect 143316 380536 143322 380548
rect 154942 380536 154948 380548
rect 155000 380536 155006 380588
rect 220722 380468 220728 380520
rect 220780 380508 220786 380520
rect 227346 380508 227352 380520
rect 220780 380480 227352 380508
rect 220780 380468 220786 380480
rect 227346 380468 227352 380480
rect 227404 380468 227410 380520
rect 220722 379448 220728 379500
rect 220780 379488 220786 379500
rect 249518 379488 249524 379500
rect 220780 379460 249524 379488
rect 220780 379448 220786 379460
rect 249518 379448 249524 379460
rect 249576 379448 249582 379500
rect 120810 379380 120816 379432
rect 120868 379420 120874 379432
rect 154850 379420 154856 379432
rect 120868 379392 154856 379420
rect 120868 379380 120874 379392
rect 154850 379380 154856 379392
rect 154908 379380 154914 379432
rect 220630 379380 220636 379432
rect 220688 379420 220694 379432
rect 235810 379420 235816 379432
rect 220688 379392 235816 379420
rect 220688 379380 220694 379392
rect 235810 379380 235816 379392
rect 235868 379380 235874 379432
rect 124950 379312 124956 379364
rect 125008 379352 125014 379364
rect 154942 379352 154948 379364
rect 125008 379324 154948 379352
rect 125008 379312 125014 379324
rect 154942 379312 154948 379324
rect 155000 379312 155006 379364
rect 220538 379312 220544 379364
rect 220596 379352 220602 379364
rect 235534 379352 235540 379364
rect 220596 379324 235540 379352
rect 220596 379312 220602 379324
rect 235534 379312 235540 379324
rect 235592 379312 235598 379364
rect 147306 379244 147312 379296
rect 147364 379284 147370 379296
rect 155034 379284 155040 379296
rect 147364 379256 155040 379284
rect 147364 379244 147370 379256
rect 155034 379244 155040 379256
rect 155092 379244 155098 379296
rect 118326 379176 118332 379228
rect 118384 379216 118390 379228
rect 154942 379216 154948 379228
rect 118384 379188 154948 379216
rect 118384 379176 118390 379188
rect 154942 379176 154948 379188
rect 155000 379176 155006 379228
rect 139118 378768 139124 378820
rect 139176 378808 139182 378820
rect 154666 378808 154672 378820
rect 139176 378780 154672 378808
rect 139176 378768 139182 378780
rect 154666 378768 154672 378780
rect 154724 378768 154730 378820
rect 220078 378156 220084 378208
rect 220136 378196 220142 378208
rect 579798 378196 579804 378208
rect 220136 378168 579804 378196
rect 220136 378156 220142 378168
rect 579798 378156 579804 378168
rect 579856 378156 579862 378208
rect 112806 378088 112812 378140
rect 112864 378128 112870 378140
rect 154942 378128 154948 378140
rect 112864 378100 154948 378128
rect 112864 378088 112870 378100
rect 154942 378088 154948 378100
rect 155000 378088 155006 378140
rect 220630 378088 220636 378140
rect 220688 378128 220694 378140
rect 235718 378128 235724 378140
rect 220688 378100 235724 378128
rect 220688 378088 220694 378100
rect 235718 378088 235724 378100
rect 235776 378088 235782 378140
rect 119706 378020 119712 378072
rect 119764 378060 119770 378072
rect 155034 378060 155040 378072
rect 119764 378032 155040 378060
rect 119764 378020 119770 378032
rect 155034 378020 155040 378032
rect 155092 378020 155098 378072
rect 220722 378020 220728 378072
rect 220780 378060 220786 378072
rect 235626 378060 235632 378072
rect 220780 378032 235632 378060
rect 220780 378020 220786 378032
rect 235626 378020 235632 378032
rect 235684 378020 235690 378072
rect 120902 377952 120908 378004
rect 120960 377992 120966 378004
rect 154758 377992 154764 378004
rect 120960 377964 154764 377992
rect 120960 377952 120966 377964
rect 154758 377952 154764 377964
rect 154816 377952 154822 378004
rect 220538 377952 220544 378004
rect 220596 377992 220602 378004
rect 233050 377992 233056 378004
rect 220596 377964 233056 377992
rect 220596 377952 220602 377964
rect 233050 377952 233056 377964
rect 233108 377952 233114 378004
rect 140314 377884 140320 377936
rect 140372 377924 140378 377936
rect 154850 377924 154856 377936
rect 140372 377896 154856 377924
rect 140372 377884 140378 377896
rect 154850 377884 154856 377896
rect 154908 377884 154914 377936
rect 144546 377816 144552 377868
rect 144604 377856 144610 377868
rect 154942 377856 154948 377868
rect 144604 377828 154948 377856
rect 144604 377816 144610 377828
rect 154942 377816 154948 377828
rect 155000 377816 155006 377868
rect 114186 376660 114192 376712
rect 114244 376700 114250 376712
rect 154942 376700 154948 376712
rect 114244 376672 154948 376700
rect 114244 376660 114250 376672
rect 154942 376660 154948 376672
rect 155000 376660 155006 376712
rect 220722 376660 220728 376712
rect 220780 376700 220786 376712
rect 252002 376700 252008 376712
rect 220780 376672 252008 376700
rect 220780 376660 220786 376672
rect 252002 376660 252008 376672
rect 252060 376660 252066 376712
rect 120994 376592 121000 376644
rect 121052 376632 121058 376644
rect 155034 376632 155040 376644
rect 121052 376604 155040 376632
rect 121052 376592 121058 376604
rect 155034 376592 155040 376604
rect 155092 376592 155098 376644
rect 219986 376592 219992 376644
rect 220044 376632 220050 376644
rect 225782 376632 225788 376644
rect 220044 376604 225788 376632
rect 220044 376592 220050 376604
rect 225782 376592 225788 376604
rect 225840 376592 225846 376644
rect 125042 376524 125048 376576
rect 125100 376564 125106 376576
rect 154850 376564 154856 376576
rect 125100 376536 154856 376564
rect 125100 376524 125106 376536
rect 154850 376524 154856 376536
rect 154908 376524 154914 376576
rect 145650 376456 145656 376508
rect 145708 376496 145714 376508
rect 154942 376496 154948 376508
rect 145708 376468 154948 376496
rect 145708 376456 145714 376468
rect 154942 376456 154948 376468
rect 155000 376456 155006 376508
rect 143350 375980 143356 376032
rect 143408 376020 143414 376032
rect 155126 376020 155132 376032
rect 143408 375992 155132 376020
rect 143408 375980 143414 375992
rect 155126 375980 155132 375992
rect 155184 375980 155190 376032
rect 219894 375980 219900 376032
rect 219952 376020 219958 376032
rect 241146 376020 241152 376032
rect 219952 375992 241152 376020
rect 219952 375980 219958 375992
rect 241146 375980 241152 375992
rect 241204 375980 241210 376032
rect 219986 375844 219992 375896
rect 220044 375884 220050 375896
rect 225874 375884 225880 375896
rect 220044 375856 225880 375884
rect 220044 375844 220050 375856
rect 225874 375844 225880 375856
rect 225932 375844 225938 375896
rect 154574 375408 154580 375420
rect 154040 375380 154580 375408
rect 112898 375300 112904 375352
rect 112956 375340 112962 375352
rect 154040 375340 154068 375380
rect 154574 375368 154580 375380
rect 154632 375368 154638 375420
rect 112956 375312 154068 375340
rect 112956 375300 112962 375312
rect 154114 375300 154120 375352
rect 154172 375340 154178 375352
rect 155034 375340 155040 375352
rect 154172 375312 155040 375340
rect 154172 375300 154178 375312
rect 155034 375300 155040 375312
rect 155092 375300 155098 375352
rect 220630 375300 220636 375352
rect 220688 375340 220694 375352
rect 250806 375340 250812 375352
rect 220688 375312 250812 375340
rect 220688 375300 220694 375312
rect 250806 375300 250812 375312
rect 250864 375300 250870 375352
rect 117130 375232 117136 375284
rect 117188 375272 117194 375284
rect 154942 375272 154948 375284
rect 117188 375244 154948 375272
rect 117188 375232 117194 375244
rect 154942 375232 154948 375244
rect 155000 375232 155006 375284
rect 220722 375232 220728 375284
rect 220780 375272 220786 375284
rect 243906 375272 243912 375284
rect 220780 375244 243912 375272
rect 220780 375232 220786 375244
rect 243906 375232 243912 375244
rect 243964 375232 243970 375284
rect 141694 375164 141700 375216
rect 141752 375204 141758 375216
rect 154850 375204 154856 375216
rect 141752 375176 154856 375204
rect 141752 375164 141758 375176
rect 154850 375164 154856 375176
rect 154908 375164 154914 375216
rect 219434 374824 219440 374876
rect 219492 374864 219498 374876
rect 225966 374864 225972 374876
rect 219492 374836 225972 374864
rect 219492 374824 219498 374836
rect 225966 374824 225972 374836
rect 226024 374824 226030 374876
rect 118418 374620 118424 374672
rect 118476 374660 118482 374672
rect 155586 374660 155592 374672
rect 118476 374632 155592 374660
rect 118476 374620 118482 374632
rect 155586 374620 155592 374632
rect 155644 374620 155650 374672
rect 125226 373940 125232 373992
rect 125284 373980 125290 373992
rect 154666 373980 154672 373992
rect 125284 373952 154672 373980
rect 125284 373940 125290 373952
rect 154666 373940 154672 373952
rect 154724 373940 154730 373992
rect 220722 373940 220728 373992
rect 220780 373980 220786 373992
rect 246850 373980 246856 373992
rect 220780 373952 246856 373980
rect 220780 373940 220786 373952
rect 246850 373940 246856 373952
rect 246908 373940 246914 373992
rect 126422 373872 126428 373924
rect 126480 373912 126486 373924
rect 154758 373912 154764 373924
rect 126480 373884 154764 373912
rect 126480 373872 126486 373884
rect 154758 373872 154764 373884
rect 154816 373872 154822 373924
rect 220630 373872 220636 373924
rect 220688 373912 220694 373924
rect 238386 373912 238392 373924
rect 220688 373884 238392 373912
rect 220688 373872 220694 373884
rect 238386 373872 238392 373884
rect 238444 373872 238450 373924
rect 129090 373804 129096 373856
rect 129148 373844 129154 373856
rect 154574 373844 154580 373856
rect 129148 373816 154580 373844
rect 129148 373804 129154 373816
rect 154574 373804 154580 373816
rect 154632 373804 154638 373856
rect 220538 373804 220544 373856
rect 220596 373844 220602 373856
rect 224402 373844 224408 373856
rect 220596 373816 224408 373844
rect 220596 373804 220602 373816
rect 224402 373804 224408 373816
rect 224460 373804 224466 373856
rect 141786 373736 141792 373788
rect 141844 373776 141850 373788
rect 154942 373776 154948 373788
rect 141844 373748 154948 373776
rect 141844 373736 141850 373748
rect 154942 373736 154948 373748
rect 155000 373736 155006 373788
rect 147398 373668 147404 373720
rect 147456 373708 147462 373720
rect 154850 373708 154856 373720
rect 147456 373680 154856 373708
rect 147456 373668 147462 373680
rect 154850 373668 154856 373680
rect 154908 373668 154914 373720
rect 114278 372512 114284 372564
rect 114336 372552 114342 372564
rect 154758 372552 154764 372564
rect 114336 372524 154764 372552
rect 114336 372512 114342 372524
rect 154758 372512 154764 372524
rect 154816 372512 154822 372564
rect 219986 372512 219992 372564
rect 220044 372552 220050 372564
rect 224770 372552 224776 372564
rect 220044 372524 224776 372552
rect 220044 372512 220050 372524
rect 224770 372512 224776 372524
rect 224828 372512 224834 372564
rect 121086 372444 121092 372496
rect 121144 372484 121150 372496
rect 154942 372484 154948 372496
rect 121144 372456 154948 372484
rect 121144 372444 121150 372456
rect 154942 372444 154948 372456
rect 155000 372444 155006 372496
rect 140406 372376 140412 372428
rect 140464 372416 140470 372428
rect 155126 372416 155132 372428
rect 140464 372388 155132 372416
rect 140464 372376 140470 372388
rect 155126 372376 155132 372388
rect 155184 372376 155190 372428
rect 140498 372308 140504 372360
rect 140556 372348 140562 372360
rect 154942 372348 154948 372360
rect 140556 372320 154948 372348
rect 140556 372308 140562 372320
rect 154942 372308 154948 372320
rect 155000 372308 155006 372360
rect 220354 372308 220360 372360
rect 220412 372348 220418 372360
rect 224494 372348 224500 372360
rect 220412 372320 224500 372348
rect 220412 372308 220418 372320
rect 224494 372308 224500 372320
rect 224552 372308 224558 372360
rect 148686 372240 148692 372292
rect 148744 372280 148750 372292
rect 154850 372280 154856 372292
rect 148744 372252 154856 372280
rect 148744 372240 148750 372252
rect 154850 372240 154856 372252
rect 154908 372240 154914 372292
rect 220446 371968 220452 372020
rect 220504 372008 220510 372020
rect 224586 372008 224592 372020
rect 220504 371980 224592 372008
rect 220504 371968 220510 371980
rect 224586 371968 224592 371980
rect 224644 371968 224650 372020
rect 218790 371832 218796 371884
rect 218848 371872 218854 371884
rect 580442 371872 580448 371884
rect 218848 371844 580448 371872
rect 218848 371832 218854 371844
rect 580442 371832 580448 371844
rect 580500 371832 580506 371884
rect 3326 371220 3332 371272
rect 3384 371260 3390 371272
rect 156690 371260 156696 371272
rect 3384 371232 156696 371260
rect 3384 371220 3390 371232
rect 156690 371220 156696 371232
rect 156748 371220 156754 371272
rect 115658 371152 115664 371204
rect 115716 371192 115722 371204
rect 154758 371192 154764 371204
rect 115716 371164 154764 371192
rect 115716 371152 115722 371164
rect 154758 371152 154764 371164
rect 154816 371152 154822 371204
rect 220538 371152 220544 371204
rect 220596 371192 220602 371204
rect 249610 371192 249616 371204
rect 220596 371164 249616 371192
rect 220596 371152 220602 371164
rect 249610 371152 249616 371164
rect 249668 371152 249674 371204
rect 127986 371084 127992 371136
rect 128044 371124 128050 371136
rect 154666 371124 154672 371136
rect 128044 371096 154672 371124
rect 128044 371084 128050 371096
rect 154666 371084 154672 371096
rect 154724 371084 154730 371136
rect 220722 371084 220728 371136
rect 220780 371124 220786 371136
rect 239766 371124 239772 371136
rect 220780 371096 239772 371124
rect 220780 371084 220786 371096
rect 239766 371084 239772 371096
rect 239824 371084 239830 371136
rect 133322 371016 133328 371068
rect 133380 371056 133386 371068
rect 154942 371056 154948 371068
rect 133380 371028 154948 371056
rect 133380 371016 133386 371028
rect 154942 371016 154948 371028
rect 155000 371016 155006 371068
rect 220630 371016 220636 371068
rect 220688 371056 220694 371068
rect 224678 371056 224684 371068
rect 220688 371028 224684 371056
rect 220688 371016 220694 371028
rect 224678 371016 224684 371028
rect 224736 371016 224742 371068
rect 135990 370948 135996 371000
rect 136048 370988 136054 371000
rect 154850 370988 154856 371000
rect 136048 370960 154856 370988
rect 136048 370948 136054 370960
rect 154850 370948 154856 370960
rect 154908 370948 154914 371000
rect 141878 370880 141884 370932
rect 141936 370920 141942 370932
rect 155126 370920 155132 370932
rect 141936 370892 155132 370920
rect 141936 370880 141942 370892
rect 155126 370880 155132 370892
rect 155184 370880 155190 370932
rect 219710 370472 219716 370524
rect 219768 370512 219774 370524
rect 242434 370512 242440 370524
rect 219768 370484 242440 370512
rect 219768 370472 219774 370484
rect 242434 370472 242440 370484
rect 242492 370472 242498 370524
rect 220538 370132 220544 370184
rect 220596 370172 220602 370184
rect 223298 370172 223304 370184
rect 220596 370144 223304 370172
rect 220596 370132 220602 370144
rect 223298 370132 223304 370144
rect 223356 370132 223362 370184
rect 114370 369792 114376 369844
rect 114428 369832 114434 369844
rect 154666 369832 154672 369844
rect 114428 369804 154672 369832
rect 114428 369792 114434 369804
rect 154666 369792 154672 369804
rect 154724 369792 154730 369844
rect 115750 369724 115756 369776
rect 115808 369764 115814 369776
rect 155126 369764 155132 369776
rect 115808 369736 155132 369764
rect 115808 369724 115814 369736
rect 155126 369724 155132 369736
rect 155184 369724 155190 369776
rect 119798 369656 119804 369708
rect 119856 369696 119862 369708
rect 154942 369696 154948 369708
rect 119856 369668 154948 369696
rect 119856 369656 119862 369668
rect 154942 369656 154948 369668
rect 155000 369656 155006 369708
rect 121178 369588 121184 369640
rect 121236 369628 121242 369640
rect 154850 369628 154856 369640
rect 121236 369600 154856 369628
rect 121236 369588 121242 369600
rect 154850 369588 154856 369600
rect 154908 369588 154914 369640
rect 220630 369588 220636 369640
rect 220688 369628 220694 369640
rect 223206 369628 223212 369640
rect 220688 369600 223212 369628
rect 220688 369588 220694 369600
rect 223206 369588 223212 369600
rect 223264 369588 223270 369640
rect 148778 369520 148784 369572
rect 148836 369560 148842 369572
rect 154758 369560 154764 369572
rect 148836 369532 154764 369560
rect 148836 369520 148842 369532
rect 154758 369520 154764 369532
rect 154816 369520 154822 369572
rect 220630 369316 220636 369368
rect 220688 369356 220694 369368
rect 227530 369356 227536 369368
rect 220688 369328 227536 369356
rect 220688 369316 220694 369328
rect 227530 369316 227536 369328
rect 227588 369316 227594 369368
rect 219986 369112 219992 369164
rect 220044 369152 220050 369164
rect 244090 369152 244096 369164
rect 220044 369124 244096 369152
rect 220044 369112 220050 369124
rect 244090 369112 244096 369124
rect 244148 369112 244154 369164
rect 151446 368432 151452 368484
rect 151504 368472 151510 368484
rect 154574 368472 154580 368484
rect 151504 368444 154580 368472
rect 151504 368432 151510 368444
rect 154574 368432 154580 368444
rect 154632 368432 154638 368484
rect 220538 368432 220544 368484
rect 220596 368472 220602 368484
rect 230106 368472 230112 368484
rect 220596 368444 230112 368472
rect 220596 368432 220602 368444
rect 230106 368432 230112 368444
rect 230164 368432 230170 368484
rect 129182 368364 129188 368416
rect 129240 368404 129246 368416
rect 154758 368404 154764 368416
rect 129240 368376 154764 368404
rect 129240 368364 129246 368376
rect 154758 368364 154764 368376
rect 154816 368364 154822 368416
rect 220722 368364 220728 368416
rect 220780 368404 220786 368416
rect 224862 368404 224868 368416
rect 220780 368376 224868 368404
rect 220780 368364 220786 368376
rect 224862 368364 224868 368376
rect 224920 368364 224926 368416
rect 140590 368296 140596 368348
rect 140648 368336 140654 368348
rect 154942 368336 154948 368348
rect 140648 368308 154948 368336
rect 140648 368296 140654 368308
rect 154942 368296 154948 368308
rect 155000 368296 155006 368348
rect 122466 368228 122472 368280
rect 122524 368268 122530 368280
rect 154850 368268 154856 368280
rect 122524 368240 154856 368268
rect 122524 368228 122530 368240
rect 154850 368228 154856 368240
rect 154908 368228 154914 368280
rect 219894 368024 219900 368076
rect 219952 368064 219958 368076
rect 227622 368064 227628 368076
rect 219952 368036 227628 368064
rect 219952 368024 219958 368036
rect 227622 368024 227628 368036
rect 227680 368024 227686 368076
rect 150066 367820 150072 367872
rect 150124 367860 150130 367872
rect 155310 367860 155316 367872
rect 150124 367832 155316 367860
rect 150124 367820 150130 367832
rect 155310 367820 155316 367832
rect 155368 367820 155374 367872
rect 118510 367752 118516 367804
rect 118568 367792 118574 367804
rect 155402 367792 155408 367804
rect 118568 367764 155408 367792
rect 118568 367752 118574 367764
rect 155402 367752 155408 367764
rect 155460 367752 155466 367804
rect 219618 367752 219624 367804
rect 219676 367792 219682 367804
rect 249702 367792 249708 367804
rect 219676 367764 249708 367792
rect 219676 367752 219682 367764
rect 249702 367752 249708 367764
rect 249760 367752 249766 367804
rect 126514 367004 126520 367056
rect 126572 367044 126578 367056
rect 155126 367044 155132 367056
rect 126572 367016 155132 367044
rect 126572 367004 126578 367016
rect 155126 367004 155132 367016
rect 155184 367004 155190 367056
rect 220538 367004 220544 367056
rect 220596 367044 220602 367056
rect 252186 367044 252192 367056
rect 220596 367016 252192 367044
rect 220596 367004 220602 367016
rect 252186 367004 252192 367016
rect 252244 367004 252250 367056
rect 128078 366936 128084 366988
rect 128136 366976 128142 366988
rect 154942 366976 154948 366988
rect 128136 366948 154948 366976
rect 128136 366936 128142 366948
rect 154942 366936 154948 366948
rect 155000 366936 155006 366988
rect 220722 366936 220728 366988
rect 220780 366976 220786 366988
rect 245286 366976 245292 366988
rect 220780 366948 245292 366976
rect 220780 366936 220786 366948
rect 245286 366936 245292 366948
rect 245344 366936 245350 366988
rect 137462 366868 137468 366920
rect 137520 366908 137526 366920
rect 154666 366908 154672 366920
rect 137520 366880 154672 366908
rect 137520 366868 137526 366880
rect 154666 366868 154672 366880
rect 154724 366868 154730 366920
rect 220630 366868 220636 366920
rect 220688 366908 220694 366920
rect 230198 366908 230204 366920
rect 220688 366880 230204 366908
rect 220688 366868 220694 366880
rect 230198 366868 230204 366880
rect 230256 366868 230262 366920
rect 144638 366800 144644 366852
rect 144696 366840 144702 366852
rect 154850 366840 154856 366852
rect 144696 366812 154856 366840
rect 144696 366800 144702 366812
rect 154850 366800 154856 366812
rect 154908 366800 154914 366852
rect 124030 366324 124036 366376
rect 124088 366364 124094 366376
rect 155218 366364 155224 366376
rect 124088 366336 155224 366364
rect 124088 366324 124094 366336
rect 155218 366324 155224 366336
rect 155276 366324 155282 366376
rect 219434 366324 219440 366376
rect 219492 366364 219498 366376
rect 250898 366364 250904 366376
rect 219492 366336 250904 366364
rect 219492 366324 219498 366336
rect 250898 366324 250904 366336
rect 250956 366324 250962 366376
rect 151538 365644 151544 365696
rect 151596 365684 151602 365696
rect 154942 365684 154948 365696
rect 151596 365656 154948 365684
rect 151596 365644 151602 365656
rect 154942 365644 154948 365656
rect 155000 365644 155006 365696
rect 220630 365644 220636 365696
rect 220688 365684 220694 365696
rect 243998 365684 244004 365696
rect 220688 365656 244004 365684
rect 220688 365644 220694 365656
rect 243998 365644 244004 365656
rect 244056 365644 244062 365696
rect 133414 365576 133420 365628
rect 133472 365616 133478 365628
rect 155126 365616 155132 365628
rect 133472 365588 155132 365616
rect 133472 365576 133478 365588
rect 155126 365576 155132 365588
rect 155184 365576 155190 365628
rect 219710 365576 219716 365628
rect 219768 365616 219774 365628
rect 230290 365616 230296 365628
rect 219768 365588 230296 365616
rect 219768 365576 219774 365588
rect 230290 365576 230296 365588
rect 230348 365576 230354 365628
rect 134794 365508 134800 365560
rect 134852 365548 134858 365560
rect 154850 365548 154856 365560
rect 134852 365520 154856 365548
rect 134852 365508 134858 365520
rect 154850 365508 154856 365520
rect 154908 365508 154914 365560
rect 137554 365440 137560 365492
rect 137612 365480 137618 365492
rect 154666 365480 154672 365492
rect 137612 365452 154672 365480
rect 137612 365440 137618 365452
rect 154666 365440 154672 365452
rect 154724 365440 154730 365492
rect 112990 365372 112996 365424
rect 113048 365412 113054 365424
rect 154758 365412 154764 365424
rect 113048 365384 154764 365412
rect 113048 365372 113054 365384
rect 154758 365372 154764 365384
rect 154816 365372 154822 365424
rect 231118 364352 231124 364404
rect 231176 364392 231182 364404
rect 579982 364392 579988 364404
rect 231176 364364 579988 364392
rect 231176 364352 231182 364364
rect 579982 364352 579988 364364
rect 580040 364352 580046 364404
rect 123938 364284 123944 364336
rect 123996 364324 124002 364336
rect 154758 364324 154764 364336
rect 123996 364296 154764 364324
rect 123996 364284 124002 364296
rect 154758 364284 154764 364296
rect 154816 364284 154822 364336
rect 220630 364284 220636 364336
rect 220688 364324 220694 364336
rect 252094 364324 252100 364336
rect 220688 364296 252100 364324
rect 220688 364284 220694 364296
rect 252094 364284 252100 364296
rect 252152 364284 252158 364336
rect 126606 364216 126612 364268
rect 126664 364256 126670 364268
rect 155034 364256 155040 364268
rect 126664 364228 155040 364256
rect 126664 364216 126670 364228
rect 155034 364216 155040 364228
rect 155092 364216 155098 364268
rect 220722 364216 220728 364268
rect 220780 364256 220786 364268
rect 248046 364256 248052 364268
rect 220780 364228 248052 364256
rect 220780 364216 220786 364228
rect 248046 364216 248052 364228
rect 248104 364216 248110 364268
rect 128170 364148 128176 364200
rect 128228 364188 128234 364200
rect 154850 364188 154856 364200
rect 128228 364160 154856 364188
rect 128228 364148 128234 364160
rect 154850 364148 154856 364160
rect 154908 364148 154914 364200
rect 220538 364148 220544 364200
rect 220596 364188 220602 364200
rect 226058 364188 226064 364200
rect 220596 364160 226064 364188
rect 220596 364148 220602 364160
rect 226058 364148 226064 364160
rect 226116 364148 226122 364200
rect 129274 364080 129280 364132
rect 129332 364120 129338 364132
rect 154942 364120 154948 364132
rect 129332 364092 154948 364120
rect 129332 364080 129338 364092
rect 154942 364080 154948 364092
rect 155000 364080 155006 364132
rect 113082 362856 113088 362908
rect 113140 362896 113146 362908
rect 154574 362896 154580 362908
rect 113140 362868 154580 362896
rect 113140 362856 113146 362868
rect 154574 362856 154580 362868
rect 154632 362856 154638 362908
rect 114462 362788 114468 362840
rect 114520 362828 114526 362840
rect 155034 362828 155040 362840
rect 114520 362800 155040 362828
rect 114520 362788 114526 362800
rect 155034 362788 155040 362800
rect 155092 362788 155098 362840
rect 220630 362788 220636 362840
rect 220688 362828 220694 362840
rect 239858 362828 239864 362840
rect 220688 362800 239864 362828
rect 220688 362788 220694 362800
rect 239858 362788 239864 362800
rect 239916 362788 239922 362840
rect 143442 362720 143448 362772
rect 143500 362760 143506 362772
rect 154850 362760 154856 362772
rect 143500 362732 154856 362760
rect 143500 362720 143506 362732
rect 154850 362720 154856 362732
rect 154908 362720 154914 362772
rect 220722 362720 220728 362772
rect 220780 362760 220786 362772
rect 238478 362760 238484 362772
rect 220780 362732 238484 362760
rect 220780 362720 220786 362732
rect 238478 362720 238484 362732
rect 238536 362720 238542 362772
rect 145834 362652 145840 362704
rect 145892 362692 145898 362704
rect 154942 362692 154948 362704
rect 145892 362664 154948 362692
rect 145892 362652 145898 362664
rect 154942 362652 154948 362664
rect 155000 362652 155006 362704
rect 220538 362652 220544 362704
rect 220596 362692 220602 362704
rect 252278 362692 252284 362704
rect 220596 362664 252284 362692
rect 220596 362652 220602 362664
rect 252278 362652 252284 362664
rect 252336 362652 252342 362704
rect 122742 362176 122748 362228
rect 122800 362216 122806 362228
rect 155402 362216 155408 362228
rect 122800 362188 155408 362216
rect 122800 362176 122806 362188
rect 155402 362176 155408 362188
rect 155460 362176 155466 362228
rect 220630 362176 220636 362228
rect 220688 362216 220694 362228
rect 239950 362216 239956 362228
rect 220688 362188 239956 362216
rect 220688 362176 220694 362188
rect 239950 362176 239956 362188
rect 240008 362176 240014 362228
rect 220446 362108 220452 362160
rect 220504 362148 220510 362160
rect 223390 362148 223396 362160
rect 220504 362120 223396 362148
rect 220504 362108 220510 362120
rect 223390 362108 223396 362120
rect 223448 362108 223454 362160
rect 115842 361496 115848 361548
rect 115900 361536 115906 361548
rect 155034 361536 155040 361548
rect 115900 361508 155040 361536
rect 115900 361496 115906 361508
rect 155034 361496 155040 361508
rect 155092 361496 155098 361548
rect 220722 361496 220728 361548
rect 220780 361536 220786 361548
rect 241238 361536 241244 361548
rect 220780 361508 241244 361536
rect 220780 361496 220786 361508
rect 241238 361496 241244 361508
rect 241296 361496 241302 361548
rect 129366 361428 129372 361480
rect 129424 361468 129430 361480
rect 154758 361468 154764 361480
rect 129424 361440 154764 361468
rect 129424 361428 129430 361440
rect 154758 361428 154764 361440
rect 154816 361428 154822 361480
rect 132126 361360 132132 361412
rect 132184 361400 132190 361412
rect 154850 361400 154856 361412
rect 132184 361372 154856 361400
rect 132184 361360 132190 361372
rect 154850 361360 154856 361372
rect 154908 361360 154914 361412
rect 133506 361292 133512 361344
rect 133564 361332 133570 361344
rect 154574 361332 154580 361344
rect 133564 361304 154580 361332
rect 133564 361292 133570 361304
rect 154574 361292 154580 361304
rect 154632 361292 154638 361344
rect 136082 361224 136088 361276
rect 136140 361264 136146 361276
rect 154942 361264 154948 361276
rect 136140 361236 154948 361264
rect 136140 361224 136146 361236
rect 154942 361224 154948 361236
rect 155000 361224 155006 361276
rect 219894 361088 219900 361140
rect 219952 361128 219958 361140
rect 223482 361128 223488 361140
rect 219952 361100 223488 361128
rect 219952 361088 219958 361100
rect 223482 361088 223488 361100
rect 223540 361088 223546 361140
rect 220446 360884 220452 360936
rect 220504 360924 220510 360936
rect 226886 360924 226892 360936
rect 220504 360896 226892 360924
rect 220504 360884 220510 360896
rect 226886 360884 226892 360896
rect 226944 360884 226950 360936
rect 220354 360816 220360 360868
rect 220412 360856 220418 360868
rect 242618 360856 242624 360868
rect 220412 360828 242624 360856
rect 220412 360816 220418 360828
rect 242618 360816 242624 360828
rect 242676 360816 242682 360868
rect 122558 360136 122564 360188
rect 122616 360176 122622 360188
rect 154574 360176 154580 360188
rect 122616 360148 154580 360176
rect 122616 360136 122622 360148
rect 154574 360136 154580 360148
rect 154632 360136 154638 360188
rect 220630 360136 220636 360188
rect 220688 360176 220694 360188
rect 252370 360176 252376 360188
rect 220688 360148 252376 360176
rect 220688 360136 220694 360148
rect 252370 360136 252376 360148
rect 252428 360136 252434 360188
rect 126698 360068 126704 360120
rect 126756 360108 126762 360120
rect 155034 360108 155040 360120
rect 126756 360080 155040 360108
rect 126756 360068 126762 360080
rect 155034 360068 155040 360080
rect 155092 360068 155098 360120
rect 219710 360068 219716 360120
rect 219768 360108 219774 360120
rect 242526 360108 242532 360120
rect 219768 360080 242532 360108
rect 219768 360068 219774 360080
rect 242526 360068 242532 360080
rect 242584 360068 242590 360120
rect 128262 360000 128268 360052
rect 128320 360040 128326 360052
rect 154942 360040 154948 360052
rect 128320 360012 154948 360040
rect 128320 360000 128326 360012
rect 154942 360000 154948 360012
rect 155000 360000 155006 360052
rect 220722 360000 220728 360052
rect 220780 360040 220786 360052
rect 231578 360040 231584 360052
rect 220780 360012 231584 360040
rect 220780 360000 220786 360012
rect 231578 360000 231584 360012
rect 231636 360000 231642 360052
rect 141970 359932 141976 359984
rect 142028 359972 142034 359984
rect 154850 359972 154856 359984
rect 142028 359944 154856 359972
rect 142028 359932 142034 359944
rect 154850 359932 154856 359944
rect 154908 359932 154914 359984
rect 147490 359864 147496 359916
rect 147548 359904 147554 359916
rect 154942 359904 154948 359916
rect 147548 359876 154948 359904
rect 147548 359864 147554 359876
rect 154942 359864 154948 359876
rect 155000 359864 155006 359916
rect 219894 359456 219900 359508
rect 219952 359496 219958 359508
rect 246206 359496 246212 359508
rect 219952 359468 246212 359496
rect 219952 359456 219958 359468
rect 246206 359456 246212 359468
rect 246264 359456 246270 359508
rect 220722 359252 220728 359304
rect 220780 359292 220786 359304
rect 226794 359292 226800 359304
rect 220780 359264 226800 359292
rect 220780 359252 220786 359264
rect 226794 359252 226800 359264
rect 226852 359252 226858 359304
rect 152918 358708 152924 358760
rect 152976 358748 152982 358760
rect 155586 358748 155592 358760
rect 152976 358720 155592 358748
rect 152976 358708 152982 358720
rect 155586 358708 155592 358720
rect 155644 358708 155650 358760
rect 220630 358708 220636 358760
rect 220688 358748 220694 358760
rect 231670 358748 231676 358760
rect 220688 358720 231676 358748
rect 220688 358708 220694 358720
rect 231670 358708 231676 358720
rect 231728 358708 231734 358760
rect 117222 358640 117228 358692
rect 117280 358680 117286 358692
rect 154942 358680 154948 358692
rect 117280 358652 154948 358680
rect 117280 358640 117286 358652
rect 154942 358640 154948 358652
rect 155000 358640 155006 358692
rect 219986 358640 219992 358692
rect 220044 358680 220050 358692
rect 228634 358680 228640 358692
rect 220044 358652 228640 358680
rect 220044 358640 220050 358652
rect 228634 358640 228640 358652
rect 228692 358640 228698 358692
rect 137646 358572 137652 358624
rect 137704 358612 137710 358624
rect 154758 358612 154764 358624
rect 137704 358584 154764 358612
rect 137704 358572 137710 358584
rect 154758 358572 154764 358584
rect 154816 358572 154822 358624
rect 115106 358504 115112 358556
rect 115164 358544 115170 358556
rect 154574 358544 154580 358556
rect 115164 358516 154580 358544
rect 115164 358504 115170 358516
rect 154574 358504 154580 358516
rect 154632 358504 154638 358556
rect 220538 358028 220544 358080
rect 220596 358068 220602 358080
rect 238570 358068 238576 358080
rect 220596 358040 238576 358068
rect 220596 358028 220602 358040
rect 238570 358028 238576 358040
rect 238628 358028 238634 358080
rect 2958 357416 2964 357468
rect 3016 357456 3022 357468
rect 156782 357456 156788 357468
rect 3016 357428 156788 357456
rect 3016 357416 3022 357428
rect 156782 357416 156788 357428
rect 156840 357416 156846 357468
rect 151630 357348 151636 357400
rect 151688 357388 151694 357400
rect 155034 357388 155040 357400
rect 151688 357360 155040 357388
rect 151688 357348 151694 357360
rect 155034 357348 155040 357360
rect 155092 357348 155098 357400
rect 220722 357348 220728 357400
rect 220780 357388 220786 357400
rect 231762 357388 231768 357400
rect 220780 357360 231768 357388
rect 220780 357348 220786 357360
rect 231762 357348 231768 357360
rect 231820 357348 231826 357400
rect 126882 357280 126888 357332
rect 126940 357320 126946 357332
rect 154758 357320 154764 357332
rect 126940 357292 154764 357320
rect 126940 357280 126946 357292
rect 154758 357280 154764 357292
rect 154816 357280 154822 357332
rect 132218 357212 132224 357264
rect 132276 357252 132282 357264
rect 154942 357252 154948 357264
rect 132276 357224 154948 357252
rect 132276 357212 132282 357224
rect 154942 357212 154948 357224
rect 155000 357212 155006 357264
rect 220630 357212 220636 357264
rect 220688 357252 220694 357264
rect 222010 357252 222016 357264
rect 220688 357224 222016 357252
rect 220688 357212 220694 357224
rect 222010 357212 222016 357224
rect 222068 357212 222074 357264
rect 149974 357144 149980 357196
rect 150032 357184 150038 357196
rect 154850 357184 154856 357196
rect 150032 357156 154856 357184
rect 150032 357144 150038 357156
rect 154850 357144 154856 357156
rect 154908 357144 154914 357196
rect 125134 357076 125140 357128
rect 125192 357116 125198 357128
rect 154942 357116 154948 357128
rect 125192 357088 154948 357116
rect 125192 357076 125198 357088
rect 154942 357076 154948 357088
rect 155000 357076 155006 357128
rect 219894 356668 219900 356720
rect 219952 356708 219958 356720
rect 248966 356708 248972 356720
rect 219952 356680 248972 356708
rect 219952 356668 219958 356680
rect 248966 356668 248972 356680
rect 249024 356668 249030 356720
rect 153010 355988 153016 356040
rect 153068 356028 153074 356040
rect 154574 356028 154580 356040
rect 153068 356000 154580 356028
rect 153068 355988 153074 356000
rect 154574 355988 154580 356000
rect 154632 355988 154638 356040
rect 220722 355988 220728 356040
rect 220780 356028 220786 356040
rect 246942 356028 246948 356040
rect 220780 356000 246948 356028
rect 220780 355988 220786 356000
rect 246942 355988 246948 356000
rect 247000 355988 247006 356040
rect 137738 355920 137744 355972
rect 137796 355960 137802 355972
rect 155034 355960 155040 355972
rect 137796 355932 155040 355960
rect 137796 355920 137802 355932
rect 155034 355920 155040 355932
rect 155092 355920 155098 355972
rect 144730 355852 144736 355904
rect 144788 355892 144794 355904
rect 154850 355892 154856 355904
rect 144788 355864 154856 355892
rect 144788 355852 144794 355864
rect 154850 355852 154856 355864
rect 154908 355852 154914 355904
rect 119890 355784 119896 355836
rect 119948 355824 119954 355836
rect 154942 355824 154948 355836
rect 119948 355796 154948 355824
rect 119948 355784 119954 355796
rect 154942 355784 154948 355796
rect 155000 355784 155006 355836
rect 219802 355784 219808 355836
rect 219860 355824 219866 355836
rect 224126 355824 224132 355836
rect 219860 355796 224132 355824
rect 219860 355784 219866 355796
rect 224126 355784 224132 355796
rect 224184 355784 224190 355836
rect 220722 355716 220728 355768
rect 220780 355756 220786 355768
rect 226150 355756 226156 355768
rect 220780 355728 226156 355756
rect 220780 355716 220786 355728
rect 226150 355716 226156 355728
rect 226208 355716 226214 355768
rect 130930 355376 130936 355428
rect 130988 355416 130994 355428
rect 155586 355416 155592 355428
rect 130988 355388 155592 355416
rect 130988 355376 130994 355388
rect 155586 355376 155592 355388
rect 155644 355376 155650 355428
rect 119246 355308 119252 355360
rect 119304 355348 119310 355360
rect 155126 355348 155132 355360
rect 119304 355320 155132 355348
rect 119304 355308 119310 355320
rect 155126 355308 155132 355320
rect 155184 355308 155190 355360
rect 112254 354628 112260 354680
rect 112312 354668 112318 354680
rect 154850 354668 154856 354680
rect 112312 354640 154856 354668
rect 112312 354628 112318 354640
rect 154850 354628 154856 354640
rect 154908 354628 154914 354680
rect 220722 354628 220728 354680
rect 220780 354668 220786 354680
rect 245378 354668 245384 354680
rect 220780 354640 245384 354668
rect 220780 354628 220786 354640
rect 245378 354628 245384 354640
rect 245436 354628 245442 354680
rect 112346 354560 112352 354612
rect 112404 354600 112410 354612
rect 154574 354600 154580 354612
rect 112404 354572 154580 354600
rect 112404 354560 112410 354572
rect 154574 354560 154580 354572
rect 154632 354560 154638 354612
rect 116394 354492 116400 354544
rect 116452 354532 116458 354544
rect 154942 354532 154948 354544
rect 116452 354504 154948 354532
rect 116452 354492 116458 354504
rect 154942 354492 154948 354504
rect 155000 354492 155006 354544
rect 133598 354424 133604 354476
rect 133656 354464 133662 354476
rect 154758 354464 154764 354476
rect 133656 354436 154764 354464
rect 133656 354424 133662 354436
rect 154758 354424 154764 354436
rect 154816 354424 154822 354476
rect 220630 354356 220636 354408
rect 220688 354396 220694 354408
rect 228726 354396 228732 354408
rect 220688 354368 228732 354396
rect 220688 354356 220694 354368
rect 228726 354356 228732 354368
rect 228784 354356 228790 354408
rect 220630 353948 220636 354000
rect 220688 353988 220694 354000
rect 251082 353988 251088 354000
rect 220688 353960 251088 353988
rect 220688 353948 220694 353960
rect 251082 353948 251088 353960
rect 251140 353948 251146 354000
rect 115014 353200 115020 353252
rect 115072 353240 115078 353252
rect 154758 353240 154764 353252
rect 115072 353212 154764 353240
rect 115072 353200 115078 353212
rect 154758 353200 154764 353212
rect 154816 353200 154822 353252
rect 220722 353200 220728 353252
rect 220780 353240 220786 353252
rect 245470 353240 245476 353252
rect 220780 353212 245476 353240
rect 220780 353200 220786 353212
rect 245470 353200 245476 353212
rect 245528 353200 245534 353252
rect 132402 353132 132408 353184
rect 132460 353172 132466 353184
rect 154942 353172 154948 353184
rect 132460 353144 154948 353172
rect 132460 353132 132466 353144
rect 154942 353132 154948 353144
rect 155000 353132 155006 353184
rect 132310 353064 132316 353116
rect 132368 353104 132374 353116
rect 154850 353104 154856 353116
rect 132368 353076 154856 353104
rect 132368 353064 132374 353076
rect 154850 353064 154856 353076
rect 154908 353064 154914 353116
rect 139210 352996 139216 353048
rect 139268 353036 139274 353048
rect 155034 353036 155040 353048
rect 139268 353008 155040 353036
rect 139268 352996 139274 353008
rect 155034 352996 155040 353008
rect 155092 352996 155098 353048
rect 142062 352928 142068 352980
rect 142120 352968 142126 352980
rect 154850 352968 154856 352980
rect 142120 352940 154856 352968
rect 142120 352928 142126 352940
rect 154850 352928 154856 352940
rect 154908 352928 154914 352980
rect 220446 352724 220452 352776
rect 220504 352764 220510 352776
rect 228818 352764 228824 352776
rect 220504 352736 228824 352764
rect 220504 352724 220510 352736
rect 228818 352724 228824 352736
rect 228876 352724 228882 352776
rect 220446 352452 220452 352504
rect 220504 352492 220510 352504
rect 222746 352492 222752 352504
rect 220504 352464 222752 352492
rect 220504 352452 220510 352464
rect 222746 352452 222752 352464
rect 222804 352452 222810 352504
rect 258718 351908 258724 351960
rect 258776 351948 258782 351960
rect 580166 351948 580172 351960
rect 258776 351920 580172 351948
rect 258776 351908 258782 351920
rect 580166 351908 580172 351920
rect 580224 351908 580230 351960
rect 119982 351840 119988 351892
rect 120040 351880 120046 351892
rect 154850 351880 154856 351892
rect 120040 351852 154856 351880
rect 120040 351840 120046 351852
rect 154850 351840 154856 351852
rect 154908 351840 154914 351892
rect 220722 351840 220728 351892
rect 220780 351880 220786 351892
rect 250990 351880 250996 351892
rect 220780 351852 250996 351880
rect 220780 351840 220786 351852
rect 250990 351840 250996 351852
rect 251048 351840 251054 351892
rect 124122 351772 124128 351824
rect 124180 351812 124186 351824
rect 154942 351812 154948 351824
rect 124180 351784 154948 351812
rect 124180 351772 124186 351784
rect 154942 351772 154948 351784
rect 155000 351772 155006 351824
rect 145926 351704 145932 351756
rect 145984 351744 145990 351756
rect 155034 351744 155040 351756
rect 145984 351716 155040 351744
rect 145984 351704 145990 351716
rect 155034 351704 155040 351716
rect 155092 351704 155098 351756
rect 148870 351636 148876 351688
rect 148928 351676 148934 351688
rect 154758 351676 154764 351688
rect 148928 351648 154764 351676
rect 148928 351636 148934 351648
rect 154758 351636 154764 351648
rect 154816 351636 154822 351688
rect 219986 351296 219992 351348
rect 220044 351336 220050 351348
rect 228910 351336 228916 351348
rect 220044 351308 228916 351336
rect 220044 351296 220050 351308
rect 228910 351296 228916 351308
rect 228968 351296 228974 351348
rect 219894 351024 219900 351076
rect 219952 351064 219958 351076
rect 226242 351064 226248 351076
rect 219952 351036 226248 351064
rect 219952 351024 219958 351036
rect 226242 351024 226248 351036
rect 226300 351024 226306 351076
rect 116486 350480 116492 350532
rect 116544 350520 116550 350532
rect 154574 350520 154580 350532
rect 116544 350492 154580 350520
rect 116544 350480 116550 350492
rect 154574 350480 154580 350492
rect 154632 350480 154638 350532
rect 220538 350480 220544 350532
rect 220596 350520 220602 350532
rect 244182 350520 244188 350532
rect 220596 350492 244188 350520
rect 220596 350480 220602 350492
rect 244182 350480 244188 350492
rect 244240 350480 244246 350532
rect 140682 350412 140688 350464
rect 140740 350452 140746 350464
rect 154942 350452 154948 350464
rect 140740 350424 154948 350452
rect 140740 350412 140746 350424
rect 154942 350412 154948 350424
rect 155000 350412 155006 350464
rect 219894 350208 219900 350260
rect 219952 350248 219958 350260
rect 229002 350248 229008 350260
rect 219952 350220 229008 350248
rect 219952 350208 219958 350220
rect 229002 350208 229008 350220
rect 229060 350208 229066 350260
rect 220722 349800 220728 349852
rect 220780 349840 220786 349852
rect 245562 349840 245568 349852
rect 220780 349812 245568 349840
rect 220780 349800 220786 349812
rect 245562 349800 245568 349812
rect 245620 349800 245626 349852
rect 138750 349188 138756 349240
rect 138808 349228 138814 349240
rect 154942 349228 154948 349240
rect 138808 349200 154948 349228
rect 138808 349188 138814 349200
rect 154942 349188 154948 349200
rect 155000 349188 155006 349240
rect 126238 349120 126244 349172
rect 126296 349160 126302 349172
rect 154850 349160 154856 349172
rect 126296 349132 154856 349160
rect 126296 349120 126302 349132
rect 154850 349120 154856 349132
rect 154908 349120 154914 349172
rect 220630 349052 220636 349104
rect 220688 349092 220694 349104
rect 248138 349092 248144 349104
rect 220688 349064 248144 349092
rect 220688 349052 220694 349064
rect 248138 349052 248144 349064
rect 248196 349052 248202 349104
rect 220538 348984 220544 349036
rect 220596 349024 220602 349036
rect 224034 349024 224040 349036
rect 220596 348996 224040 349024
rect 220596 348984 220602 348996
rect 224034 348984 224040 348996
rect 224092 348984 224098 349036
rect 220538 348372 220544 348424
rect 220596 348412 220602 348424
rect 236638 348412 236644 348424
rect 220596 348384 236644 348412
rect 220596 348372 220602 348384
rect 236638 348372 236644 348384
rect 236696 348372 236702 348424
rect 220446 348032 220452 348084
rect 220504 348072 220510 348084
rect 223942 348072 223948 348084
rect 220504 348044 223948 348072
rect 220504 348032 220510 348044
rect 223942 348032 223948 348044
rect 224000 348032 224006 348084
rect 122650 347964 122656 348016
rect 122708 348004 122714 348016
rect 154850 348004 154856 348016
rect 122708 347976 154856 348004
rect 122708 347964 122714 347976
rect 154850 347964 154856 347976
rect 154908 347964 154914 348016
rect 119430 347896 119436 347948
rect 119488 347936 119494 347948
rect 154942 347936 154948 347948
rect 119488 347908 154948 347936
rect 119488 347896 119494 347908
rect 154942 347896 154948 347908
rect 155000 347896 155006 347948
rect 119522 347828 119528 347880
rect 119580 347868 119586 347880
rect 154758 347868 154764 347880
rect 119580 347840 154764 347868
rect 119580 347828 119586 347840
rect 154758 347828 154764 347840
rect 154816 347828 154822 347880
rect 116670 347760 116676 347812
rect 116728 347800 116734 347812
rect 155034 347800 155040 347812
rect 116728 347772 155040 347800
rect 116728 347760 116734 347772
rect 155034 347760 155040 347772
rect 155092 347760 155098 347812
rect 220446 347692 220452 347744
rect 220504 347732 220510 347744
rect 234154 347732 234160 347744
rect 220504 347704 234160 347732
rect 220504 347692 220510 347704
rect 234154 347692 234160 347704
rect 234212 347692 234218 347744
rect 220722 347624 220728 347676
rect 220780 347664 220786 347676
rect 233970 347664 233976 347676
rect 220780 347636 233976 347664
rect 220780 347624 220786 347636
rect 233970 347624 233976 347636
rect 234028 347624 234034 347676
rect 220630 347556 220636 347608
rect 220688 347596 220694 347608
rect 231026 347596 231032 347608
rect 220688 347568 231032 347596
rect 220688 347556 220694 347568
rect 231026 347556 231032 347568
rect 231084 347556 231090 347608
rect 118234 347012 118240 347064
rect 118292 347052 118298 347064
rect 154942 347052 154948 347064
rect 118292 347024 154948 347052
rect 118292 347012 118298 347024
rect 154942 347012 154948 347024
rect 155000 347012 155006 347064
rect 142982 346604 142988 346656
rect 143040 346644 143046 346656
rect 154850 346644 154856 346656
rect 143040 346616 154856 346644
rect 143040 346604 143046 346616
rect 154850 346604 154856 346616
rect 154908 346604 154914 346656
rect 136174 346536 136180 346588
rect 136232 346576 136238 346588
rect 154942 346576 154948 346588
rect 136232 346548 154948 346576
rect 136232 346536 136238 346548
rect 154942 346536 154948 346548
rect 155000 346536 155006 346588
rect 116578 346468 116584 346520
rect 116636 346508 116642 346520
rect 155034 346508 155040 346520
rect 116636 346480 155040 346508
rect 116636 346468 116642 346480
rect 155034 346468 155040 346480
rect 155092 346468 155098 346520
rect 113910 346400 113916 346452
rect 113968 346440 113974 346452
rect 154574 346440 154580 346452
rect 113968 346412 154580 346440
rect 113968 346400 113974 346412
rect 154574 346400 154580 346412
rect 154632 346400 154638 346452
rect 220630 346332 220636 346384
rect 220688 346372 220694 346384
rect 252462 346372 252468 346384
rect 220688 346344 252468 346372
rect 220688 346332 220694 346344
rect 252462 346332 252468 346344
rect 252520 346332 252526 346384
rect 220722 346264 220728 346316
rect 220780 346304 220786 346316
rect 229738 346304 229744 346316
rect 220780 346276 229744 346304
rect 220780 346264 220786 346276
rect 229738 346264 229744 346276
rect 229796 346264 229802 346316
rect 220722 345924 220728 345976
rect 220780 345964 220786 345976
rect 222102 345964 222108 345976
rect 220780 345936 222108 345964
rect 220780 345924 220786 345936
rect 222102 345924 222108 345936
rect 222160 345924 222166 345976
rect 122098 345652 122104 345704
rect 122156 345692 122162 345704
rect 154850 345692 154856 345704
rect 122156 345664 154856 345692
rect 122156 345652 122162 345664
rect 154850 345652 154856 345664
rect 154908 345652 154914 345704
rect 141510 345176 141516 345228
rect 141568 345216 141574 345228
rect 154942 345216 154948 345228
rect 141568 345188 154948 345216
rect 141568 345176 141574 345188
rect 154942 345176 154948 345188
rect 155000 345176 155006 345228
rect 113818 345108 113824 345160
rect 113876 345148 113882 345160
rect 155034 345148 155040 345160
rect 113876 345120 155040 345148
rect 113876 345108 113882 345120
rect 155034 345108 155040 345120
rect 155092 345108 155098 345160
rect 3050 345040 3056 345092
rect 3108 345080 3114 345092
rect 135990 345080 135996 345092
rect 3108 345052 135996 345080
rect 3108 345040 3114 345052
rect 135990 345040 135996 345052
rect 136048 345040 136054 345092
rect 140130 345040 140136 345092
rect 140188 345080 140194 345092
rect 154942 345080 154948 345092
rect 140188 345052 154948 345080
rect 140188 345040 140194 345052
rect 154942 345040 154948 345052
rect 155000 345040 155006 345092
rect 220630 344972 220636 345024
rect 220688 345012 220694 345024
rect 250438 345012 250444 345024
rect 220688 344984 250444 345012
rect 220688 344972 220694 344984
rect 250438 344972 250444 344984
rect 250496 344972 250502 345024
rect 220722 344904 220728 344956
rect 220780 344944 220786 344956
rect 231210 344944 231216 344956
rect 220780 344916 231216 344944
rect 220780 344904 220786 344916
rect 231210 344904 231216 344916
rect 231268 344904 231274 344956
rect 219894 343884 219900 343936
rect 219952 343924 219958 343936
rect 226978 343924 226984 343936
rect 219952 343896 226984 343924
rect 219952 343884 219958 343896
rect 226978 343884 226984 343896
rect 227036 343884 227042 343936
rect 131758 343816 131764 343868
rect 131816 343856 131822 343868
rect 154574 343856 154580 343868
rect 131816 343828 154580 343856
rect 131816 343816 131822 343828
rect 154574 343816 154580 343828
rect 154632 343816 154638 343868
rect 123478 343748 123484 343800
rect 123536 343788 123542 343800
rect 154942 343788 154948 343800
rect 123536 343760 154948 343788
rect 123536 343748 123542 343760
rect 154942 343748 154948 343760
rect 155000 343748 155006 343800
rect 120718 343680 120724 343732
rect 120776 343720 120782 343732
rect 155034 343720 155040 343732
rect 120776 343692 155040 343720
rect 120776 343680 120782 343692
rect 155034 343680 155040 343692
rect 155092 343680 155098 343732
rect 119338 343612 119344 343664
rect 119396 343652 119402 343664
rect 154850 343652 154856 343664
rect 119396 343624 154856 343652
rect 119396 343612 119402 343624
rect 154850 343612 154856 343624
rect 154908 343612 154914 343664
rect 220722 343544 220728 343596
rect 220780 343584 220786 343596
rect 247770 343584 247776 343596
rect 220780 343556 247776 343584
rect 220780 343544 220786 343556
rect 247770 343544 247776 343556
rect 247828 343544 247834 343596
rect 220630 343340 220636 343392
rect 220688 343380 220694 343392
rect 222838 343380 222844 343392
rect 220688 343352 222844 343380
rect 220688 343340 220694 343352
rect 222838 343340 222844 343352
rect 222896 343340 222902 343392
rect 115198 342864 115204 342916
rect 115256 342904 115262 342916
rect 154574 342904 154580 342916
rect 115256 342876 154580 342904
rect 115256 342864 115262 342876
rect 154574 342864 154580 342876
rect 154632 342864 154638 342916
rect 220446 342524 220452 342576
rect 220504 342564 220510 342576
rect 221734 342564 221740 342576
rect 220504 342536 221740 342564
rect 220504 342524 220510 342536
rect 221734 342524 221740 342536
rect 221792 342524 221798 342576
rect 144546 342388 144552 342440
rect 144604 342428 144610 342440
rect 154850 342428 154856 342440
rect 144604 342400 154856 342428
rect 144604 342388 144610 342400
rect 154850 342388 154856 342400
rect 154908 342388 154914 342440
rect 139210 342320 139216 342372
rect 139268 342360 139274 342372
rect 154942 342360 154948 342372
rect 139268 342332 154948 342360
rect 139268 342320 139274 342332
rect 154942 342320 154948 342332
rect 155000 342320 155006 342372
rect 115842 342252 115848 342304
rect 115900 342292 115906 342304
rect 155034 342292 155040 342304
rect 115900 342264 155040 342292
rect 115900 342252 115906 342264
rect 155034 342252 155040 342264
rect 155092 342252 155098 342304
rect 220722 342116 220728 342168
rect 220780 342156 220786 342168
rect 251910 342156 251916 342168
rect 220780 342128 251916 342156
rect 220780 342116 220786 342128
rect 251910 342116 251916 342128
rect 251968 342116 251974 342168
rect 219802 341912 219808 341964
rect 219860 341952 219866 341964
rect 221642 341952 221648 341964
rect 219860 341924 221648 341952
rect 219860 341912 219866 341924
rect 221642 341912 221648 341924
rect 221700 341912 221706 341964
rect 128170 341096 128176 341148
rect 128228 341136 128234 341148
rect 154942 341136 154948 341148
rect 128228 341108 154948 341136
rect 128228 341096 128234 341108
rect 154942 341096 154948 341108
rect 155000 341096 155006 341148
rect 124030 341028 124036 341080
rect 124088 341068 124094 341080
rect 154758 341068 154764 341080
rect 124088 341040 154764 341068
rect 124088 341028 124094 341040
rect 154758 341028 154764 341040
rect 154816 341028 154822 341080
rect 121178 340960 121184 341012
rect 121236 341000 121242 341012
rect 155034 341000 155040 341012
rect 121236 340972 155040 341000
rect 121236 340960 121242 340972
rect 155034 340960 155040 340972
rect 155092 340960 155098 341012
rect 117130 340892 117136 340944
rect 117188 340932 117194 340944
rect 154850 340932 154856 340944
rect 117188 340904 154856 340932
rect 117188 340892 117194 340904
rect 154850 340892 154856 340904
rect 154908 340892 154914 340944
rect 219526 340824 219532 340876
rect 219584 340864 219590 340876
rect 249150 340864 249156 340876
rect 219584 340836 249156 340864
rect 219584 340824 219590 340836
rect 249150 340824 249156 340836
rect 249208 340824 249214 340876
rect 219894 340484 219900 340536
rect 219952 340524 219958 340536
rect 227070 340524 227076 340536
rect 219952 340496 227076 340524
rect 219952 340484 219958 340496
rect 227070 340484 227076 340496
rect 227128 340484 227134 340536
rect 155310 340144 155316 340196
rect 155368 340184 155374 340196
rect 155586 340184 155592 340196
rect 155368 340156 155592 340184
rect 155368 340144 155374 340156
rect 155586 340144 155592 340156
rect 155644 340144 155650 340196
rect 147490 339736 147496 339788
rect 147548 339776 147554 339788
rect 154942 339776 154948 339788
rect 147548 339748 154948 339776
rect 147548 339736 147554 339748
rect 154942 339736 154948 339748
rect 155000 339736 155006 339788
rect 141786 339668 141792 339720
rect 141844 339708 141850 339720
rect 154850 339708 154856 339720
rect 141844 339680 154856 339708
rect 141844 339668 141850 339680
rect 154850 339668 154856 339680
rect 154908 339668 154914 339720
rect 137278 339600 137284 339652
rect 137336 339640 137342 339652
rect 155034 339640 155040 339652
rect 137336 339612 155040 339640
rect 137336 339600 137342 339612
rect 155034 339600 155040 339612
rect 155092 339600 155098 339652
rect 134702 339532 134708 339584
rect 134760 339572 134766 339584
rect 154942 339572 154948 339584
rect 134760 339544 154948 339572
rect 134760 339532 134766 339544
rect 154942 339532 154948 339544
rect 155000 339532 155006 339584
rect 133230 339464 133236 339516
rect 133288 339504 133294 339516
rect 154758 339504 154764 339516
rect 133288 339476 154764 339504
rect 133288 339464 133294 339476
rect 154758 339464 154764 339476
rect 154816 339464 154822 339516
rect 220722 339396 220728 339448
rect 220780 339436 220786 339448
rect 251726 339436 251732 339448
rect 220780 339408 251732 339436
rect 220780 339396 220786 339408
rect 251726 339396 251732 339408
rect 251784 339396 251790 339448
rect 220630 339328 220636 339380
rect 220688 339368 220694 339380
rect 251634 339368 251640 339380
rect 220688 339340 251640 339368
rect 220688 339328 220694 339340
rect 251634 339328 251640 339340
rect 251692 339328 251698 339380
rect 220446 339260 220452 339312
rect 220504 339300 220510 339312
rect 234246 339300 234252 339312
rect 220504 339272 234252 339300
rect 220504 339260 220510 339272
rect 234246 339260 234252 339272
rect 234304 339260 234310 339312
rect 117222 338716 117228 338768
rect 117280 338756 117286 338768
rect 154574 338756 154580 338768
rect 117280 338728 154580 338756
rect 117280 338716 117286 338728
rect 154574 338716 154580 338728
rect 154632 338716 154638 338768
rect 148870 338308 148876 338360
rect 148928 338348 148934 338360
rect 154942 338348 154948 338360
rect 148928 338320 154948 338348
rect 148928 338308 148934 338320
rect 154942 338308 154948 338320
rect 155000 338308 155006 338360
rect 144730 338240 144736 338292
rect 144788 338280 144794 338292
rect 154850 338280 154856 338292
rect 144788 338252 154856 338280
rect 144788 338240 144794 338252
rect 154850 338240 154856 338252
rect 154908 338240 154914 338292
rect 126790 338172 126796 338224
rect 126848 338212 126854 338224
rect 154666 338212 154672 338224
rect 126848 338184 154672 338212
rect 126848 338172 126854 338184
rect 154666 338172 154672 338184
rect 154724 338172 154730 338224
rect 125134 338104 125140 338156
rect 125192 338144 125198 338156
rect 155034 338144 155040 338156
rect 125192 338116 155040 338144
rect 125192 338104 125198 338116
rect 155034 338104 155040 338116
rect 155092 338104 155098 338156
rect 119890 337356 119896 337408
rect 119948 337396 119954 337408
rect 155126 337396 155132 337408
rect 119948 337368 155132 337396
rect 119948 337356 119954 337368
rect 155126 337356 155132 337368
rect 155184 337356 155190 337408
rect 112254 337016 112260 337068
rect 112312 337056 112318 337068
rect 154574 337056 154580 337068
rect 112312 337028 154580 337056
rect 112312 337016 112318 337028
rect 154574 337016 154580 337028
rect 154632 337016 154638 337068
rect 143350 336948 143356 337000
rect 143408 336988 143414 337000
rect 154850 336988 154856 337000
rect 143408 336960 154856 336988
rect 143408 336948 143414 336960
rect 154850 336948 154856 336960
rect 154908 336948 154914 337000
rect 139118 336880 139124 336932
rect 139176 336920 139182 336932
rect 154758 336920 154764 336932
rect 139176 336892 154764 336920
rect 139176 336880 139182 336892
rect 154758 336880 154764 336892
rect 154816 336880 154822 336932
rect 220538 336880 220544 336932
rect 220596 336920 220602 336932
rect 227070 336920 227076 336932
rect 220596 336892 227076 336920
rect 220596 336880 220602 336892
rect 227070 336880 227076 336892
rect 227128 336880 227134 336932
rect 133598 336812 133604 336864
rect 133656 336852 133662 336864
rect 154942 336852 154948 336864
rect 133656 336824 154948 336852
rect 133656 336812 133662 336824
rect 154942 336812 154948 336824
rect 155000 336812 155006 336864
rect 220722 336812 220728 336864
rect 220780 336852 220786 336864
rect 233970 336852 233976 336864
rect 220780 336824 233976 336852
rect 220780 336812 220786 336824
rect 233970 336812 233976 336824
rect 234028 336812 234034 336864
rect 151538 336744 151544 336796
rect 151596 336784 151602 336796
rect 155034 336784 155040 336796
rect 151596 336756 155040 336784
rect 151596 336744 151602 336756
rect 155034 336744 155040 336756
rect 155092 336744 155098 336796
rect 220630 336744 220636 336796
rect 220688 336784 220694 336796
rect 247770 336784 247776 336796
rect 220688 336756 247776 336784
rect 220688 336744 220694 336756
rect 247770 336744 247776 336756
rect 247828 336744 247834 336796
rect 220630 336064 220636 336116
rect 220688 336104 220694 336116
rect 223942 336104 223948 336116
rect 220688 336076 223948 336104
rect 220688 336064 220694 336076
rect 223942 336064 223948 336076
rect 224000 336064 224006 336116
rect 119798 335588 119804 335640
rect 119856 335628 119862 335640
rect 154758 335628 154764 335640
rect 119856 335600 154764 335628
rect 119856 335588 119862 335600
rect 154758 335588 154764 335600
rect 154816 335588 154822 335640
rect 145926 335520 145932 335572
rect 145984 335560 145990 335572
rect 155034 335560 155040 335572
rect 145984 335532 155040 335560
rect 145984 335520 145990 335532
rect 155034 335520 155040 335532
rect 155092 335520 155098 335572
rect 220722 335520 220728 335572
rect 220780 335560 220786 335572
rect 222930 335560 222936 335572
rect 220780 335532 222936 335560
rect 220780 335520 220786 335532
rect 222930 335520 222936 335532
rect 222988 335520 222994 335572
rect 133506 335452 133512 335504
rect 133564 335492 133570 335504
rect 154850 335492 154856 335504
rect 133564 335464 154856 335492
rect 133564 335452 133570 335464
rect 154850 335452 154856 335464
rect 154908 335452 154914 335504
rect 220538 335452 220544 335504
rect 220596 335492 220602 335504
rect 246574 335492 246580 335504
rect 220596 335464 246580 335492
rect 220596 335452 220602 335464
rect 246574 335452 246580 335464
rect 246632 335452 246638 335504
rect 128078 335384 128084 335436
rect 128136 335424 128142 335436
rect 154666 335424 154672 335436
rect 128136 335396 154672 335424
rect 128136 335384 128142 335396
rect 154666 335384 154672 335396
rect 154724 335384 154730 335436
rect 151446 335316 151452 335368
rect 151504 335356 151510 335368
rect 154942 335356 154948 335368
rect 151504 335328 154948 335356
rect 151504 335316 151510 335328
rect 154942 335316 154948 335328
rect 155000 335316 155006 335368
rect 155218 335316 155224 335368
rect 155276 335356 155282 335368
rect 155678 335356 155684 335368
rect 155276 335328 155684 335356
rect 155276 335316 155282 335328
rect 155678 335316 155684 335328
rect 155736 335316 155742 335368
rect 140590 334636 140596 334688
rect 140648 334676 140654 334688
rect 155034 334676 155040 334688
rect 140648 334648 155040 334676
rect 140648 334636 140654 334648
rect 155034 334636 155040 334648
rect 155092 334636 155098 334688
rect 115106 334568 115112 334620
rect 115164 334608 115170 334620
rect 155494 334608 155500 334620
rect 115164 334580 155500 334608
rect 115164 334568 115170 334580
rect 155494 334568 155500 334580
rect 155552 334568 155558 334620
rect 219894 334568 219900 334620
rect 219952 334608 219958 334620
rect 229830 334608 229836 334620
rect 219952 334580 229836 334608
rect 219952 334568 219958 334580
rect 229830 334568 229836 334580
rect 229888 334568 229894 334620
rect 132218 334092 132224 334144
rect 132276 334132 132282 334144
rect 154942 334132 154948 334144
rect 132276 334104 154948 334132
rect 132276 334092 132282 334104
rect 154942 334092 154948 334104
rect 155000 334092 155006 334144
rect 148778 334024 148784 334076
rect 148836 334064 148842 334076
rect 154758 334064 154764 334076
rect 148836 334036 154764 334064
rect 148836 334024 148842 334036
rect 154758 334024 154764 334036
rect 154816 334024 154822 334076
rect 219986 334024 219992 334076
rect 220044 334064 220050 334076
rect 222838 334064 222844 334076
rect 220044 334036 222844 334064
rect 220044 334024 220050 334036
rect 222838 334024 222844 334036
rect 222896 334024 222902 334076
rect 153010 333956 153016 334008
rect 153068 333996 153074 334008
rect 155126 333996 155132 334008
rect 153068 333968 155132 333996
rect 153068 333956 153074 333968
rect 155126 333956 155132 333968
rect 155184 333956 155190 334008
rect 220354 333956 220360 334008
rect 220412 333996 220418 334008
rect 249610 333996 249616 334008
rect 220412 333968 249616 333996
rect 220412 333956 220418 333968
rect 249610 333956 249616 333968
rect 249668 333956 249674 334008
rect 117958 333208 117964 333260
rect 118016 333248 118022 333260
rect 155402 333248 155408 333260
rect 118016 333220 155408 333248
rect 118016 333208 118022 333220
rect 155402 333208 155408 333220
rect 155460 333208 155466 333260
rect 219802 333072 219808 333124
rect 219860 333112 219866 333124
rect 227714 333112 227720 333124
rect 219860 333084 227720 333112
rect 219860 333072 219866 333084
rect 227714 333072 227720 333084
rect 227772 333072 227778 333124
rect 114462 332868 114468 332920
rect 114520 332908 114526 332920
rect 154758 332908 154764 332920
rect 114520 332880 154764 332908
rect 114520 332868 114526 332880
rect 154758 332868 154764 332880
rect 154816 332868 154822 332920
rect 145834 332800 145840 332852
rect 145892 332840 145898 332852
rect 154574 332840 154580 332852
rect 145892 332812 154580 332840
rect 145892 332800 145898 332812
rect 154574 332800 154580 332812
rect 154632 332800 154638 332852
rect 140498 332732 140504 332784
rect 140556 332772 140562 332784
rect 154942 332772 154948 332784
rect 140556 332744 154948 332772
rect 140556 332732 140562 332744
rect 154942 332732 154948 332744
rect 155000 332732 155006 332784
rect 129366 332664 129372 332716
rect 129424 332704 129430 332716
rect 154850 332704 154856 332716
rect 129424 332676 154856 332704
rect 129424 332664 129430 332676
rect 154850 332664 154856 332676
rect 154908 332664 154914 332716
rect 220630 332664 220636 332716
rect 220688 332704 220694 332716
rect 235626 332704 235632 332716
rect 220688 332676 235632 332704
rect 220688 332664 220694 332676
rect 235626 332664 235632 332676
rect 235684 332664 235690 332716
rect 220722 332596 220728 332648
rect 220780 332636 220786 332648
rect 244918 332636 244924 332648
rect 220780 332608 244924 332636
rect 220780 332596 220786 332608
rect 244918 332596 244924 332608
rect 244976 332596 244982 332648
rect 220446 331848 220452 331900
rect 220504 331888 220510 331900
rect 248138 331888 248144 331900
rect 220504 331860 248144 331888
rect 220504 331848 220510 331860
rect 248138 331848 248144 331860
rect 248196 331848 248202 331900
rect 219894 331576 219900 331628
rect 219952 331616 219958 331628
rect 227530 331616 227536 331628
rect 219952 331588 227536 331616
rect 219952 331576 219958 331588
rect 227530 331576 227536 331588
rect 227588 331576 227594 331628
rect 150066 331440 150072 331492
rect 150124 331480 150130 331492
rect 154942 331480 154948 331492
rect 150124 331452 154948 331480
rect 150124 331440 150130 331452
rect 154942 331440 154948 331452
rect 155000 331440 155006 331492
rect 219894 331440 219900 331492
rect 219952 331480 219958 331492
rect 224126 331480 224132 331492
rect 219952 331452 224132 331480
rect 219952 331440 219958 331452
rect 224126 331440 224132 331452
rect 224184 331440 224190 331492
rect 132126 331372 132132 331424
rect 132184 331412 132190 331424
rect 154850 331412 154856 331424
rect 132184 331384 154856 331412
rect 132184 331372 132190 331384
rect 154850 331372 154856 331384
rect 154908 331372 154914 331424
rect 129274 331304 129280 331356
rect 129332 331344 129338 331356
rect 154942 331344 154948 331356
rect 129332 331316 154948 331344
rect 129332 331304 129338 331316
rect 154942 331304 154948 331316
rect 155000 331304 155006 331356
rect 115750 331236 115756 331288
rect 115808 331276 115814 331288
rect 155034 331276 155040 331288
rect 115808 331248 155040 331276
rect 115808 331236 115814 331248
rect 155034 331236 155040 331248
rect 155092 331236 155098 331288
rect 220538 331236 220544 331288
rect 220596 331276 220602 331288
rect 254946 331276 254952 331288
rect 220596 331248 254952 331276
rect 220596 331236 220602 331248
rect 254946 331236 254952 331248
rect 255004 331236 255010 331288
rect 147398 330488 147404 330540
rect 147456 330528 147462 330540
rect 154758 330528 154764 330540
rect 147456 330500 154764 330528
rect 147456 330488 147462 330500
rect 154758 330488 154764 330500
rect 154816 330488 154822 330540
rect 144638 330012 144644 330064
rect 144696 330052 144702 330064
rect 154942 330052 154948 330064
rect 144696 330024 154948 330052
rect 144696 330012 144702 330024
rect 154942 330012 154948 330024
rect 155000 330012 155006 330064
rect 137646 329944 137652 329996
rect 137704 329984 137710 329996
rect 154850 329984 154856 329996
rect 137704 329956 154856 329984
rect 137704 329944 137710 329956
rect 154850 329944 154856 329956
rect 154908 329944 154914 329996
rect 219710 329944 219716 329996
rect 219768 329984 219774 329996
rect 228910 329984 228916 329996
rect 219768 329956 228916 329984
rect 219768 329944 219774 329956
rect 228910 329944 228916 329956
rect 228968 329944 228974 329996
rect 122558 329876 122564 329928
rect 122616 329916 122622 329928
rect 155034 329916 155040 329928
rect 122616 329888 155040 329916
rect 122616 329876 122622 329888
rect 155034 329876 155040 329888
rect 155092 329876 155098 329928
rect 220538 329876 220544 329928
rect 220596 329916 220602 329928
rect 231670 329916 231676 329928
rect 220596 329888 231676 329916
rect 220596 329876 220602 329888
rect 231670 329876 231676 329888
rect 231728 329876 231734 329928
rect 115658 329808 115664 329860
rect 115716 329848 115722 329860
rect 155126 329848 155132 329860
rect 115716 329820 155132 329848
rect 115716 329808 115722 329820
rect 155126 329808 155132 329820
rect 155184 329808 155190 329860
rect 220722 329808 220728 329860
rect 220780 329848 220786 329860
rect 250438 329848 250444 329860
rect 220780 329820 250444 329848
rect 220780 329808 220786 329820
rect 250438 329808 250444 329820
rect 250496 329808 250502 329860
rect 220630 329060 220636 329112
rect 220688 329100 220694 329112
rect 241238 329100 241244 329112
rect 220688 329072 241244 329100
rect 220688 329060 220694 329072
rect 241238 329060 241244 329072
rect 241296 329060 241302 329112
rect 219526 328992 219532 329044
rect 219584 329032 219590 329044
rect 224862 329032 224868 329044
rect 219584 329004 224868 329032
rect 219584 328992 219590 329004
rect 224862 328992 224868 329004
rect 224920 328992 224926 329044
rect 152918 328720 152924 328772
rect 152976 328760 152982 328772
rect 154574 328760 154580 328772
rect 152976 328732 154580 328760
rect 152976 328720 152982 328732
rect 154574 328720 154580 328732
rect 154632 328720 154638 328772
rect 149974 328652 149980 328704
rect 150032 328692 150038 328704
rect 154942 328692 154948 328704
rect 150032 328664 154948 328692
rect 150032 328652 150038 328664
rect 154942 328652 154948 328664
rect 155000 328652 155006 328704
rect 140406 328584 140412 328636
rect 140464 328624 140470 328636
rect 154850 328624 154856 328636
rect 140464 328596 154856 328624
rect 140464 328584 140470 328596
rect 154850 328584 154856 328596
rect 154908 328584 154914 328636
rect 132034 328516 132040 328568
rect 132092 328556 132098 328568
rect 154574 328556 154580 328568
rect 132092 328528 154580 328556
rect 132092 328516 132098 328528
rect 154574 328516 154580 328528
rect 154632 328516 154638 328568
rect 220722 328516 220728 328568
rect 220780 328556 220786 328568
rect 231578 328556 231584 328568
rect 220780 328528 231584 328556
rect 220780 328516 220786 328528
rect 231578 328516 231584 328528
rect 231636 328516 231642 328568
rect 112346 328448 112352 328500
rect 112404 328488 112410 328500
rect 155034 328488 155040 328500
rect 112404 328460 155040 328488
rect 112404 328448 112410 328460
rect 155034 328448 155040 328460
rect 155092 328448 155098 328500
rect 220538 328448 220544 328500
rect 220596 328488 220602 328500
rect 255958 328488 255964 328500
rect 220596 328460 255964 328488
rect 220596 328448 220602 328460
rect 255958 328448 255964 328460
rect 256016 328448 256022 328500
rect 220262 327904 220268 327956
rect 220320 327944 220326 327956
rect 228818 327944 228824 327956
rect 220320 327916 228824 327944
rect 220320 327904 220326 327916
rect 228818 327904 228824 327916
rect 228876 327904 228882 327956
rect 3418 327700 3424 327752
rect 3476 327740 3482 327752
rect 158254 327740 158260 327752
rect 3476 327712 158260 327740
rect 3476 327700 3482 327712
rect 158254 327700 158260 327712
rect 158312 327700 158318 327752
rect 227714 327700 227720 327752
rect 227772 327740 227778 327752
rect 257338 327740 257344 327752
rect 227772 327712 257344 327740
rect 227772 327700 227778 327712
rect 257338 327700 257344 327712
rect 257396 327700 257402 327752
rect 143258 327292 143264 327344
rect 143316 327332 143322 327344
rect 154758 327332 154764 327344
rect 143316 327304 154764 327332
rect 143316 327292 143322 327304
rect 154758 327292 154764 327304
rect 154816 327292 154822 327344
rect 121086 327224 121092 327276
rect 121144 327264 121150 327276
rect 154942 327264 154948 327276
rect 121144 327236 154948 327264
rect 121144 327224 121150 327236
rect 154942 327224 154948 327236
rect 155000 327224 155006 327276
rect 118050 327156 118056 327208
rect 118108 327196 118114 327208
rect 154850 327196 154856 327208
rect 118108 327168 154856 327196
rect 118108 327156 118114 327168
rect 154850 327156 154856 327168
rect 154908 327156 154914 327208
rect 220262 327156 220268 327208
rect 220320 327196 220326 327208
rect 226058 327196 226064 327208
rect 220320 327168 226064 327196
rect 220320 327156 220326 327168
rect 226058 327156 226064 327168
rect 226116 327156 226122 327208
rect 117038 327088 117044 327140
rect 117096 327128 117102 327140
rect 155034 327128 155040 327140
rect 117096 327100 155040 327128
rect 117096 327088 117102 327100
rect 155034 327088 155040 327100
rect 155092 327088 155098 327140
rect 220722 327088 220728 327140
rect 220780 327128 220786 327140
rect 238294 327128 238300 327140
rect 220780 327100 238300 327128
rect 220780 327088 220786 327100
rect 238294 327088 238300 327100
rect 238352 327088 238358 327140
rect 113082 325932 113088 325984
rect 113140 325972 113146 325984
rect 154850 325972 154856 325984
rect 113140 325944 154856 325972
rect 113140 325932 113146 325944
rect 154850 325932 154856 325944
rect 154908 325932 154914 325984
rect 137554 325864 137560 325916
rect 137612 325904 137618 325916
rect 154942 325904 154948 325916
rect 137612 325876 154948 325904
rect 137612 325864 137618 325876
rect 154942 325864 154948 325876
rect 155000 325864 155006 325916
rect 220354 325864 220360 325916
rect 220412 325904 220418 325916
rect 224770 325904 224776 325916
rect 220412 325876 224776 325904
rect 220412 325864 220418 325876
rect 224770 325864 224776 325876
rect 224828 325864 224834 325916
rect 131942 325796 131948 325848
rect 132000 325836 132006 325848
rect 154574 325836 154580 325848
rect 132000 325808 154580 325836
rect 132000 325796 132006 325808
rect 154574 325796 154580 325808
rect 154632 325796 154638 325848
rect 112990 325728 112996 325780
rect 113048 325768 113054 325780
rect 154758 325768 154764 325780
rect 113048 325740 154764 325768
rect 113048 325728 113054 325740
rect 154758 325728 154764 325740
rect 154816 325728 154822 325780
rect 220722 325728 220728 325780
rect 220780 325768 220786 325780
rect 228726 325768 228732 325780
rect 220780 325740 228732 325768
rect 220780 325728 220786 325740
rect 228726 325728 228732 325740
rect 228784 325728 228790 325780
rect 151354 325660 151360 325712
rect 151412 325700 151418 325712
rect 155034 325700 155040 325712
rect 151412 325672 155040 325700
rect 151412 325660 151418 325672
rect 155034 325660 155040 325672
rect 155092 325660 155098 325712
rect 220630 325660 220636 325712
rect 220688 325700 220694 325712
rect 236914 325700 236920 325712
rect 220688 325672 236920 325700
rect 220688 325660 220694 325672
rect 236914 325660 236920 325672
rect 236972 325660 236978 325712
rect 3510 324912 3516 324964
rect 3568 324952 3574 324964
rect 140038 324952 140044 324964
rect 3568 324924 140044 324952
rect 3568 324912 3574 324924
rect 140038 324912 140044 324924
rect 140096 324912 140102 324964
rect 219526 324912 219532 324964
rect 219584 324952 219590 324964
rect 234338 324952 234344 324964
rect 219584 324924 234344 324952
rect 219584 324912 219590 324924
rect 234338 324912 234344 324924
rect 234396 324912 234402 324964
rect 112898 324572 112904 324624
rect 112956 324612 112962 324624
rect 154942 324612 154948 324624
rect 112956 324584 154948 324612
rect 112956 324572 112962 324584
rect 154942 324572 154948 324584
rect 155000 324572 155006 324624
rect 220722 324572 220728 324624
rect 220780 324612 220786 324624
rect 220780 324584 229094 324612
rect 220780 324572 220786 324584
rect 123938 324504 123944 324556
rect 123996 324544 124002 324556
rect 155034 324544 155040 324556
rect 123996 324516 155040 324544
rect 123996 324504 124002 324516
rect 155034 324504 155040 324516
rect 155092 324504 155098 324556
rect 122466 324436 122472 324488
rect 122524 324476 122530 324488
rect 154850 324476 154856 324488
rect 122524 324448 154856 324476
rect 122524 324436 122530 324448
rect 154850 324436 154856 324448
rect 154908 324436 154914 324488
rect 220262 324436 220268 324488
rect 220320 324476 220326 324488
rect 225966 324476 225972 324488
rect 220320 324448 225972 324476
rect 220320 324436 220326 324448
rect 225966 324436 225972 324448
rect 226024 324436 226030 324488
rect 120994 324368 121000 324420
rect 121052 324408 121058 324420
rect 154758 324408 154764 324420
rect 121052 324380 154764 324408
rect 121052 324368 121058 324380
rect 154758 324368 154764 324380
rect 154816 324368 154822 324420
rect 220354 324368 220360 324420
rect 220412 324408 220418 324420
rect 229066 324408 229094 324584
rect 235534 324408 235540 324420
rect 220412 324380 224816 324408
rect 229066 324380 235540 324408
rect 220412 324368 220418 324380
rect 149882 324300 149888 324352
rect 149940 324340 149946 324352
rect 154942 324340 154948 324352
rect 149940 324312 154948 324340
rect 149940 324300 149946 324312
rect 154942 324300 154948 324312
rect 155000 324300 155006 324352
rect 219894 324300 219900 324352
rect 219952 324340 219958 324352
rect 224678 324340 224684 324352
rect 219952 324312 224684 324340
rect 219952 324300 219958 324312
rect 224678 324300 224684 324312
rect 224736 324300 224742 324352
rect 224788 324340 224816 324380
rect 235534 324368 235540 324380
rect 235592 324368 235598 324420
rect 580166 324340 580172 324352
rect 224788 324312 580172 324340
rect 580166 324300 580172 324312
rect 580224 324300 580230 324352
rect 3602 323552 3608 323604
rect 3660 323592 3666 323604
rect 157886 323592 157892 323604
rect 3660 323564 157892 323592
rect 3660 323552 3666 323564
rect 157886 323552 157892 323564
rect 157944 323552 157950 323604
rect 219710 323280 219716 323332
rect 219768 323320 219774 323332
rect 228634 323320 228640 323332
rect 219768 323292 228640 323320
rect 219768 323280 219774 323292
rect 228634 323280 228640 323292
rect 228692 323280 228698 323332
rect 112806 323212 112812 323264
rect 112864 323252 112870 323264
rect 154942 323252 154948 323264
rect 112864 323224 154948 323252
rect 112864 323212 112870 323224
rect 154942 323212 154948 323224
rect 155000 323212 155006 323264
rect 137462 323144 137468 323196
rect 137520 323184 137526 323196
rect 155034 323184 155040 323196
rect 137520 323156 155040 323184
rect 137520 323144 137526 323156
rect 155034 323144 155040 323156
rect 155092 323144 155098 323196
rect 130838 323076 130844 323128
rect 130896 323116 130902 323128
rect 154942 323116 154948 323128
rect 130896 323088 154948 323116
rect 130896 323076 130902 323088
rect 154942 323076 154948 323088
rect 155000 323076 155006 323128
rect 220262 323076 220268 323128
rect 220320 323116 220326 323128
rect 224586 323116 224592 323128
rect 220320 323088 224592 323116
rect 220320 323076 220326 323088
rect 224586 323076 224592 323088
rect 224644 323076 224650 323128
rect 114370 323008 114376 323060
rect 114428 323048 114434 323060
rect 154850 323048 154856 323060
rect 114428 323020 154856 323048
rect 114428 323008 114434 323020
rect 154850 323008 154856 323020
rect 154908 323008 154914 323060
rect 220722 323008 220728 323060
rect 220780 323048 220786 323060
rect 224034 323048 224040 323060
rect 220780 323020 224040 323048
rect 220780 323008 220786 323020
rect 224034 323008 224040 323020
rect 224092 323008 224098 323060
rect 220630 322940 220636 322992
rect 220688 322980 220694 322992
rect 231486 322980 231492 322992
rect 220688 322952 231492 322980
rect 220688 322940 220694 322952
rect 231486 322940 231492 322952
rect 231544 322940 231550 322992
rect 3786 322260 3792 322312
rect 3844 322300 3850 322312
rect 142890 322300 142896 322312
rect 3844 322272 142896 322300
rect 3844 322260 3850 322272
rect 142890 322260 142896 322272
rect 142948 322260 142954 322312
rect 3694 322192 3700 322244
rect 3752 322232 3758 322244
rect 152550 322232 152556 322244
rect 3752 322204 152556 322232
rect 3752 322192 3758 322204
rect 152550 322192 152556 322204
rect 152608 322192 152614 322244
rect 147306 321784 147312 321836
rect 147364 321824 147370 321836
rect 154850 321824 154856 321836
rect 147364 321796 154856 321824
rect 147364 321784 147370 321796
rect 154850 321784 154856 321796
rect 154908 321784 154914 321836
rect 126698 321716 126704 321768
rect 126756 321756 126762 321768
rect 155034 321756 155040 321768
rect 126756 321728 155040 321756
rect 126756 321716 126762 321728
rect 155034 321716 155040 321728
rect 155092 321716 155098 321768
rect 220538 321716 220544 321768
rect 220596 321756 220602 321768
rect 236822 321756 236828 321768
rect 220596 321728 236828 321756
rect 220596 321716 220602 321728
rect 236822 321716 236828 321728
rect 236880 321716 236886 321768
rect 116946 321648 116952 321700
rect 117004 321688 117010 321700
rect 154942 321688 154948 321700
rect 117004 321660 154948 321688
rect 117004 321648 117010 321660
rect 154942 321648 154948 321660
rect 155000 321648 155006 321700
rect 220722 321648 220728 321700
rect 220780 321688 220786 321700
rect 250714 321688 250720 321700
rect 220780 321660 250720 321688
rect 220780 321648 220786 321660
rect 250714 321648 250720 321660
rect 250772 321648 250778 321700
rect 115566 321580 115572 321632
rect 115624 321620 115630 321632
rect 154758 321620 154764 321632
rect 115624 321592 154764 321620
rect 115624 321580 115630 321592
rect 154758 321580 154764 321592
rect 154816 321580 154822 321632
rect 220630 321580 220636 321632
rect 220688 321620 220694 321632
rect 256326 321620 256332 321632
rect 220688 321592 256332 321620
rect 220688 321580 220694 321592
rect 256326 321580 256332 321592
rect 256384 321580 256390 321632
rect 228358 320900 228364 320952
rect 228416 320940 228422 320952
rect 580902 320940 580908 320952
rect 228416 320912 580908 320940
rect 228416 320900 228422 320912
rect 580902 320900 580908 320912
rect 580960 320900 580966 320952
rect 218974 320832 218980 320884
rect 219032 320872 219038 320884
rect 580718 320872 580724 320884
rect 219032 320844 580724 320872
rect 219032 320832 219038 320844
rect 580718 320832 580724 320844
rect 580776 320832 580782 320884
rect 220262 320560 220268 320612
rect 220320 320600 220326 320612
rect 222746 320600 222752 320612
rect 220320 320572 222752 320600
rect 220320 320560 220326 320572
rect 222746 320560 222752 320572
rect 222804 320560 222810 320612
rect 144454 320424 144460 320476
rect 144512 320464 144518 320476
rect 154942 320464 154948 320476
rect 144512 320436 154948 320464
rect 144512 320424 144518 320436
rect 154942 320424 154948 320436
rect 155000 320424 155006 320476
rect 143166 320356 143172 320408
rect 143224 320396 143230 320408
rect 154850 320396 154856 320408
rect 143224 320368 154856 320396
rect 143224 320356 143230 320368
rect 154850 320356 154856 320368
rect 154908 320356 154914 320408
rect 133414 320288 133420 320340
rect 133472 320328 133478 320340
rect 154758 320328 154764 320340
rect 133472 320300 154764 320328
rect 133472 320288 133478 320300
rect 154758 320288 154764 320300
rect 154816 320288 154822 320340
rect 133322 320220 133328 320272
rect 133380 320260 133386 320272
rect 154942 320260 154948 320272
rect 133380 320232 154948 320260
rect 133380 320220 133386 320232
rect 154942 320220 154948 320232
rect 155000 320220 155006 320272
rect 220262 320220 220268 320272
rect 220320 320260 220326 320272
rect 242342 320260 242348 320272
rect 220320 320232 242348 320260
rect 220320 320220 220326 320232
rect 242342 320220 242348 320232
rect 242400 320220 242406 320272
rect 112714 320152 112720 320204
rect 112772 320192 112778 320204
rect 155034 320192 155040 320204
rect 112772 320164 155040 320192
rect 112772 320152 112778 320164
rect 155034 320152 155040 320164
rect 155092 320152 155098 320204
rect 220722 320152 220728 320204
rect 220780 320192 220786 320204
rect 249518 320192 249524 320204
rect 220780 320164 249524 320192
rect 220780 320152 220786 320164
rect 249518 320152 249524 320164
rect 249576 320152 249582 320204
rect 220170 320016 220176 320068
rect 220228 320056 220234 320068
rect 220228 320028 220308 320056
rect 220228 320016 220234 320028
rect 220280 319864 220308 320028
rect 220262 319812 220268 319864
rect 220320 319812 220326 319864
rect 220446 319744 220452 319796
rect 220504 319784 220510 319796
rect 223482 319784 223488 319796
rect 220504 319756 223488 319784
rect 220504 319744 220510 319756
rect 223482 319744 223488 319756
rect 223540 319744 223546 319796
rect 229922 319676 229928 319728
rect 229980 319716 229986 319728
rect 580350 319716 580356 319728
rect 229980 319688 580356 319716
rect 229980 319676 229986 319688
rect 580350 319676 580356 319688
rect 580408 319676 580414 319728
rect 229738 319608 229744 319660
rect 229796 319648 229802 319660
rect 580258 319648 580264 319660
rect 229796 319620 580264 319648
rect 229796 319608 229802 319620
rect 580258 319608 580264 319620
rect 580316 319608 580322 319660
rect 226978 319540 226984 319592
rect 227036 319580 227042 319592
rect 580534 319580 580540 319592
rect 227036 319552 580540 319580
rect 227036 319540 227042 319552
rect 580534 319540 580540 319552
rect 580592 319540 580598 319592
rect 221642 319472 221648 319524
rect 221700 319512 221706 319524
rect 580810 319512 580816 319524
rect 221700 319484 580816 319512
rect 221700 319472 221706 319484
rect 580810 319472 580816 319484
rect 580868 319472 580874 319524
rect 118142 319404 118148 319456
rect 118200 319444 118206 319456
rect 154666 319444 154672 319456
rect 118200 319416 154672 319444
rect 118200 319404 118206 319416
rect 154666 319404 154672 319416
rect 154724 319404 154730 319456
rect 219158 319404 219164 319456
rect 219216 319444 219222 319456
rect 580626 319444 580632 319456
rect 219216 319416 580632 319444
rect 219216 319404 219222 319416
rect 580626 319404 580632 319416
rect 580684 319404 580690 319456
rect 148686 318996 148692 319048
rect 148744 319036 148750 319048
rect 154850 319036 154856 319048
rect 148744 319008 154856 319036
rect 148744 318996 148750 319008
rect 154850 318996 154856 319008
rect 154908 318996 154914 319048
rect 220722 318996 220728 319048
rect 220780 319036 220786 319048
rect 252002 319036 252008 319048
rect 220780 319008 252008 319036
rect 220780 318996 220786 319008
rect 252002 318996 252008 319008
rect 252060 318996 252066 319048
rect 130746 318928 130752 318980
rect 130804 318968 130810 318980
rect 154758 318968 154764 318980
rect 130804 318940 154764 318968
rect 130804 318928 130810 318940
rect 154758 318928 154764 318940
rect 154816 318928 154822 318980
rect 127986 318860 127992 318912
rect 128044 318900 128050 318912
rect 154942 318900 154948 318912
rect 128044 318872 154948 318900
rect 128044 318860 128050 318872
rect 154942 318860 154948 318872
rect 155000 318860 155006 318912
rect 220446 318860 220452 318912
rect 220504 318900 220510 318912
rect 223390 318900 223396 318912
rect 220504 318872 223396 318900
rect 220504 318860 220510 318872
rect 223390 318860 223396 318872
rect 223448 318860 223454 318912
rect 3418 318792 3424 318844
rect 3476 318832 3482 318844
rect 30006 318832 30012 318844
rect 3476 318804 30012 318832
rect 3476 318792 3482 318804
rect 30006 318792 30012 318804
rect 30064 318792 30070 318844
rect 114278 318792 114284 318844
rect 114336 318832 114342 318844
rect 155034 318832 155040 318844
rect 114336 318804 155040 318832
rect 114336 318792 114342 318804
rect 155034 318792 155040 318804
rect 155092 318792 155098 318844
rect 220354 318792 220360 318844
rect 220412 318832 220418 318844
rect 223298 318832 223304 318844
rect 220412 318804 223304 318832
rect 220412 318792 220418 318804
rect 223298 318792 223304 318804
rect 223356 318792 223362 318844
rect 254578 318792 254584 318844
rect 254636 318832 254642 318844
rect 580442 318832 580448 318844
rect 254636 318804 580448 318832
rect 254636 318792 254642 318804
rect 580442 318792 580448 318804
rect 580500 318792 580506 318844
rect 219986 318384 219992 318436
rect 220044 318424 220050 318436
rect 221826 318424 221832 318436
rect 220044 318396 221832 318424
rect 220044 318384 220050 318396
rect 221826 318384 221832 318396
rect 221884 318384 221890 318436
rect 122374 318044 122380 318096
rect 122432 318084 122438 318096
rect 154574 318084 154580 318096
rect 122432 318056 154580 318084
rect 122432 318044 122438 318056
rect 154574 318044 154580 318056
rect 154632 318044 154638 318096
rect 148594 317704 148600 317756
rect 148652 317744 148658 317756
rect 154850 317744 154856 317756
rect 148652 317716 154856 317744
rect 148652 317704 148658 317716
rect 154850 317704 154856 317716
rect 154908 317704 154914 317756
rect 145650 317636 145656 317688
rect 145708 317676 145714 317688
rect 154942 317676 154948 317688
rect 145708 317648 154948 317676
rect 145708 317636 145714 317648
rect 154942 317636 154948 317648
rect 155000 317636 155006 317688
rect 139026 317568 139032 317620
rect 139084 317608 139090 317620
rect 155034 317608 155040 317620
rect 139084 317580 155040 317608
rect 139084 317568 139090 317580
rect 155034 317568 155040 317580
rect 155092 317568 155098 317620
rect 122282 317500 122288 317552
rect 122340 317540 122346 317552
rect 154758 317540 154764 317552
rect 122340 317512 154764 317540
rect 122340 317500 122346 317512
rect 154758 317500 154764 317512
rect 154816 317500 154822 317552
rect 220630 317500 220636 317552
rect 220688 317540 220694 317552
rect 239674 317540 239680 317552
rect 220688 317512 239680 317540
rect 220688 317500 220694 317512
rect 239674 317500 239680 317512
rect 239732 317500 239738 317552
rect 119706 317432 119712 317484
rect 119764 317472 119770 317484
rect 154666 317472 154672 317484
rect 119764 317444 154672 317472
rect 119764 317432 119770 317444
rect 154666 317432 154672 317444
rect 154724 317432 154730 317484
rect 220722 317432 220728 317484
rect 220780 317472 220786 317484
rect 256234 317472 256240 317484
rect 220780 317444 256240 317472
rect 220780 317432 220786 317444
rect 256234 317432 256240 317444
rect 256292 317432 256298 317484
rect 220630 316480 220636 316532
rect 220688 316520 220694 316532
rect 225874 316520 225880 316532
rect 220688 316492 225880 316520
rect 220688 316480 220694 316492
rect 225874 316480 225880 316492
rect 225932 316480 225938 316532
rect 152826 316344 152832 316396
rect 152884 316384 152890 316396
rect 154574 316384 154580 316396
rect 152884 316356 154580 316384
rect 152884 316344 152890 316356
rect 154574 316344 154580 316356
rect 154632 316344 154638 316396
rect 115474 316276 115480 316328
rect 115532 316316 115538 316328
rect 154850 316316 154856 316328
rect 115532 316288 154856 316316
rect 115532 316276 115538 316288
rect 154850 316276 154856 316288
rect 154908 316276 154914 316328
rect 147214 316208 147220 316260
rect 147272 316248 147278 316260
rect 154758 316248 154764 316260
rect 147272 316220 154764 316248
rect 147272 316208 147278 316220
rect 154758 316208 154764 316220
rect 154816 316208 154822 316260
rect 130654 316140 130660 316192
rect 130712 316180 130718 316192
rect 155034 316180 155040 316192
rect 130712 316152 155040 316180
rect 130712 316140 130718 316152
rect 155034 316140 155040 316152
rect 155092 316140 155098 316192
rect 126606 316072 126612 316124
rect 126664 316112 126670 316124
rect 154942 316112 154948 316124
rect 126664 316084 154948 316112
rect 126664 316072 126670 316084
rect 154942 316072 154948 316084
rect 155000 316072 155006 316124
rect 220446 316072 220452 316124
rect 220504 316112 220510 316124
rect 248046 316112 248052 316124
rect 220504 316084 248052 316112
rect 220504 316072 220510 316084
rect 248046 316072 248052 316084
rect 248104 316072 248110 316124
rect 220722 316004 220728 316056
rect 220780 316044 220786 316056
rect 254854 316044 254860 316056
rect 220780 316016 254860 316044
rect 220780 316004 220786 316016
rect 254854 316004 254860 316016
rect 254912 316004 254918 316056
rect 127894 314848 127900 314900
rect 127952 314888 127958 314900
rect 155034 314888 155040 314900
rect 127952 314860 155040 314888
rect 127952 314848 127958 314860
rect 155034 314848 155040 314860
rect 155092 314848 155098 314900
rect 219986 314848 219992 314900
rect 220044 314888 220050 314900
rect 227346 314888 227352 314900
rect 220044 314860 227352 314888
rect 220044 314848 220050 314860
rect 227346 314848 227352 314860
rect 227404 314848 227410 314900
rect 125042 314780 125048 314832
rect 125100 314820 125106 314832
rect 154850 314820 154856 314832
rect 125100 314792 154856 314820
rect 125100 314780 125106 314792
rect 154850 314780 154856 314792
rect 154908 314780 154914 314832
rect 220538 314780 220544 314832
rect 220596 314820 220602 314832
rect 223206 314820 223212 314832
rect 220596 314792 223212 314820
rect 220596 314780 220602 314792
rect 223206 314780 223212 314792
rect 223264 314780 223270 314832
rect 123846 314712 123852 314764
rect 123904 314752 123910 314764
rect 154758 314752 154764 314764
rect 123904 314724 154764 314752
rect 123904 314712 123910 314724
rect 154758 314712 154764 314724
rect 154816 314712 154822 314764
rect 220630 314712 220636 314764
rect 220688 314752 220694 314764
rect 230198 314752 230204 314764
rect 220688 314724 230204 314752
rect 220688 314712 220694 314724
rect 230198 314712 230204 314724
rect 230256 314712 230262 314764
rect 122190 314644 122196 314696
rect 122248 314684 122254 314696
rect 154942 314684 154948 314696
rect 122248 314656 154948 314684
rect 122248 314644 122254 314656
rect 154942 314644 154948 314656
rect 155000 314644 155006 314696
rect 220722 314644 220728 314696
rect 220780 314684 220786 314696
rect 243906 314684 243912 314696
rect 220780 314656 243912 314684
rect 220780 314644 220786 314656
rect 243906 314644 243912 314656
rect 243964 314644 243970 314696
rect 111794 314576 111800 314628
rect 111852 314616 111858 314628
rect 138750 314616 138756 314628
rect 111852 314588 138756 314616
rect 111852 314576 111858 314588
rect 138750 314576 138756 314588
rect 138808 314576 138814 314628
rect 147122 313556 147128 313608
rect 147180 313596 147186 313608
rect 154942 313596 154948 313608
rect 147180 313568 154948 313596
rect 147180 313556 147186 313568
rect 154942 313556 154948 313568
rect 155000 313556 155006 313608
rect 134610 313488 134616 313540
rect 134668 313528 134674 313540
rect 154574 313528 154580 313540
rect 134668 313500 154580 313528
rect 134668 313488 134674 313500
rect 154574 313488 154580 313500
rect 154632 313488 154638 313540
rect 130562 313420 130568 313472
rect 130620 313460 130626 313472
rect 154942 313460 154948 313472
rect 130620 313432 154948 313460
rect 130620 313420 130626 313432
rect 154942 313420 154948 313432
rect 155000 313420 155006 313472
rect 220722 313420 220728 313472
rect 220780 313460 220786 313472
rect 230106 313460 230112 313472
rect 220780 313432 230112 313460
rect 220780 313420 220786 313432
rect 230106 313420 230112 313432
rect 230164 313420 230170 313472
rect 115382 313352 115388 313404
rect 115440 313392 115446 313404
rect 154850 313392 154856 313404
rect 115440 313364 154856 313392
rect 115440 313352 115446 313364
rect 154850 313352 154856 313364
rect 154908 313352 154914 313404
rect 220446 313352 220452 313404
rect 220504 313392 220510 313404
rect 239582 313392 239588 313404
rect 220504 313364 239588 313392
rect 220504 313352 220510 313364
rect 239582 313352 239588 313364
rect 239640 313352 239646 313404
rect 112622 313284 112628 313336
rect 112680 313324 112686 313336
rect 154758 313324 154764 313336
rect 112680 313296 154764 313324
rect 112680 313284 112686 313296
rect 154758 313284 154764 313296
rect 154816 313284 154822 313336
rect 220630 313284 220636 313336
rect 220688 313324 220694 313336
rect 249426 313324 249432 313336
rect 220688 313296 249432 313324
rect 220688 313284 220694 313296
rect 249426 313284 249432 313296
rect 249484 313284 249490 313336
rect 111794 313216 111800 313268
rect 111852 313256 111858 313268
rect 126238 313256 126244 313268
rect 111852 313228 126244 313256
rect 111852 313216 111858 313228
rect 126238 313216 126244 313228
rect 126296 313216 126302 313268
rect 111886 313148 111892 313200
rect 111944 313188 111950 313200
rect 117958 313188 117964 313200
rect 111944 313160 117964 313188
rect 111944 313148 111950 313160
rect 117958 313148 117964 313160
rect 118016 313148 118022 313200
rect 227070 312536 227076 312588
rect 227128 312576 227134 312588
rect 257706 312576 257712 312588
rect 227128 312548 257712 312576
rect 227128 312536 227134 312548
rect 257706 312536 257712 312548
rect 257764 312536 257770 312588
rect 220446 312400 220452 312452
rect 220504 312440 220510 312452
rect 224494 312440 224500 312452
rect 220504 312412 224500 312440
rect 220504 312400 220510 312412
rect 224494 312400 224500 312412
rect 224552 312400 224558 312452
rect 219894 312196 219900 312248
rect 219952 312236 219958 312248
rect 227254 312236 227260 312248
rect 219952 312208 227260 312236
rect 219952 312196 219958 312208
rect 227254 312196 227260 312208
rect 227312 312196 227318 312248
rect 123754 312128 123760 312180
rect 123812 312168 123818 312180
rect 154942 312168 154948 312180
rect 123812 312140 154948 312168
rect 123812 312128 123818 312140
rect 154942 312128 154948 312140
rect 155000 312128 155006 312180
rect 133138 312060 133144 312112
rect 133196 312100 133202 312112
rect 154574 312100 154580 312112
rect 133196 312072 154580 312100
rect 133196 312060 133202 312072
rect 154574 312060 154580 312072
rect 154632 312060 154638 312112
rect 127802 311992 127808 312044
rect 127860 312032 127866 312044
rect 154758 312032 154764 312044
rect 127860 312004 154764 312032
rect 127860 311992 127866 312004
rect 154758 311992 154764 312004
rect 154816 311992 154822 312044
rect 126514 311924 126520 311976
rect 126572 311964 126578 311976
rect 154850 311964 154856 311976
rect 126572 311936 154856 311964
rect 126572 311924 126578 311936
rect 154850 311924 154856 311936
rect 154908 311924 154914 311976
rect 220722 311924 220728 311976
rect 220780 311964 220786 311976
rect 225782 311964 225788 311976
rect 220780 311936 225788 311964
rect 220780 311924 220786 311936
rect 225782 311924 225788 311936
rect 225840 311924 225846 311976
rect 152734 311856 152740 311908
rect 152792 311896 152798 311908
rect 154574 311896 154580 311908
rect 152792 311868 154580 311896
rect 152792 311856 152798 311868
rect 154574 311856 154580 311868
rect 154632 311856 154638 311908
rect 220446 311856 220452 311908
rect 220504 311896 220510 311908
rect 235442 311896 235448 311908
rect 220504 311868 235448 311896
rect 220504 311856 220510 311868
rect 235442 311856 235448 311868
rect 235500 311856 235506 311908
rect 111886 311788 111892 311840
rect 111944 311828 111950 311840
rect 122650 311828 122656 311840
rect 111944 311800 122656 311828
rect 111944 311788 111950 311800
rect 122650 311788 122656 311800
rect 122708 311788 122714 311840
rect 229830 311788 229836 311840
rect 229888 311828 229894 311840
rect 256694 311828 256700 311840
rect 229888 311800 256700 311828
rect 229888 311788 229894 311800
rect 256694 311788 256700 311800
rect 256752 311788 256758 311840
rect 111794 311720 111800 311772
rect 111852 311760 111858 311772
rect 116670 311760 116676 311772
rect 111852 311732 116676 311760
rect 111852 311720 111858 311732
rect 116670 311720 116676 311732
rect 116728 311720 116734 311772
rect 154666 311176 154672 311228
rect 154724 311216 154730 311228
rect 155402 311216 155408 311228
rect 154724 311188 155408 311216
rect 154724 311176 154730 311188
rect 155402 311176 155408 311188
rect 155460 311176 155466 311228
rect 116854 311108 116860 311160
rect 116912 311148 116918 311160
rect 155586 311148 155592 311160
rect 116912 311120 155592 311148
rect 116912 311108 116918 311120
rect 155586 311108 155592 311120
rect 155644 311108 155650 311160
rect 114186 310768 114192 310820
rect 114244 310808 114250 310820
rect 154850 310808 154856 310820
rect 114244 310780 154856 310808
rect 114244 310768 114250 310780
rect 154850 310768 154856 310780
rect 154908 310768 154914 310820
rect 145742 310700 145748 310752
rect 145800 310740 145806 310752
rect 154942 310740 154948 310752
rect 145800 310712 154948 310740
rect 145800 310700 145806 310712
rect 154942 310700 154948 310712
rect 155000 310700 155006 310752
rect 138934 310632 138940 310684
rect 138992 310672 138998 310684
rect 154850 310672 154856 310684
rect 138992 310644 154856 310672
rect 138992 310632 138998 310644
rect 154850 310632 154856 310644
rect 154908 310632 154914 310684
rect 220538 310632 220544 310684
rect 220596 310672 220602 310684
rect 227438 310672 227444 310684
rect 220596 310644 227444 310672
rect 220596 310632 220602 310644
rect 227438 310632 227444 310644
rect 227496 310632 227502 310684
rect 119614 310564 119620 310616
rect 119672 310604 119678 310616
rect 154758 310604 154764 310616
rect 119672 310576 154764 310604
rect 119672 310564 119678 310576
rect 154758 310564 154764 310576
rect 154816 310564 154822 310616
rect 220722 310564 220728 310616
rect 220780 310604 220786 310616
rect 230014 310604 230020 310616
rect 220780 310576 230020 310604
rect 220780 310564 220786 310576
rect 230014 310564 230020 310576
rect 230072 310564 230078 310616
rect 151262 310496 151268 310548
rect 151320 310536 151326 310548
rect 155034 310536 155040 310548
rect 151320 310508 155040 310536
rect 151320 310496 151326 310508
rect 155034 310496 155040 310508
rect 155092 310496 155098 310548
rect 220630 310496 220636 310548
rect 220688 310536 220694 310548
rect 245102 310536 245108 310548
rect 220688 310508 245108 310536
rect 220688 310496 220694 310508
rect 245102 310496 245108 310508
rect 245160 310496 245166 310548
rect 111794 310428 111800 310480
rect 111852 310468 111858 310480
rect 119522 310468 119528 310480
rect 111852 310440 119528 310468
rect 111852 310428 111858 310440
rect 119522 310428 119528 310440
rect 119580 310428 119586 310480
rect 111886 310360 111892 310412
rect 111944 310400 111950 310412
rect 119430 310400 119436 310412
rect 111944 310372 119436 310400
rect 111944 310360 111950 310372
rect 119430 310360 119436 310372
rect 119488 310360 119494 310412
rect 233970 309748 233976 309800
rect 234028 309788 234034 309800
rect 256786 309788 256792 309800
rect 234028 309760 256792 309788
rect 234028 309748 234034 309760
rect 256786 309748 256792 309760
rect 256844 309748 256850 309800
rect 144362 309408 144368 309460
rect 144420 309448 144426 309460
rect 154850 309448 154856 309460
rect 144420 309420 154856 309448
rect 144420 309408 144426 309420
rect 154850 309408 154856 309420
rect 154908 309408 154914 309460
rect 220630 309408 220636 309460
rect 220688 309448 220694 309460
rect 224402 309448 224408 309460
rect 220688 309420 224408 309448
rect 220688 309408 220694 309420
rect 224402 309408 224408 309420
rect 224460 309408 224466 309460
rect 130470 309340 130476 309392
rect 130528 309380 130534 309392
rect 154758 309380 154764 309392
rect 130528 309352 154764 309380
rect 130528 309340 130534 309352
rect 154758 309340 154764 309352
rect 154816 309340 154822 309392
rect 127710 309272 127716 309324
rect 127768 309312 127774 309324
rect 154942 309312 154948 309324
rect 127768 309284 154948 309312
rect 127768 309272 127774 309284
rect 154942 309272 154948 309284
rect 155000 309272 155006 309324
rect 126422 309204 126428 309256
rect 126480 309244 126486 309256
rect 154574 309244 154580 309256
rect 126480 309216 154580 309244
rect 126480 309204 126486 309216
rect 154574 309204 154580 309216
rect 154632 309204 154638 309256
rect 220538 309204 220544 309256
rect 220596 309244 220602 309256
rect 234246 309244 234252 309256
rect 220596 309216 234252 309244
rect 220596 309204 220602 309216
rect 234246 309204 234252 309216
rect 234304 309204 234310 309256
rect 124950 309136 124956 309188
rect 125008 309176 125014 309188
rect 154942 309176 154948 309188
rect 125008 309148 154948 309176
rect 125008 309136 125014 309148
rect 154942 309136 154948 309148
rect 155000 309136 155006 309188
rect 220722 309136 220728 309188
rect 220780 309176 220786 309188
rect 246758 309176 246764 309188
rect 220780 309148 246764 309176
rect 220780 309136 220786 309148
rect 246758 309136 246764 309148
rect 246816 309136 246822 309188
rect 111794 309068 111800 309120
rect 111852 309108 111858 309120
rect 118234 309108 118240 309120
rect 111852 309080 118240 309108
rect 111852 309068 111858 309080
rect 118234 309068 118240 309080
rect 118292 309068 118298 309120
rect 247770 309068 247776 309120
rect 247828 309108 247834 309120
rect 256694 309108 256700 309120
rect 247828 309080 256700 309108
rect 247828 309068 247834 309080
rect 256694 309068 256700 309080
rect 256752 309068 256758 309120
rect 111886 309000 111892 309052
rect 111944 309040 111950 309052
rect 116578 309040 116584 309052
rect 111944 309012 116584 309040
rect 111944 309000 111950 309012
rect 116578 309000 116584 309012
rect 116636 309000 116642 309052
rect 149790 307980 149796 308032
rect 149848 308020 149854 308032
rect 154942 308020 154948 308032
rect 149848 307992 154948 308020
rect 149848 307980 149854 307992
rect 154942 307980 154948 307992
rect 155000 307980 155006 308032
rect 219894 307980 219900 308032
rect 219952 308020 219958 308032
rect 225690 308020 225696 308032
rect 219952 307992 225696 308020
rect 219952 307980 219958 307992
rect 225690 307980 225696 307992
rect 225748 307980 225754 308032
rect 141694 307912 141700 307964
rect 141752 307952 141758 307964
rect 154758 307952 154764 307964
rect 141752 307924 154764 307952
rect 141752 307912 141758 307924
rect 154758 307912 154764 307924
rect 154816 307912 154822 307964
rect 220722 307912 220728 307964
rect 220780 307952 220786 307964
rect 232682 307952 232688 307964
rect 220780 307924 232688 307952
rect 220780 307912 220786 307924
rect 232682 307912 232688 307924
rect 232740 307912 232746 307964
rect 123570 307844 123576 307896
rect 123628 307884 123634 307896
rect 155034 307884 155040 307896
rect 123628 307856 155040 307884
rect 123628 307844 123634 307856
rect 155034 307844 155040 307856
rect 155092 307844 155098 307896
rect 220630 307844 220636 307896
rect 220688 307884 220694 307896
rect 238202 307884 238208 307896
rect 220688 307856 238208 307884
rect 220688 307844 220694 307856
rect 238202 307844 238208 307856
rect 238260 307844 238266 307896
rect 117958 307776 117964 307828
rect 118016 307816 118022 307828
rect 154850 307816 154856 307828
rect 118016 307788 154856 307816
rect 118016 307776 118022 307788
rect 154850 307776 154856 307788
rect 154908 307776 154914 307828
rect 219710 307776 219716 307828
rect 219768 307816 219774 307828
rect 242250 307816 242256 307828
rect 219768 307788 242256 307816
rect 219768 307776 219774 307788
rect 242250 307776 242256 307788
rect 242308 307776 242314 307828
rect 111794 307708 111800 307760
rect 111852 307748 111858 307760
rect 142982 307748 142988 307760
rect 111852 307720 142988 307748
rect 111852 307708 111858 307720
rect 142982 307708 142988 307720
rect 143040 307708 143046 307760
rect 111794 307504 111800 307556
rect 111852 307544 111858 307556
rect 113910 307544 113916 307556
rect 111852 307516 113916 307544
rect 111852 307504 111858 307516
rect 113910 307504 113916 307516
rect 113968 307504 113974 307556
rect 148502 306620 148508 306672
rect 148560 306660 148566 306672
rect 155034 306660 155040 306672
rect 148560 306632 155040 306660
rect 148560 306620 148566 306632
rect 155034 306620 155040 306632
rect 155092 306620 155098 306672
rect 143074 306552 143080 306604
rect 143132 306592 143138 306604
rect 154942 306592 154948 306604
rect 143132 306564 154948 306592
rect 143132 306552 143138 306564
rect 154942 306552 154948 306564
rect 155000 306552 155006 306604
rect 130378 306484 130384 306536
rect 130436 306524 130442 306536
rect 154850 306524 154856 306536
rect 130436 306496 154856 306524
rect 130436 306484 130442 306496
rect 154850 306484 154856 306496
rect 154908 306484 154914 306536
rect 155034 306484 155040 306536
rect 155092 306524 155098 306536
rect 155678 306524 155684 306536
rect 155092 306496 155684 306524
rect 155092 306484 155098 306496
rect 155678 306484 155684 306496
rect 155736 306484 155742 306536
rect 220538 306484 220544 306536
rect 220596 306524 220602 306536
rect 232866 306524 232872 306536
rect 220596 306496 232872 306524
rect 220596 306484 220602 306496
rect 232866 306484 232872 306496
rect 232924 306484 232930 306536
rect 126330 306416 126336 306468
rect 126388 306456 126394 306468
rect 154942 306456 154948 306468
rect 126388 306428 154948 306456
rect 126388 306416 126394 306428
rect 154942 306416 154948 306428
rect 155000 306416 155006 306468
rect 155310 306416 155316 306468
rect 155368 306416 155374 306468
rect 220722 306416 220728 306468
rect 220780 306456 220786 306468
rect 238110 306456 238116 306468
rect 220780 306428 238116 306456
rect 220780 306416 220786 306428
rect 238110 306416 238116 306428
rect 238168 306416 238174 306468
rect 112070 306348 112076 306400
rect 112128 306388 112134 306400
rect 154758 306388 154764 306400
rect 112128 306360 154764 306388
rect 112128 306348 112134 306360
rect 154758 306348 154764 306360
rect 154816 306348 154822 306400
rect 154850 306348 154856 306400
rect 154908 306388 154914 306400
rect 155328 306388 155356 306416
rect 154908 306360 155356 306388
rect 154908 306348 154914 306360
rect 220630 306348 220636 306400
rect 220688 306388 220694 306400
rect 247954 306388 247960 306400
rect 220688 306360 247960 306388
rect 220688 306348 220694 306360
rect 247954 306348 247960 306360
rect 248012 306348 248018 306400
rect 111794 306280 111800 306332
rect 111852 306320 111858 306332
rect 136174 306320 136180 306332
rect 111852 306292 136180 306320
rect 111852 306280 111858 306292
rect 136174 306280 136180 306292
rect 136232 306280 136238 306332
rect 111886 306212 111892 306264
rect 111944 306252 111950 306264
rect 122098 306252 122104 306264
rect 111944 306224 122104 306252
rect 111944 306212 111950 306224
rect 122098 306212 122104 306224
rect 122156 306212 122162 306264
rect 136082 305600 136088 305652
rect 136140 305640 136146 305652
rect 155494 305640 155500 305652
rect 136140 305612 155500 305640
rect 136140 305600 136146 305612
rect 155494 305600 155500 305612
rect 155552 305600 155558 305652
rect 244918 305600 244924 305652
rect 244976 305640 244982 305652
rect 257614 305640 257620 305652
rect 244976 305612 257620 305640
rect 244976 305600 244982 305612
rect 257614 305600 257620 305612
rect 257672 305600 257678 305652
rect 154574 305532 154580 305584
rect 154632 305572 154638 305584
rect 155678 305572 155684 305584
rect 154632 305544 155684 305572
rect 154632 305532 154638 305544
rect 155678 305532 155684 305544
rect 155736 305532 155742 305584
rect 154942 305464 154948 305516
rect 155000 305504 155006 305516
rect 155310 305504 155316 305516
rect 155000 305476 155316 305504
rect 155000 305464 155006 305476
rect 155310 305464 155316 305476
rect 155368 305464 155374 305516
rect 220722 305328 220728 305380
rect 220780 305368 220786 305380
rect 224310 305368 224316 305380
rect 220780 305340 224316 305368
rect 220780 305328 220786 305340
rect 224310 305328 224316 305340
rect 224368 305328 224374 305380
rect 155126 305192 155132 305244
rect 155184 305232 155190 305244
rect 155402 305232 155408 305244
rect 155184 305204 155408 305232
rect 155184 305192 155190 305204
rect 155402 305192 155408 305204
rect 155460 305192 155466 305244
rect 127618 305124 127624 305176
rect 127676 305164 127682 305176
rect 154850 305164 154856 305176
rect 127676 305136 154856 305164
rect 127676 305124 127682 305136
rect 154850 305124 154856 305136
rect 154908 305124 154914 305176
rect 220722 305124 220728 305176
rect 220780 305164 220786 305176
rect 243814 305164 243820 305176
rect 220780 305136 243820 305164
rect 220780 305124 220786 305136
rect 243814 305124 243820 305136
rect 243872 305124 243878 305176
rect 124858 305056 124864 305108
rect 124916 305096 124922 305108
rect 154758 305096 154764 305108
rect 124916 305068 154764 305096
rect 124916 305056 124922 305068
rect 154758 305056 154764 305068
rect 154816 305056 154822 305108
rect 220630 305056 220636 305108
rect 220688 305096 220694 305108
rect 245010 305096 245016 305108
rect 220688 305068 245016 305096
rect 220688 305056 220694 305068
rect 245010 305056 245016 305068
rect 245068 305056 245074 305108
rect 3234 304988 3240 305040
rect 3292 305028 3298 305040
rect 30098 305028 30104 305040
rect 3292 305000 30104 305028
rect 3292 304988 3298 305000
rect 30098 304988 30104 305000
rect 30156 304988 30162 305040
rect 114094 304988 114100 305040
rect 114152 305028 114158 305040
rect 154942 305028 154948 305040
rect 114152 305000 154948 305028
rect 114152 304988 114158 305000
rect 154942 304988 154948 305000
rect 155000 304988 155006 305040
rect 220538 304988 220544 305040
rect 220596 305028 220602 305040
rect 246666 305028 246672 305040
rect 220596 305000 246672 305028
rect 220596 304988 220602 305000
rect 246666 304988 246672 305000
rect 246724 304988 246730 305040
rect 111886 304920 111892 304972
rect 111944 304960 111950 304972
rect 141510 304960 141516 304972
rect 111944 304932 141516 304960
rect 111944 304920 111950 304932
rect 141510 304920 141516 304932
rect 141568 304920 141574 304972
rect 111794 304852 111800 304904
rect 111852 304892 111858 304904
rect 113818 304892 113824 304904
rect 111852 304864 113824 304892
rect 111852 304852 111858 304864
rect 113818 304852 113824 304864
rect 113876 304852 113882 304904
rect 112070 304444 112076 304496
rect 112128 304484 112134 304496
rect 112530 304484 112536 304496
rect 112128 304456 112536 304484
rect 112128 304444 112134 304456
rect 112530 304444 112536 304456
rect 112588 304444 112594 304496
rect 119522 304240 119528 304292
rect 119580 304280 119586 304292
rect 155126 304280 155132 304292
rect 119580 304252 155132 304280
rect 119580 304240 119586 304252
rect 155126 304240 155132 304252
rect 155184 304240 155190 304292
rect 115290 303832 115296 303884
rect 115348 303872 115354 303884
rect 154942 303872 154948 303884
rect 115348 303844 154948 303872
rect 115348 303832 115354 303844
rect 154942 303832 154948 303844
rect 155000 303832 155006 303884
rect 140314 303764 140320 303816
rect 140372 303804 140378 303816
rect 154574 303804 154580 303816
rect 140372 303776 154580 303804
rect 140372 303764 140378 303776
rect 154574 303764 154580 303776
rect 154632 303764 154638 303816
rect 220630 303764 220636 303816
rect 220688 303804 220694 303816
rect 231394 303804 231400 303816
rect 220688 303776 231400 303804
rect 220688 303764 220694 303776
rect 231394 303764 231400 303776
rect 231452 303764 231458 303816
rect 116762 303696 116768 303748
rect 116820 303736 116826 303748
rect 154850 303736 154856 303748
rect 116820 303708 154856 303736
rect 116820 303696 116826 303708
rect 154850 303696 154856 303708
rect 154908 303696 154914 303748
rect 220722 303696 220728 303748
rect 220780 303736 220786 303748
rect 239490 303736 239496 303748
rect 220780 303708 239496 303736
rect 220780 303696 220786 303708
rect 239490 303696 239496 303708
rect 239548 303696 239554 303748
rect 152642 303628 152648 303680
rect 152700 303668 152706 303680
rect 155494 303668 155500 303680
rect 152700 303640 155500 303668
rect 152700 303628 152706 303640
rect 155494 303628 155500 303640
rect 155552 303628 155558 303680
rect 220446 303628 220452 303680
rect 220504 303668 220510 303680
rect 250622 303668 250628 303680
rect 220504 303640 250628 303668
rect 220504 303628 220510 303640
rect 250622 303628 250628 303640
rect 250680 303628 250686 303680
rect 111886 303560 111892 303612
rect 111944 303600 111950 303612
rect 155310 303600 155316 303612
rect 111944 303572 155316 303600
rect 111944 303560 111950 303572
rect 155310 303560 155316 303572
rect 155368 303560 155374 303612
rect 223942 303560 223948 303612
rect 224000 303600 224006 303612
rect 256694 303600 256700 303612
rect 224000 303572 256700 303600
rect 224000 303560 224006 303572
rect 256694 303560 256700 303572
rect 256752 303560 256758 303612
rect 111794 303492 111800 303544
rect 111852 303532 111858 303544
rect 117222 303532 117228 303544
rect 111852 303504 117228 303532
rect 111852 303492 111858 303504
rect 117222 303492 117228 303504
rect 117280 303492 117286 303544
rect 141602 302880 141608 302932
rect 141660 302920 141666 302932
rect 154758 302920 154764 302932
rect 141660 302892 154764 302920
rect 141660 302880 141666 302892
rect 154758 302880 154764 302892
rect 154816 302880 154822 302932
rect 114002 302472 114008 302524
rect 114060 302512 114066 302524
rect 154942 302512 154948 302524
rect 114060 302484 154948 302512
rect 114060 302472 114066 302484
rect 154942 302472 154948 302484
rect 155000 302472 155006 302524
rect 138750 302404 138756 302456
rect 138808 302444 138814 302456
rect 154666 302444 154672 302456
rect 138808 302416 154672 302444
rect 138808 302404 138814 302416
rect 154666 302404 154672 302416
rect 154724 302404 154730 302456
rect 129182 302336 129188 302388
rect 129240 302376 129246 302388
rect 155126 302376 155132 302388
rect 129240 302348 155132 302376
rect 129240 302336 129246 302348
rect 155126 302336 155132 302348
rect 155184 302336 155190 302388
rect 219894 302336 219900 302388
rect 219952 302376 219958 302388
rect 224218 302376 224224 302388
rect 219952 302348 224224 302376
rect 219952 302336 219958 302348
rect 224218 302336 224224 302348
rect 224276 302336 224282 302388
rect 126238 302268 126244 302320
rect 126296 302308 126302 302320
rect 154850 302308 154856 302320
rect 126296 302280 154856 302308
rect 126296 302268 126302 302280
rect 154850 302268 154856 302280
rect 154908 302268 154914 302320
rect 220538 302268 220544 302320
rect 220596 302308 220602 302320
rect 241146 302308 241152 302320
rect 220596 302280 241152 302308
rect 220596 302268 220602 302280
rect 241146 302268 241152 302280
rect 241204 302268 241210 302320
rect 220722 302200 220728 302252
rect 220780 302240 220786 302252
rect 241054 302240 241060 302252
rect 220780 302212 241060 302240
rect 220780 302200 220786 302212
rect 241054 302200 241060 302212
rect 241112 302200 241118 302252
rect 111794 302132 111800 302184
rect 111852 302172 111858 302184
rect 140130 302172 140136 302184
rect 111852 302144 140136 302172
rect 111852 302132 111858 302144
rect 140130 302132 140136 302144
rect 140188 302132 140194 302184
rect 111886 302064 111892 302116
rect 111944 302104 111950 302116
rect 120718 302104 120724 302116
rect 111944 302076 120724 302104
rect 111944 302064 111950 302076
rect 120718 302064 120724 302076
rect 120776 302064 120782 302116
rect 154114 301384 154120 301436
rect 154172 301424 154178 301436
rect 154574 301424 154580 301436
rect 154172 301396 154580 301424
rect 154172 301384 154178 301396
rect 154574 301384 154580 301396
rect 154632 301384 154638 301436
rect 140222 301044 140228 301096
rect 140280 301084 140286 301096
rect 154574 301084 154580 301096
rect 140280 301056 154580 301084
rect 140280 301044 140286 301056
rect 154574 301044 154580 301056
rect 154632 301044 154638 301096
rect 219986 301044 219992 301096
rect 220044 301084 220050 301096
rect 232590 301084 232596 301096
rect 220044 301056 232596 301084
rect 220044 301044 220050 301056
rect 232590 301044 232596 301056
rect 232648 301044 232654 301096
rect 137370 300976 137376 301028
rect 137428 301016 137434 301028
rect 154850 301016 154856 301028
rect 137428 300988 154856 301016
rect 137428 300976 137434 300988
rect 154850 300976 154856 300988
rect 154908 300976 154914 301028
rect 220722 300976 220728 301028
rect 220780 301016 220786 301028
rect 233970 301016 233976 301028
rect 220780 300988 233976 301016
rect 220780 300976 220786 300988
rect 233970 300976 233976 300988
rect 234028 300976 234034 301028
rect 120810 300908 120816 300960
rect 120868 300948 120874 300960
rect 154758 300948 154764 300960
rect 120868 300920 154764 300948
rect 120868 300908 120874 300920
rect 154758 300908 154764 300920
rect 154816 300908 154822 300960
rect 220538 300908 220544 300960
rect 220596 300948 220602 300960
rect 234154 300948 234160 300960
rect 220596 300920 234160 300948
rect 220596 300908 220602 300920
rect 234154 300908 234160 300920
rect 234212 300908 234218 300960
rect 119430 300840 119436 300892
rect 119488 300880 119494 300892
rect 154666 300880 154672 300892
rect 119488 300852 154672 300880
rect 119488 300840 119494 300852
rect 154666 300840 154672 300852
rect 154724 300840 154730 300892
rect 220630 300840 220636 300892
rect 220688 300880 220694 300892
rect 256142 300880 256148 300892
rect 220688 300852 256148 300880
rect 220688 300840 220694 300852
rect 256142 300840 256148 300852
rect 256200 300840 256206 300892
rect 111978 300772 111984 300824
rect 112036 300812 112042 300824
rect 131758 300812 131764 300824
rect 112036 300784 131764 300812
rect 112036 300772 112042 300784
rect 131758 300772 131764 300784
rect 131816 300772 131822 300824
rect 246574 300772 246580 300824
rect 246632 300812 246638 300824
rect 256694 300812 256700 300824
rect 246632 300784 256700 300812
rect 246632 300772 246638 300784
rect 256694 300772 256700 300784
rect 256752 300772 256758 300824
rect 111886 300704 111892 300756
rect 111944 300744 111950 300756
rect 123478 300744 123484 300756
rect 111944 300716 123484 300744
rect 111944 300704 111950 300716
rect 123478 300704 123484 300716
rect 123536 300704 123542 300756
rect 111794 300636 111800 300688
rect 111852 300676 111858 300688
rect 119338 300676 119344 300688
rect 111852 300648 119344 300676
rect 111852 300636 111858 300648
rect 119338 300636 119344 300648
rect 119396 300636 119402 300688
rect 142982 299684 142988 299736
rect 143040 299724 143046 299736
rect 154666 299724 154672 299736
rect 143040 299696 154672 299724
rect 143040 299684 143046 299696
rect 154666 299684 154672 299696
rect 154724 299684 154730 299736
rect 141510 299616 141516 299668
rect 141568 299656 141574 299668
rect 154574 299656 154580 299668
rect 141568 299628 154580 299656
rect 141568 299616 141574 299628
rect 154574 299616 154580 299628
rect 154632 299616 154638 299668
rect 131850 299548 131856 299600
rect 131908 299588 131914 299600
rect 154758 299588 154764 299600
rect 131908 299560 154764 299588
rect 131908 299548 131914 299560
rect 154758 299548 154764 299560
rect 154816 299548 154822 299600
rect 220630 299548 220636 299600
rect 220688 299588 220694 299600
rect 236638 299588 236644 299600
rect 220688 299560 236644 299588
rect 220688 299548 220694 299560
rect 236638 299548 236644 299560
rect 236696 299548 236702 299600
rect 113910 299480 113916 299532
rect 113968 299520 113974 299532
rect 154850 299520 154856 299532
rect 113968 299492 154856 299520
rect 113968 299480 113974 299492
rect 154850 299480 154856 299492
rect 154908 299480 154914 299532
rect 220722 299480 220728 299532
rect 220780 299520 220786 299532
rect 251910 299520 251916 299532
rect 220780 299492 251916 299520
rect 220780 299480 220786 299492
rect 251910 299480 251916 299492
rect 251968 299480 251974 299532
rect 222930 299412 222936 299464
rect 222988 299452 222994 299464
rect 256694 299452 256700 299464
rect 222988 299424 256700 299452
rect 222988 299412 222994 299424
rect 256694 299412 256700 299424
rect 256752 299412 256758 299464
rect 111794 299140 111800 299192
rect 111852 299180 111858 299192
rect 115198 299180 115204 299192
rect 111852 299152 115204 299180
rect 111852 299140 111858 299152
rect 115198 299140 115204 299152
rect 115256 299140 115262 299192
rect 111794 298800 111800 298852
rect 111852 298840 111858 298852
rect 115842 298840 115848 298852
rect 111852 298812 115848 298840
rect 111852 298800 111858 298812
rect 115842 298800 115848 298812
rect 115900 298800 115906 298852
rect 123662 298732 123668 298784
rect 123720 298772 123726 298784
rect 155494 298772 155500 298784
rect 123720 298744 155500 298772
rect 123720 298732 123726 298744
rect 155494 298732 155500 298744
rect 155552 298732 155558 298784
rect 148410 298324 148416 298376
rect 148468 298364 148474 298376
rect 154942 298364 154948 298376
rect 148468 298336 154948 298364
rect 148468 298324 148474 298336
rect 154942 298324 154948 298336
rect 155000 298324 155006 298376
rect 149698 298256 149704 298308
rect 149756 298296 149762 298308
rect 154850 298296 154856 298308
rect 149756 298268 154856 298296
rect 149756 298256 149762 298268
rect 154850 298256 154856 298268
rect 154908 298256 154914 298308
rect 219986 298256 219992 298308
rect 220044 298296 220050 298308
rect 223114 298296 223120 298308
rect 220044 298268 223120 298296
rect 220044 298256 220050 298268
rect 223114 298256 223120 298268
rect 223172 298256 223178 298308
rect 144270 298188 144276 298240
rect 144328 298228 144334 298240
rect 154574 298228 154580 298240
rect 144328 298200 154580 298228
rect 144328 298188 144334 298200
rect 154574 298188 154580 298200
rect 154632 298188 154638 298240
rect 220538 298188 220544 298240
rect 220596 298228 220602 298240
rect 231302 298228 231308 298240
rect 220596 298200 231308 298228
rect 220596 298188 220602 298200
rect 231302 298188 231308 298200
rect 231360 298188 231366 298240
rect 123478 298120 123484 298172
rect 123536 298160 123542 298172
rect 154758 298160 154764 298172
rect 123536 298132 154764 298160
rect 123536 298120 123542 298132
rect 154758 298120 154764 298132
rect 154816 298120 154822 298172
rect 220722 298120 220728 298172
rect 220780 298160 220786 298172
rect 254762 298160 254768 298172
rect 220780 298132 254768 298160
rect 220780 298120 220786 298132
rect 254762 298120 254768 298132
rect 254820 298120 254826 298172
rect 111886 298052 111892 298104
rect 111944 298092 111950 298104
rect 144546 298092 144552 298104
rect 111944 298064 144552 298092
rect 111944 298052 111950 298064
rect 144546 298052 144552 298064
rect 144604 298052 144610 298104
rect 111794 297916 111800 297968
rect 111852 297956 111858 297968
rect 115106 297956 115112 297968
rect 111852 297928 115112 297956
rect 111852 297916 111858 297928
rect 115106 297916 115112 297928
rect 115164 297916 115170 297968
rect 220722 297576 220728 297628
rect 220780 297616 220786 297628
rect 223022 297616 223028 297628
rect 220780 297588 223028 297616
rect 220780 297576 220786 297588
rect 223022 297576 223028 297588
rect 223080 297576 223086 297628
rect 147030 297372 147036 297424
rect 147088 297412 147094 297424
rect 154666 297412 154672 297424
rect 147088 297384 154672 297412
rect 147088 297372 147094 297384
rect 154666 297372 154672 297384
rect 154724 297372 154730 297424
rect 151630 297168 151636 297220
rect 151688 297208 151694 297220
rect 155402 297208 155408 297220
rect 151688 297180 155408 297208
rect 151688 297168 151694 297180
rect 155402 297168 155408 297180
rect 155460 297168 155466 297220
rect 138842 296828 138848 296880
rect 138900 296868 138906 296880
rect 154574 296868 154580 296880
rect 138900 296840 154580 296868
rect 138900 296828 138906 296840
rect 154574 296828 154580 296840
rect 154632 296828 154638 296880
rect 116670 296760 116676 296812
rect 116728 296800 116734 296812
rect 154758 296800 154764 296812
rect 116728 296772 154764 296800
rect 116728 296760 116734 296772
rect 154758 296760 154764 296772
rect 154816 296760 154822 296812
rect 220722 296760 220728 296812
rect 220780 296800 220786 296812
rect 246574 296800 246580 296812
rect 220780 296772 246580 296800
rect 220780 296760 220786 296772
rect 246574 296760 246580 296772
rect 246632 296760 246638 296812
rect 115198 296692 115204 296744
rect 115256 296732 115262 296744
rect 154942 296732 154948 296744
rect 115256 296704 154948 296732
rect 115256 296692 115262 296704
rect 154942 296692 154948 296704
rect 155000 296692 155006 296744
rect 220630 296692 220636 296744
rect 220688 296732 220694 296744
rect 247862 296732 247868 296744
rect 220688 296704 247868 296732
rect 220688 296692 220694 296704
rect 247862 296692 247868 296704
rect 247920 296692 247926 296744
rect 111794 296624 111800 296676
rect 111852 296664 111858 296676
rect 155218 296664 155224 296676
rect 111852 296636 155224 296664
rect 111852 296624 111858 296636
rect 155218 296624 155224 296636
rect 155276 296624 155282 296676
rect 220262 296624 220268 296676
rect 220320 296664 220326 296676
rect 256694 296664 256700 296676
rect 220320 296636 256700 296664
rect 220320 296624 220326 296636
rect 256694 296624 256700 296636
rect 256752 296624 256758 296676
rect 111886 296556 111892 296608
rect 111944 296596 111950 296608
rect 139210 296596 139216 296608
rect 111944 296568 139216 296596
rect 111944 296556 111950 296568
rect 139210 296556 139216 296568
rect 139268 296556 139274 296608
rect 145558 295604 145564 295656
rect 145616 295644 145622 295656
rect 154574 295644 154580 295656
rect 145616 295616 154580 295644
rect 145616 295604 145622 295616
rect 154574 295604 154580 295616
rect 154632 295604 154638 295656
rect 131758 295536 131764 295588
rect 131816 295576 131822 295588
rect 154850 295576 154856 295588
rect 131816 295548 154856 295576
rect 131816 295536 131822 295548
rect 154850 295536 154856 295548
rect 154908 295536 154914 295588
rect 129090 295468 129096 295520
rect 129148 295508 129154 295520
rect 154758 295508 154764 295520
rect 129148 295480 154764 295508
rect 129148 295468 129154 295480
rect 154758 295468 154764 295480
rect 154816 295468 154822 295520
rect 219894 295468 219900 295520
rect 219952 295508 219958 295520
rect 228542 295508 228548 295520
rect 219952 295480 228548 295508
rect 219952 295468 219958 295480
rect 228542 295468 228548 295480
rect 228600 295468 228606 295520
rect 128998 295400 129004 295452
rect 129056 295440 129062 295452
rect 154666 295440 154672 295452
rect 129056 295412 154672 295440
rect 129056 295400 129062 295412
rect 154666 295400 154672 295412
rect 154724 295400 154730 295452
rect 220630 295400 220636 295452
rect 220688 295440 220694 295452
rect 231210 295440 231216 295452
rect 220688 295412 231216 295440
rect 220688 295400 220694 295412
rect 231210 295400 231216 295412
rect 231268 295400 231274 295452
rect 113818 295332 113824 295384
rect 113876 295372 113882 295384
rect 154942 295372 154948 295384
rect 113876 295344 154948 295372
rect 113876 295332 113882 295344
rect 154942 295332 154948 295344
rect 155000 295332 155006 295384
rect 220722 295332 220728 295384
rect 220780 295372 220786 295384
rect 256050 295372 256056 295384
rect 220780 295344 256056 295372
rect 220780 295332 220786 295344
rect 256050 295332 256056 295344
rect 256108 295332 256114 295384
rect 111886 295264 111892 295316
rect 111944 295304 111950 295316
rect 128170 295304 128176 295316
rect 111944 295276 128176 295304
rect 111944 295264 111950 295276
rect 128170 295264 128176 295276
rect 128228 295264 128234 295316
rect 222838 295264 222844 295316
rect 222896 295304 222902 295316
rect 256694 295304 256700 295316
rect 222896 295276 256700 295304
rect 222896 295264 222902 295276
rect 256694 295264 256700 295276
rect 256752 295264 256758 295316
rect 111794 295196 111800 295248
rect 111852 295236 111858 295248
rect 124030 295236 124036 295248
rect 111852 295208 124036 295236
rect 111852 295196 111858 295208
rect 124030 295196 124036 295208
rect 124088 295196 124094 295248
rect 151170 294244 151176 294296
rect 151228 294284 151234 294296
rect 154850 294284 154856 294296
rect 151228 294256 154856 294284
rect 151228 294244 151234 294256
rect 154850 294244 154856 294256
rect 154908 294244 154914 294296
rect 140130 294176 140136 294228
rect 140188 294216 140194 294228
rect 154666 294216 154672 294228
rect 140188 294188 154672 294216
rect 140188 294176 140194 294188
rect 154666 294176 154672 294188
rect 154724 294176 154730 294228
rect 220262 294176 220268 294228
rect 220320 294216 220326 294228
rect 225598 294216 225604 294228
rect 220320 294188 225604 294216
rect 220320 294176 220326 294188
rect 225598 294176 225604 294188
rect 225656 294176 225662 294228
rect 122098 294108 122104 294160
rect 122156 294148 122162 294160
rect 154574 294148 154580 294160
rect 122156 294120 154580 294148
rect 122156 294108 122162 294120
rect 154574 294108 154580 294120
rect 154632 294108 154638 294160
rect 220722 294108 220728 294160
rect 220780 294148 220786 294160
rect 254670 294148 254676 294160
rect 220780 294120 254676 294148
rect 220780 294108 220786 294120
rect 254670 294108 254676 294120
rect 254728 294108 254734 294160
rect 120902 294040 120908 294092
rect 120960 294080 120966 294092
rect 154758 294080 154764 294092
rect 120960 294052 154764 294080
rect 120960 294040 120966 294052
rect 154758 294040 154764 294052
rect 154816 294040 154822 294092
rect 112438 293972 112444 294024
rect 112496 294012 112502 294024
rect 154574 294012 154580 294024
rect 112496 293984 154580 294012
rect 112496 293972 112502 293984
rect 154574 293972 154580 293984
rect 154632 293972 154638 294024
rect 219894 293972 219900 294024
rect 219952 294012 219958 294024
rect 222930 294012 222936 294024
rect 219952 293984 222936 294012
rect 219952 293972 219958 293984
rect 222930 293972 222936 293984
rect 222988 293972 222994 294024
rect 111794 293904 111800 293956
rect 111852 293944 111858 293956
rect 121178 293944 121184 293956
rect 111852 293916 121184 293944
rect 111852 293904 111858 293916
rect 121178 293904 121184 293916
rect 121236 293904 121242 293956
rect 111886 293836 111892 293888
rect 111944 293876 111950 293888
rect 117130 293876 117136 293888
rect 111944 293848 117136 293876
rect 111944 293836 111950 293848
rect 117130 293836 117136 293848
rect 117188 293836 117194 293888
rect 250438 292748 250444 292800
rect 250496 292788 250502 292800
rect 257430 292788 257436 292800
rect 250496 292760 257436 292788
rect 250496 292748 250502 292760
rect 257430 292748 257436 292760
rect 257488 292748 257494 292800
rect 120718 292680 120724 292732
rect 120776 292720 120782 292732
rect 154574 292720 154580 292732
rect 120776 292692 154580 292720
rect 120776 292680 120782 292692
rect 154574 292680 154580 292692
rect 154632 292680 154638 292732
rect 220538 292680 220544 292732
rect 220596 292720 220602 292732
rect 228450 292720 228456 292732
rect 220596 292692 228456 292720
rect 220596 292680 220602 292692
rect 228450 292680 228456 292692
rect 228508 292680 228514 292732
rect 119338 292612 119344 292664
rect 119396 292652 119402 292664
rect 154666 292652 154672 292664
rect 119396 292624 154672 292652
rect 119396 292612 119402 292624
rect 154666 292612 154672 292624
rect 154724 292612 154730 292664
rect 154942 292612 154948 292664
rect 155000 292652 155006 292664
rect 155310 292652 155316 292664
rect 155000 292624 155316 292652
rect 155000 292612 155006 292624
rect 155310 292612 155316 292624
rect 155368 292612 155374 292664
rect 220722 292612 220728 292664
rect 220780 292652 220786 292664
rect 243722 292652 243728 292664
rect 220780 292624 243728 292652
rect 220780 292612 220786 292624
rect 243722 292612 243728 292624
rect 243780 292612 243786 292664
rect 116578 292544 116584 292596
rect 116636 292584 116642 292596
rect 154574 292584 154580 292596
rect 116636 292556 154580 292584
rect 116636 292544 116642 292556
rect 154574 292544 154580 292556
rect 154632 292544 154638 292596
rect 220630 292544 220636 292596
rect 220688 292584 220694 292596
rect 249334 292584 249340 292596
rect 220688 292556 249340 292584
rect 220688 292544 220694 292556
rect 249334 292544 249340 292556
rect 249392 292544 249398 292596
rect 111886 292476 111892 292528
rect 111944 292516 111950 292528
rect 137278 292516 137284 292528
rect 111944 292488 137284 292516
rect 111944 292476 111950 292488
rect 137278 292476 137284 292488
rect 137336 292476 137342 292528
rect 249610 292476 249616 292528
rect 249668 292516 249674 292528
rect 256694 292516 256700 292528
rect 249668 292488 256700 292516
rect 249668 292476 249674 292488
rect 256694 292476 256700 292488
rect 256752 292476 256758 292528
rect 111794 292408 111800 292460
rect 111852 292448 111858 292460
rect 119890 292448 119896 292460
rect 111852 292420 119896 292448
rect 111852 292408 111858 292420
rect 119890 292408 119896 292420
rect 119948 292408 119954 292460
rect 144546 291796 144552 291848
rect 144604 291836 144610 291848
rect 155126 291836 155132 291848
rect 144604 291808 155132 291836
rect 144604 291796 144610 291808
rect 155126 291796 155132 291808
rect 155184 291796 155190 291848
rect 219894 291320 219900 291372
rect 219952 291360 219958 291372
rect 227162 291360 227168 291372
rect 219952 291332 227168 291360
rect 219952 291320 219958 291332
rect 227162 291320 227168 291332
rect 227220 291320 227226 291372
rect 220630 291252 220636 291304
rect 220688 291292 220694 291304
rect 249150 291292 249156 291304
rect 220688 291264 249156 291292
rect 220688 291252 220694 291264
rect 249150 291252 249156 291264
rect 249208 291252 249214 291304
rect 220722 291184 220728 291236
rect 220780 291224 220786 291236
rect 250530 291224 250536 291236
rect 220780 291196 250536 291224
rect 220780 291184 220786 291196
rect 250530 291184 250536 291196
rect 250588 291184 250594 291236
rect 111886 291116 111892 291168
rect 111944 291156 111950 291168
rect 147490 291156 147496 291168
rect 111944 291128 147496 291156
rect 111944 291116 111950 291128
rect 147490 291116 147496 291128
rect 147548 291116 147554 291168
rect 248138 291116 248144 291168
rect 248196 291156 248202 291168
rect 256694 291156 256700 291168
rect 248196 291128 256700 291156
rect 248196 291116 248202 291128
rect 256694 291116 256700 291128
rect 256752 291116 256758 291168
rect 111794 291048 111800 291100
rect 111852 291088 111858 291100
rect 133230 291088 133236 291100
rect 111852 291060 133236 291088
rect 111852 291048 111858 291060
rect 133230 291048 133236 291060
rect 133288 291048 133294 291100
rect 137278 290436 137284 290488
rect 137336 290476 137342 290488
rect 154666 290476 154672 290488
rect 137336 290448 154672 290476
rect 137336 290436 137342 290448
rect 154666 290436 154672 290448
rect 154724 290436 154730 290488
rect 220722 289960 220728 290012
rect 220780 290000 220786 290012
rect 235350 290000 235356 290012
rect 220780 289972 235356 290000
rect 220780 289960 220786 289972
rect 235350 289960 235356 289972
rect 235408 289960 235414 290012
rect 220630 289892 220636 289944
rect 220688 289932 220694 289944
rect 244918 289932 244924 289944
rect 220688 289904 244924 289932
rect 220688 289892 220694 289904
rect 244918 289892 244924 289904
rect 244976 289892 244982 289944
rect 220722 289824 220728 289876
rect 220780 289864 220786 289876
rect 247770 289864 247776 289876
rect 220780 289836 247776 289864
rect 220780 289824 220786 289836
rect 247770 289824 247776 289836
rect 247828 289824 247834 289876
rect 111794 289756 111800 289808
rect 111852 289796 111858 289808
rect 141786 289796 141792 289808
rect 111852 289768 141792 289796
rect 111852 289756 111858 289768
rect 141786 289756 141792 289768
rect 141844 289756 141850 289808
rect 255958 289756 255964 289808
rect 256016 289796 256022 289808
rect 257798 289796 257804 289808
rect 256016 289768 257804 289796
rect 256016 289756 256022 289768
rect 257798 289756 257804 289768
rect 257856 289756 257862 289808
rect 111886 289688 111892 289740
rect 111944 289728 111950 289740
rect 134702 289728 134708 289740
rect 111944 289700 134708 289728
rect 111944 289688 111950 289700
rect 134702 289688 134708 289700
rect 134760 289688 134766 289740
rect 220538 288532 220544 288584
rect 220596 288572 220602 288584
rect 229830 288572 229836 288584
rect 220596 288544 229836 288572
rect 220596 288532 220602 288544
rect 229830 288532 229836 288544
rect 229888 288532 229894 288584
rect 220630 288464 220636 288516
rect 220688 288504 220694 288516
rect 236730 288504 236736 288516
rect 220688 288476 236736 288504
rect 220688 288464 220694 288476
rect 236730 288464 236736 288476
rect 236788 288464 236794 288516
rect 220722 288396 220728 288448
rect 220780 288436 220786 288448
rect 250438 288436 250444 288448
rect 220780 288408 250444 288436
rect 220780 288396 220786 288408
rect 250438 288396 250444 288408
rect 250496 288396 250502 288448
rect 111886 288328 111892 288380
rect 111944 288368 111950 288380
rect 144730 288368 144736 288380
rect 111944 288340 144736 288368
rect 111944 288328 111950 288340
rect 144730 288328 144736 288340
rect 144788 288328 144794 288380
rect 235626 288328 235632 288380
rect 235684 288368 235690 288380
rect 256694 288368 256700 288380
rect 235684 288340 256700 288368
rect 235684 288328 235690 288340
rect 256694 288328 256700 288340
rect 256752 288328 256758 288380
rect 111794 288260 111800 288312
rect 111852 288300 111858 288312
rect 126790 288300 126796 288312
rect 111852 288272 126796 288300
rect 111852 288260 111858 288272
rect 126790 288260 126796 288272
rect 126848 288260 126854 288312
rect 220722 287376 220728 287428
rect 220780 287416 220786 287428
rect 227070 287416 227076 287428
rect 220780 287388 227076 287416
rect 220780 287376 220786 287388
rect 227070 287376 227076 287388
rect 227128 287376 227134 287428
rect 220630 287104 220636 287156
rect 220688 287144 220694 287156
rect 235258 287144 235264 287156
rect 220688 287116 235264 287144
rect 220688 287104 220694 287116
rect 235258 287104 235264 287116
rect 235316 287104 235322 287156
rect 219526 287036 219532 287088
rect 219584 287076 219590 287088
rect 242158 287076 242164 287088
rect 219584 287048 242164 287076
rect 219584 287036 219590 287048
rect 242158 287036 242164 287048
rect 242216 287036 242222 287088
rect 111886 286968 111892 287020
rect 111944 287008 111950 287020
rect 148870 287008 148876 287020
rect 111944 286980 148876 287008
rect 111944 286968 111950 286980
rect 148870 286968 148876 286980
rect 148928 286968 148934 287020
rect 111794 286900 111800 286952
rect 111852 286940 111858 286952
rect 125134 286940 125140 286952
rect 111852 286912 125140 286940
rect 111852 286900 111858 286912
rect 125134 286900 125140 286912
rect 125192 286900 125198 286952
rect 219894 286696 219900 286748
rect 219952 286736 219958 286748
rect 222838 286736 222844 286748
rect 219952 286708 222844 286736
rect 219952 286696 219958 286708
rect 222838 286696 222844 286708
rect 222896 286696 222902 286748
rect 219894 286084 219900 286136
rect 219952 286124 219958 286136
rect 221734 286124 221740 286136
rect 219952 286096 221740 286124
rect 219952 286084 219958 286096
rect 221734 286084 221740 286096
rect 221792 286084 221798 286136
rect 220722 285880 220728 285932
rect 220780 285920 220786 285932
rect 255958 285920 255964 285932
rect 220780 285892 255964 285920
rect 220780 285880 220786 285892
rect 255958 285880 255964 285892
rect 256016 285880 256022 285932
rect 220630 285744 220636 285796
rect 220688 285784 220694 285796
rect 232774 285784 232780 285796
rect 220688 285756 232780 285784
rect 220688 285744 220694 285756
rect 232774 285744 232780 285756
rect 232832 285744 232838 285796
rect 111794 285608 111800 285660
rect 111852 285648 111858 285660
rect 140590 285648 140596 285660
rect 111852 285620 140596 285648
rect 111852 285608 111858 285620
rect 140590 285608 140596 285620
rect 140648 285608 140654 285660
rect 111886 285540 111892 285592
rect 111944 285580 111950 285592
rect 139118 285580 139124 285592
rect 111944 285552 139124 285580
rect 111944 285540 111950 285552
rect 139118 285540 139124 285552
rect 139176 285540 139182 285592
rect 111886 284248 111892 284300
rect 111944 284288 111950 284300
rect 151538 284288 151544 284300
rect 111944 284260 151544 284288
rect 111944 284248 111950 284260
rect 151538 284248 151544 284260
rect 151596 284248 151602 284300
rect 111794 284180 111800 284232
rect 111852 284220 111858 284232
rect 143350 284220 143356 284232
rect 111852 284192 143356 284220
rect 111852 284180 111858 284192
rect 143350 284180 143356 284192
rect 143408 284180 143414 284232
rect 224034 283568 224040 283620
rect 224092 283608 224098 283620
rect 257338 283608 257344 283620
rect 224092 283580 257344 283608
rect 224092 283568 224098 283580
rect 257338 283568 257344 283580
rect 257396 283568 257402 283620
rect 111794 282820 111800 282872
rect 111852 282860 111858 282872
rect 133598 282860 133604 282872
rect 111852 282832 133604 282860
rect 111852 282820 111858 282832
rect 133598 282820 133604 282832
rect 133656 282820 133662 282872
rect 227530 282820 227536 282872
rect 227588 282860 227594 282872
rect 256694 282860 256700 282872
rect 227588 282832 256700 282860
rect 227588 282820 227594 282832
rect 256694 282820 256700 282832
rect 256752 282820 256758 282872
rect 133230 282140 133236 282192
rect 133288 282180 133294 282192
rect 154942 282180 154948 282192
rect 133288 282152 154948 282180
rect 133288 282140 133294 282152
rect 154942 282140 154948 282152
rect 155000 282140 155006 282192
rect 111886 281460 111892 281512
rect 111944 281500 111950 281512
rect 128078 281500 128084 281512
rect 111944 281472 128084 281500
rect 111944 281460 111950 281472
rect 128078 281460 128084 281472
rect 128136 281460 128142 281512
rect 111794 281392 111800 281444
rect 111852 281432 111858 281444
rect 119798 281432 119804 281444
rect 111852 281404 119804 281432
rect 111852 281392 111858 281404
rect 119798 281392 119804 281404
rect 119856 281392 119862 281444
rect 111794 280100 111800 280152
rect 111852 280140 111858 280152
rect 145926 280140 145932 280152
rect 111852 280112 145932 280140
rect 111852 280100 111858 280112
rect 145926 280100 145932 280112
rect 145984 280100 145990 280152
rect 254946 280100 254952 280152
rect 255004 280140 255010 280152
rect 256694 280140 256700 280152
rect 255004 280112 256700 280140
rect 255004 280100 255010 280112
rect 256694 280100 256700 280112
rect 256752 280100 256758 280152
rect 111886 280032 111892 280084
rect 111944 280072 111950 280084
rect 133506 280072 133512 280084
rect 111944 280044 133512 280072
rect 111944 280032 111950 280044
rect 133506 280032 133512 280044
rect 133564 280032 133570 280084
rect 111886 278672 111892 278724
rect 111944 278712 111950 278724
rect 154114 278712 154120 278724
rect 111944 278684 154120 278712
rect 111944 278672 111950 278684
rect 154114 278672 154120 278684
rect 154172 278672 154178 278724
rect 224126 278672 224132 278724
rect 224184 278712 224190 278724
rect 256694 278712 256700 278724
rect 224184 278684 256700 278712
rect 224184 278672 224190 278684
rect 256694 278672 256700 278684
rect 256752 278672 256758 278724
rect 111794 278604 111800 278656
rect 111852 278644 111858 278656
rect 151446 278644 151452 278656
rect 111852 278616 151452 278644
rect 111852 278604 111858 278616
rect 151446 278604 151452 278616
rect 151504 278604 151510 278656
rect 111794 277312 111800 277364
rect 111852 277352 111858 277364
rect 155862 277352 155868 277364
rect 111852 277324 155868 277352
rect 111852 277312 111858 277324
rect 155862 277312 155868 277324
rect 155920 277312 155926 277364
rect 111886 277244 111892 277296
rect 111944 277284 111950 277296
rect 148778 277284 148784 277296
rect 111944 277256 148784 277284
rect 111944 277244 111950 277256
rect 148778 277244 148784 277256
rect 148836 277244 148842 277296
rect 111794 275952 111800 276004
rect 111852 275992 111858 276004
rect 153010 275992 153016 276004
rect 111852 275964 153016 275992
rect 111852 275952 111858 275964
rect 153010 275952 153016 275964
rect 153068 275952 153074 276004
rect 231670 275952 231676 276004
rect 231728 275992 231734 276004
rect 256694 275992 256700 276004
rect 231728 275964 256700 275992
rect 231728 275952 231734 275964
rect 256694 275952 256700 275964
rect 256752 275952 256758 276004
rect 111886 275884 111892 275936
rect 111944 275924 111950 275936
rect 132218 275924 132224 275936
rect 111944 275896 132224 275924
rect 111944 275884 111950 275896
rect 132218 275884 132224 275896
rect 132276 275884 132282 275936
rect 111886 274592 111892 274644
rect 111944 274632 111950 274644
rect 140498 274632 140504 274644
rect 111944 274604 140504 274632
rect 111944 274592 111950 274604
rect 140498 274592 140504 274604
rect 140556 274592 140562 274644
rect 228910 274592 228916 274644
rect 228968 274632 228974 274644
rect 256694 274632 256700 274644
rect 228968 274604 256700 274632
rect 228968 274592 228974 274604
rect 256694 274592 256700 274604
rect 256752 274592 256758 274644
rect 111794 274524 111800 274576
rect 111852 274564 111858 274576
rect 129366 274564 129372 274576
rect 111852 274536 129372 274564
rect 111852 274524 111858 274536
rect 129366 274524 129372 274536
rect 129424 274524 129430 274576
rect 111886 273164 111892 273216
rect 111944 273204 111950 273216
rect 154022 273204 154028 273216
rect 111944 273176 154028 273204
rect 111944 273164 111950 273176
rect 154022 273164 154028 273176
rect 154080 273164 154086 273216
rect 111794 273028 111800 273080
rect 111852 273068 111858 273080
rect 114462 273068 114468 273080
rect 111852 273040 114468 273068
rect 111852 273028 111858 273040
rect 114462 273028 114468 273040
rect 114520 273028 114526 273080
rect 551278 271872 551284 271924
rect 551336 271912 551342 271924
rect 580166 271912 580172 271924
rect 551336 271884 580172 271912
rect 551336 271872 551342 271884
rect 580166 271872 580172 271884
rect 580224 271872 580230 271924
rect 111886 271804 111892 271856
rect 111944 271844 111950 271856
rect 147398 271844 147404 271856
rect 111944 271816 147404 271844
rect 111944 271804 111950 271816
rect 147398 271804 147404 271816
rect 147456 271804 147462 271856
rect 111794 271736 111800 271788
rect 111852 271776 111858 271788
rect 145834 271776 145840 271788
rect 111852 271748 145840 271776
rect 111852 271736 111858 271748
rect 145834 271736 145840 271748
rect 145892 271736 145898 271788
rect 111794 270444 111800 270496
rect 111852 270484 111858 270496
rect 155770 270484 155776 270496
rect 111852 270456 155776 270484
rect 111852 270444 111858 270456
rect 155770 270444 155776 270456
rect 155828 270444 155834 270496
rect 241238 270444 241244 270496
rect 241296 270484 241302 270496
rect 256694 270484 256700 270496
rect 241296 270456 256700 270484
rect 241296 270444 241302 270456
rect 256694 270444 256700 270456
rect 256752 270444 256758 270496
rect 111886 270376 111892 270428
rect 111944 270416 111950 270428
rect 150066 270416 150072 270428
rect 111944 270388 150072 270416
rect 111944 270376 111950 270388
rect 150066 270376 150072 270388
rect 150124 270376 150130 270428
rect 111886 269016 111892 269068
rect 111944 269056 111950 269068
rect 132126 269056 132132 269068
rect 111944 269028 132132 269056
rect 111944 269016 111950 269028
rect 132126 269016 132132 269028
rect 132184 269016 132190 269068
rect 111794 268948 111800 269000
rect 111852 268988 111858 269000
rect 115750 268988 115756 269000
rect 111852 268960 115756 268988
rect 111852 268948 111858 268960
rect 115750 268948 115756 268960
rect 115808 268948 115814 269000
rect 111794 267656 111800 267708
rect 111852 267696 111858 267708
rect 129274 267696 129280 267708
rect 111852 267668 129280 267696
rect 111852 267656 111858 267668
rect 129274 267656 129280 267668
rect 129332 267656 129338 267708
rect 111886 267588 111892 267640
rect 111944 267628 111950 267640
rect 122558 267628 122564 267640
rect 111944 267600 122564 267628
rect 111944 267588 111950 267600
rect 122558 267588 122564 267600
rect 122616 267588 122622 267640
rect 232866 266976 232872 267028
rect 232924 267016 232930 267028
rect 257430 267016 257436 267028
rect 232924 266988 257436 267016
rect 232924 266976 232930 266988
rect 257430 266976 257436 266988
rect 257488 266976 257494 267028
rect 3050 266364 3056 266416
rect 3108 266404 3114 266416
rect 30190 266404 30196 266416
rect 3108 266376 30196 266404
rect 3108 266364 3114 266376
rect 30190 266364 30196 266376
rect 30248 266364 30254 266416
rect 160370 266364 160376 266416
rect 160428 266404 160434 266416
rect 161566 266404 161572 266416
rect 160428 266376 161572 266404
rect 160428 266364 160434 266376
rect 161566 266364 161572 266376
rect 161624 266364 161630 266416
rect 111886 266296 111892 266348
rect 111944 266336 111950 266348
rect 137646 266336 137652 266348
rect 111944 266308 137652 266336
rect 111944 266296 111950 266308
rect 137646 266296 137652 266308
rect 137704 266296 137710 266348
rect 224862 266296 224868 266348
rect 224920 266336 224926 266348
rect 256694 266336 256700 266348
rect 224920 266308 256700 266336
rect 224920 266296 224926 266308
rect 256694 266296 256700 266308
rect 256752 266296 256758 266348
rect 111794 266228 111800 266280
rect 111852 266268 111858 266280
rect 115658 266268 115664 266280
rect 111852 266240 115664 266268
rect 111852 266228 111858 266240
rect 115658 266228 115664 266240
rect 115716 266228 115722 266280
rect 111886 264868 111892 264920
rect 111944 264908 111950 264920
rect 152918 264908 152924 264920
rect 111944 264880 152924 264908
rect 111944 264868 111950 264880
rect 152918 264868 152924 264880
rect 152976 264868 152982 264920
rect 231578 264868 231584 264920
rect 231636 264908 231642 264920
rect 256694 264908 256700 264920
rect 231636 264880 256700 264908
rect 231636 264868 231642 264880
rect 256694 264868 256700 264880
rect 256752 264868 256758 264920
rect 111794 264800 111800 264852
rect 111852 264840 111858 264852
rect 144638 264840 144644 264852
rect 111852 264812 144644 264840
rect 111852 264800 111858 264812
rect 144638 264800 144644 264812
rect 144696 264800 144702 264852
rect 111886 263508 111892 263560
rect 111944 263548 111950 263560
rect 151630 263548 151636 263560
rect 111944 263520 151636 263548
rect 111944 263508 111950 263520
rect 151630 263508 151636 263520
rect 151688 263508 151694 263560
rect 111794 263440 111800 263492
rect 111852 263480 111858 263492
rect 140406 263480 140412 263492
rect 111852 263452 140412 263480
rect 111852 263440 111858 263452
rect 140406 263440 140412 263452
rect 140464 263440 140470 263492
rect 161474 262896 161480 262948
rect 161532 262936 161538 262948
rect 162394 262936 162400 262948
rect 161532 262908 162400 262936
rect 161532 262896 161538 262908
rect 162394 262896 162400 262908
rect 162452 262896 162458 262948
rect 168374 262896 168380 262948
rect 168432 262936 168438 262948
rect 169018 262936 169024 262948
rect 168432 262908 169024 262936
rect 168432 262896 168438 262908
rect 169018 262896 169024 262908
rect 169076 262896 169082 262948
rect 169754 262896 169760 262948
rect 169812 262936 169818 262948
rect 170674 262936 170680 262948
rect 169812 262908 170680 262936
rect 169812 262896 169818 262908
rect 170674 262896 170680 262908
rect 170732 262896 170738 262948
rect 173894 262896 173900 262948
rect 173952 262936 173958 262948
rect 174814 262936 174820 262948
rect 173952 262908 174820 262936
rect 173952 262896 173958 262908
rect 174814 262896 174820 262908
rect 174872 262896 174878 262948
rect 176654 262896 176660 262948
rect 176712 262936 176718 262948
rect 177298 262936 177304 262948
rect 176712 262908 177304 262936
rect 176712 262896 176718 262908
rect 177298 262896 177304 262908
rect 177356 262896 177362 262948
rect 178034 262896 178040 262948
rect 178092 262936 178098 262948
rect 178954 262936 178960 262948
rect 178092 262908 178960 262936
rect 178092 262896 178098 262908
rect 178954 262896 178960 262908
rect 179012 262896 179018 262948
rect 186314 262896 186320 262948
rect 186372 262936 186378 262948
rect 187234 262936 187240 262948
rect 186372 262908 187240 262936
rect 186372 262896 186378 262908
rect 187234 262896 187240 262908
rect 187292 262896 187298 262948
rect 190454 262896 190460 262948
rect 190512 262936 190518 262948
rect 191374 262936 191380 262948
rect 190512 262908 191380 262936
rect 190512 262896 190518 262908
rect 191374 262896 191380 262908
rect 191432 262896 191438 262948
rect 111794 262148 111800 262200
rect 111852 262188 111858 262200
rect 149974 262188 149980 262200
rect 111852 262160 149980 262188
rect 111852 262148 111858 262160
rect 149974 262148 149980 262160
rect 150032 262148 150038 262200
rect 228818 262148 228824 262200
rect 228876 262188 228882 262200
rect 256694 262188 256700 262200
rect 228876 262160 256700 262188
rect 228876 262148 228882 262160
rect 256694 262148 256700 262160
rect 256752 262148 256758 262200
rect 194594 261264 194600 261316
rect 194652 261304 194658 261316
rect 195514 261304 195520 261316
rect 194652 261276 195520 261304
rect 194652 261264 194658 261276
rect 195514 261264 195520 261276
rect 195572 261264 195578 261316
rect 202874 261264 202880 261316
rect 202932 261304 202938 261316
rect 203794 261304 203800 261316
rect 202932 261276 203800 261304
rect 202932 261264 202938 261276
rect 203794 261264 203800 261276
rect 203852 261264 203858 261316
rect 112898 261060 112904 261112
rect 112956 261060 112962 261112
rect 112916 260964 112944 261060
rect 113082 260992 113088 261044
rect 113140 260992 113146 261044
rect 112990 260964 112996 260976
rect 112916 260936 112996 260964
rect 112990 260924 112996 260936
rect 113048 260924 113054 260976
rect 112898 260856 112904 260908
rect 112956 260896 112962 260908
rect 113100 260896 113128 260992
rect 112956 260868 113128 260896
rect 112956 260856 112962 260868
rect 111794 260788 111800 260840
rect 111852 260828 111858 260840
rect 132034 260828 132040 260840
rect 111852 260800 132040 260828
rect 111852 260788 111858 260800
rect 132034 260788 132040 260800
rect 132092 260788 132098 260840
rect 226058 260788 226064 260840
rect 226116 260828 226122 260840
rect 256694 260828 256700 260840
rect 226116 260800 256700 260828
rect 226116 260788 226122 260800
rect 256694 260788 256700 260800
rect 256752 260788 256758 260840
rect 111886 260720 111892 260772
rect 111944 260760 111950 260772
rect 117038 260760 117044 260772
rect 111944 260732 117044 260760
rect 111944 260720 111950 260732
rect 117038 260720 117044 260732
rect 117096 260720 117102 260772
rect 112254 260652 112260 260704
rect 112312 260692 112318 260704
rect 113174 260692 113180 260704
rect 112312 260664 113180 260692
rect 112312 260652 112318 260664
rect 113174 260652 113180 260664
rect 113232 260652 113238 260704
rect 215294 260380 215300 260432
rect 215352 260420 215358 260432
rect 216214 260420 216220 260432
rect 215352 260392 216220 260420
rect 215352 260380 215358 260392
rect 216214 260380 216220 260392
rect 216272 260380 216278 260432
rect 111886 259360 111892 259412
rect 111944 259400 111950 259412
rect 118050 259400 118056 259412
rect 111944 259372 118056 259400
rect 111944 259360 111950 259372
rect 118050 259360 118056 259372
rect 118108 259360 118114 259412
rect 111794 259292 111800 259344
rect 111852 259332 111858 259344
rect 118142 259332 118148 259344
rect 111852 259304 118148 259332
rect 111852 259292 111858 259304
rect 118142 259292 118148 259304
rect 118200 259292 118206 259344
rect 551370 258068 551376 258120
rect 551428 258108 551434 258120
rect 580166 258108 580172 258120
rect 551428 258080 580172 258108
rect 551428 258068 551434 258080
rect 580166 258068 580172 258080
rect 580224 258068 580230 258120
rect 111886 258000 111892 258052
rect 111944 258040 111950 258052
rect 143258 258040 143264 258052
rect 111944 258012 143264 258040
rect 111944 258000 111950 258012
rect 143258 258000 143264 258012
rect 143316 258000 143322 258052
rect 238294 258000 238300 258052
rect 238352 258040 238358 258052
rect 256694 258040 256700 258052
rect 238352 258012 256700 258040
rect 238352 258000 238358 258012
rect 256694 258000 256700 258012
rect 256752 258000 256758 258052
rect 111794 257932 111800 257984
rect 111852 257972 111858 257984
rect 121086 257972 121092 257984
rect 111852 257944 121092 257972
rect 111852 257932 111858 257944
rect 121086 257932 121092 257944
rect 121144 257932 121150 257984
rect 111794 256640 111800 256692
rect 111852 256680 111858 256692
rect 137554 256680 137560 256692
rect 111852 256652 137560 256680
rect 111852 256640 111858 256652
rect 137554 256640 137560 256652
rect 137612 256640 137618 256692
rect 234338 256640 234344 256692
rect 234396 256680 234402 256692
rect 256694 256680 256700 256692
rect 234396 256652 256700 256680
rect 234396 256640 234402 256652
rect 256694 256640 256700 256652
rect 256752 256640 256758 256692
rect 111794 255212 111800 255264
rect 111852 255252 111858 255264
rect 151354 255252 151360 255264
rect 111852 255224 151360 255252
rect 111852 255212 111858 255224
rect 151354 255212 151360 255224
rect 151412 255212 151418 255264
rect 3510 253920 3516 253972
rect 3568 253960 3574 253972
rect 26878 253960 26884 253972
rect 3568 253932 26884 253960
rect 3568 253920 3574 253932
rect 26878 253920 26884 253932
rect 26936 253920 26942 253972
rect 111794 253852 111800 253904
rect 111852 253892 111858 253904
rect 131942 253892 131948 253904
rect 111852 253864 131948 253892
rect 111852 253852 111858 253864
rect 131942 253852 131948 253864
rect 132000 253852 132006 253904
rect 236914 253852 236920 253904
rect 236972 253892 236978 253904
rect 256694 253892 256700 253904
rect 236972 253864 256700 253892
rect 236972 253852 236978 253864
rect 256694 253852 256700 253864
rect 256752 253852 256758 253904
rect 111886 253784 111892 253836
rect 111944 253824 111950 253836
rect 123938 253824 123944 253836
rect 111944 253796 123944 253824
rect 111944 253784 111950 253796
rect 123938 253784 123944 253796
rect 123996 253784 124002 253836
rect 111794 253716 111800 253768
rect 111852 253756 111858 253768
rect 120994 253756 121000 253768
rect 111852 253728 121000 253756
rect 111852 253716 111858 253728
rect 120994 253716 121000 253728
rect 121052 253716 121058 253768
rect 112346 252968 112352 253020
rect 112404 253008 112410 253020
rect 112714 253008 112720 253020
rect 112404 252980 112720 253008
rect 112404 252968 112410 252980
rect 112714 252968 112720 252980
rect 112772 252968 112778 253020
rect 111794 252492 111800 252544
rect 111852 252532 111858 252544
rect 122466 252532 122472 252544
rect 111852 252504 122472 252532
rect 111852 252492 111858 252504
rect 122466 252492 122472 252504
rect 122524 252492 122530 252544
rect 224770 252492 224776 252544
rect 224828 252532 224834 252544
rect 256694 252532 256700 252544
rect 224828 252504 256700 252532
rect 224828 252492 224834 252504
rect 256694 252492 256700 252504
rect 256752 252492 256758 252544
rect 111794 251132 111800 251184
rect 111852 251172 111858 251184
rect 149882 251172 149888 251184
rect 111852 251144 149888 251172
rect 111852 251132 111858 251144
rect 149882 251132 149888 251144
rect 149940 251132 149946 251184
rect 111886 251064 111892 251116
rect 111944 251104 111950 251116
rect 137462 251104 137468 251116
rect 111944 251076 137468 251104
rect 111944 251064 111950 251076
rect 137462 251064 137468 251076
rect 137520 251064 137526 251116
rect 111794 249704 111800 249756
rect 111852 249744 111858 249756
rect 153930 249744 153936 249756
rect 111852 249716 153936 249744
rect 111852 249704 111858 249716
rect 153930 249704 153936 249716
rect 153988 249704 153994 249756
rect 228726 249704 228732 249756
rect 228784 249744 228790 249756
rect 256694 249744 256700 249756
rect 228784 249716 256700 249744
rect 228784 249704 228790 249716
rect 256694 249704 256700 249716
rect 256752 249704 256758 249756
rect 111886 248344 111892 248396
rect 111944 248384 111950 248396
rect 130838 248384 130844 248396
rect 111944 248356 130844 248384
rect 111944 248344 111950 248356
rect 130838 248344 130844 248356
rect 130896 248344 130902 248396
rect 225966 248344 225972 248396
rect 226024 248384 226030 248396
rect 256694 248384 256700 248396
rect 226024 248356 256700 248384
rect 226024 248344 226030 248356
rect 256694 248344 256700 248356
rect 256752 248344 256758 248396
rect 111794 248276 111800 248328
rect 111852 248316 111858 248328
rect 114370 248316 114376 248328
rect 111852 248288 114376 248316
rect 111852 248276 111858 248288
rect 114370 248276 114376 248288
rect 114428 248276 114434 248328
rect 111886 246984 111892 247036
rect 111944 247024 111950 247036
rect 126698 247024 126704 247036
rect 111944 246996 126704 247024
rect 111944 246984 111950 246996
rect 126698 246984 126704 246996
rect 126756 246984 126762 247036
rect 111794 246916 111800 246968
rect 111852 246956 111858 246968
rect 115566 246956 115572 246968
rect 111852 246928 115572 246956
rect 111852 246916 111858 246928
rect 115566 246916 115572 246928
rect 115624 246916 115630 246968
rect 112898 246304 112904 246356
rect 112956 246344 112962 246356
rect 152826 246344 152832 246356
rect 112956 246316 152832 246344
rect 112956 246304 112962 246316
rect 152826 246304 152832 246316
rect 152884 246304 152890 246356
rect 111794 245556 111800 245608
rect 111852 245596 111858 245608
rect 147306 245596 147312 245608
rect 111852 245568 147312 245596
rect 111852 245556 111858 245568
rect 147306 245556 147312 245568
rect 147364 245556 147370 245608
rect 224678 245556 224684 245608
rect 224736 245596 224742 245608
rect 256694 245596 256700 245608
rect 224736 245568 256700 245596
rect 224736 245556 224742 245568
rect 256694 245556 256700 245568
rect 256752 245556 256758 245608
rect 111886 245488 111892 245540
rect 111944 245528 111950 245540
rect 116946 245528 116952 245540
rect 111944 245500 116952 245528
rect 111944 245488 111950 245500
rect 116946 245488 116952 245500
rect 117004 245488 117010 245540
rect 111794 244196 111800 244248
rect 111852 244236 111858 244248
rect 122374 244236 122380 244248
rect 111852 244208 122380 244236
rect 111852 244196 111858 244208
rect 122374 244196 122380 244208
rect 122432 244196 122438 244248
rect 235534 244196 235540 244248
rect 235592 244236 235598 244248
rect 256694 244236 256700 244248
rect 235592 244208 256700 244236
rect 235592 244196 235598 244208
rect 256694 244196 256700 244208
rect 256752 244196 256758 244248
rect 111978 243516 111984 243568
rect 112036 243556 112042 243568
rect 144454 243556 144460 243568
rect 112036 243528 144460 243556
rect 112036 243516 112042 243528
rect 144454 243516 144460 243528
rect 144512 243516 144518 243568
rect 111794 242836 111800 242888
rect 111852 242876 111858 242888
rect 133414 242876 133420 242888
rect 111852 242848 133420 242876
rect 111852 242836 111858 242848
rect 133414 242836 133420 242848
rect 133472 242836 133478 242888
rect 111886 242156 111892 242208
rect 111944 242196 111950 242208
rect 143166 242196 143172 242208
rect 111944 242168 143172 242196
rect 111944 242156 111950 242168
rect 143166 242156 143172 242168
rect 143224 242156 143230 242208
rect 111794 241408 111800 241460
rect 111852 241448 111858 241460
rect 133322 241448 133328 241460
rect 111852 241420 133328 241448
rect 111852 241408 111858 241420
rect 133322 241408 133328 241420
rect 133380 241408 133386 241460
rect 224586 241408 224592 241460
rect 224644 241448 224650 241460
rect 256694 241448 256700 241460
rect 224644 241420 256700 241448
rect 224644 241408 224650 241420
rect 256694 241408 256700 241420
rect 256752 241408 256758 241460
rect 112346 240728 112352 240780
rect 112404 240768 112410 240780
rect 119706 240768 119712 240780
rect 112404 240740 119712 240768
rect 112404 240728 112410 240740
rect 119706 240728 119712 240740
rect 119764 240728 119770 240780
rect 111794 240048 111800 240100
rect 111852 240088 111858 240100
rect 148686 240088 148692 240100
rect 111852 240060 148692 240088
rect 111852 240048 111858 240060
rect 148686 240048 148692 240060
rect 148744 240048 148750 240100
rect 231486 240048 231492 240100
rect 231544 240088 231550 240100
rect 256694 240088 256700 240100
rect 231544 240060 256700 240088
rect 231544 240048 231550 240060
rect 256694 240048 256700 240060
rect 256752 240048 256758 240100
rect 111886 239980 111892 240032
rect 111944 240020 111950 240032
rect 130746 240020 130752 240032
rect 111944 239992 130752 240020
rect 111944 239980 111950 239992
rect 130746 239980 130752 239992
rect 130804 239980 130810 240032
rect 111794 238688 111800 238740
rect 111852 238728 111858 238740
rect 127986 238728 127992 238740
rect 111852 238700 127992 238728
rect 111852 238688 111858 238700
rect 127986 238688 127992 238700
rect 128044 238688 128050 238740
rect 111886 238484 111892 238536
rect 111944 238524 111950 238536
rect 114278 238524 114284 238536
rect 111944 238496 114284 238524
rect 111944 238484 111950 238496
rect 114278 238484 114284 238496
rect 114336 238484 114342 238536
rect 227438 238008 227444 238060
rect 227496 238048 227502 238060
rect 257798 238048 257804 238060
rect 227496 238020 257804 238048
rect 227496 238008 227502 238020
rect 257798 238008 257804 238020
rect 257856 238008 257862 238060
rect 111794 237328 111800 237380
rect 111852 237368 111858 237380
rect 136082 237368 136088 237380
rect 111852 237340 136088 237368
rect 111852 237328 111858 237340
rect 136082 237328 136088 237340
rect 136140 237328 136146 237380
rect 228634 237328 228640 237380
rect 228692 237368 228698 237380
rect 256694 237368 256700 237380
rect 228692 237340 256700 237368
rect 228692 237328 228698 237340
rect 256694 237328 256700 237340
rect 256752 237328 256758 237380
rect 111886 236648 111892 236700
rect 111944 236688 111950 236700
rect 139026 236688 139032 236700
rect 111944 236660 139032 236688
rect 111944 236648 111950 236660
rect 139026 236648 139032 236660
rect 139084 236648 139090 236700
rect 111794 235900 111800 235952
rect 111852 235940 111858 235952
rect 122282 235940 122288 235952
rect 111852 235912 122288 235940
rect 111852 235900 111858 235912
rect 122282 235900 122288 235912
rect 122340 235900 122346 235952
rect 111886 235220 111892 235272
rect 111944 235260 111950 235272
rect 145650 235260 145656 235272
rect 111944 235232 145656 235260
rect 111944 235220 111950 235232
rect 145650 235220 145656 235232
rect 145708 235220 145714 235272
rect 111794 234540 111800 234592
rect 111852 234580 111858 234592
rect 148594 234580 148600 234592
rect 111852 234552 148600 234580
rect 111852 234540 111858 234552
rect 148594 234540 148600 234552
rect 148652 234540 148658 234592
rect 112346 233928 112352 233980
rect 112404 233968 112410 233980
rect 112622 233968 112628 233980
rect 112404 233940 112628 233968
rect 112404 233928 112410 233940
rect 112622 233928 112628 233940
rect 112680 233928 112686 233980
rect 111794 233860 111800 233912
rect 111852 233900 111858 233912
rect 147214 233900 147220 233912
rect 111852 233872 147220 233900
rect 111852 233860 111858 233872
rect 147214 233860 147220 233872
rect 147272 233860 147278 233912
rect 232774 233860 232780 233912
rect 232832 233900 232838 233912
rect 257338 233900 257344 233912
rect 232832 233872 257344 233900
rect 232832 233860 232838 233872
rect 257338 233860 257344 233872
rect 257396 233860 257402 233912
rect 236822 233180 236828 233232
rect 236880 233220 236886 233232
rect 256694 233220 256700 233232
rect 236880 233192 256700 233220
rect 236880 233180 236886 233192
rect 256694 233180 256700 233192
rect 256752 233180 256758 233232
rect 111794 232908 111800 232960
rect 111852 232948 111858 232960
rect 115474 232948 115480 232960
rect 111852 232920 115480 232948
rect 111852 232908 111858 232920
rect 115474 232908 115480 232920
rect 115532 232908 115538 232960
rect 112806 232500 112812 232552
rect 112864 232540 112870 232552
rect 145742 232540 145748 232552
rect 112864 232512 145748 232540
rect 112864 232500 112870 232512
rect 145742 232500 145748 232512
rect 145800 232500 145806 232552
rect 551462 231820 551468 231872
rect 551520 231860 551526 231872
rect 579614 231860 579620 231872
rect 551520 231832 579620 231860
rect 551520 231820 551526 231832
rect 579614 231820 579620 231832
rect 579672 231820 579678 231872
rect 111794 231752 111800 231804
rect 111852 231792 111858 231804
rect 130654 231792 130660 231804
rect 111852 231764 130660 231792
rect 111852 231752 111858 231764
rect 130654 231752 130660 231764
rect 130712 231752 130718 231804
rect 112898 231072 112904 231124
rect 112956 231112 112962 231124
rect 119614 231112 119620 231124
rect 112956 231084 119620 231112
rect 112956 231072 112962 231084
rect 119614 231072 119620 231084
rect 119672 231072 119678 231124
rect 111794 230392 111800 230444
rect 111852 230432 111858 230444
rect 127894 230432 127900 230444
rect 111852 230404 127900 230432
rect 111852 230392 111858 230404
rect 127894 230392 127900 230404
rect 127952 230392 127958 230444
rect 111886 230324 111892 230376
rect 111944 230364 111950 230376
rect 126606 230364 126612 230376
rect 111944 230336 126612 230364
rect 111944 230324 111950 230336
rect 126606 230324 126612 230336
rect 126664 230324 126670 230376
rect 111794 229032 111800 229084
rect 111852 229072 111858 229084
rect 125042 229072 125048 229084
rect 111852 229044 125048 229072
rect 111852 229032 111858 229044
rect 125042 229032 125048 229044
rect 125100 229032 125106 229084
rect 111886 228964 111892 229016
rect 111944 229004 111950 229016
rect 123846 229004 123852 229016
rect 111944 228976 123852 229004
rect 111944 228964 111950 228976
rect 123846 228964 123852 228976
rect 123904 228964 123910 229016
rect 250714 228964 250720 229016
rect 250772 229004 250778 229016
rect 256694 229004 256700 229016
rect 250772 228976 256700 229004
rect 250772 228964 250778 228976
rect 256694 228964 256700 228976
rect 256752 228964 256758 229016
rect 111794 227672 111800 227724
rect 111852 227712 111858 227724
rect 122190 227712 122196 227724
rect 111852 227684 122196 227712
rect 111852 227672 111858 227684
rect 122190 227672 122196 227684
rect 122248 227672 122254 227724
rect 222746 227672 222752 227724
rect 222804 227712 222810 227724
rect 256694 227712 256700 227724
rect 222804 227684 256700 227712
rect 222804 227672 222810 227684
rect 256694 227672 256700 227684
rect 256752 227672 256758 227724
rect 111886 227604 111892 227656
rect 111944 227644 111950 227656
rect 116854 227644 116860 227656
rect 111944 227616 116860 227644
rect 111944 227604 111950 227616
rect 116854 227604 116860 227616
rect 116912 227604 116918 227656
rect 111794 225972 111800 226024
rect 111852 226012 111858 226024
rect 115382 226012 115388 226024
rect 111852 225984 115388 226012
rect 111852 225972 111858 225984
rect 115382 225972 115388 225984
rect 115440 225972 115446 226024
rect 111794 224884 111800 224936
rect 111852 224924 111858 224936
rect 144546 224924 144552 224936
rect 111852 224896 144552 224924
rect 111852 224884 111858 224896
rect 144546 224884 144552 224896
rect 144604 224884 144610 224936
rect 249518 224884 249524 224936
rect 249576 224924 249582 224936
rect 256694 224924 256700 224936
rect 249576 224896 256700 224924
rect 249576 224884 249582 224896
rect 256694 224884 256700 224896
rect 256752 224884 256758 224936
rect 111886 224816 111892 224868
rect 111944 224856 111950 224868
rect 134610 224856 134616 224868
rect 111944 224828 134616 224856
rect 111944 224816 111950 224828
rect 134610 224816 134616 224828
rect 134668 224816 134674 224868
rect 112806 224408 112812 224460
rect 112864 224448 112870 224460
rect 112990 224448 112996 224460
rect 112864 224420 112996 224448
rect 112864 224408 112870 224420
rect 112990 224408 112996 224420
rect 113048 224408 113054 224460
rect 111794 223524 111800 223576
rect 111852 223564 111858 223576
rect 147122 223564 147128 223576
rect 111852 223536 147128 223564
rect 111852 223524 111858 223536
rect 147122 223524 147128 223536
rect 147180 223524 147186 223576
rect 242342 223524 242348 223576
rect 242400 223564 242406 223576
rect 256694 223564 256700 223576
rect 242400 223536 256700 223564
rect 242400 223524 242406 223536
rect 256694 223524 256700 223536
rect 256752 223524 256758 223576
rect 111886 223456 111892 223508
rect 111944 223496 111950 223508
rect 130562 223496 130568 223508
rect 111944 223468 130568 223496
rect 111944 223456 111950 223468
rect 130562 223456 130568 223468
rect 130620 223456 130626 223508
rect 111794 222096 111800 222148
rect 111852 222136 111858 222148
rect 127802 222136 127808 222148
rect 111852 222108 127808 222136
rect 111852 222096 111858 222108
rect 127802 222096 127808 222108
rect 127860 222096 127866 222148
rect 111886 222028 111892 222080
rect 111944 222068 111950 222080
rect 126514 222068 126520 222080
rect 111944 222040 126520 222068
rect 111944 222028 111950 222040
rect 126514 222028 126520 222040
rect 126572 222028 126578 222080
rect 111794 220736 111800 220788
rect 111852 220776 111858 220788
rect 133138 220776 133144 220788
rect 111852 220748 133144 220776
rect 111852 220736 111858 220748
rect 133138 220736 133144 220748
rect 133196 220736 133202 220788
rect 223482 220736 223488 220788
rect 223540 220776 223546 220788
rect 256694 220776 256700 220788
rect 223540 220748 256700 220776
rect 223540 220736 223546 220748
rect 256694 220736 256700 220748
rect 256752 220736 256758 220788
rect 111886 220668 111892 220720
rect 111944 220708 111950 220720
rect 123754 220708 123760 220720
rect 111944 220680 123760 220708
rect 111944 220668 111950 220680
rect 123754 220668 123760 220680
rect 123812 220668 123818 220720
rect 112622 220056 112628 220108
rect 112680 220096 112686 220108
rect 152734 220096 152740 220108
rect 112680 220068 152740 220096
rect 112680 220056 112686 220068
rect 152734 220056 152740 220068
rect 152792 220056 152798 220108
rect 223390 219376 223396 219428
rect 223448 219416 223454 219428
rect 256694 219416 256700 219428
rect 223448 219388 256700 219416
rect 223448 219376 223454 219388
rect 256694 219376 256700 219388
rect 256752 219376 256758 219428
rect 111886 218696 111892 218748
rect 111944 218736 111950 218748
rect 151262 218736 151268 218748
rect 111944 218708 151268 218736
rect 111944 218696 111950 218708
rect 151262 218696 151268 218708
rect 151320 218696 151326 218748
rect 551554 218016 551560 218068
rect 551612 218056 551618 218068
rect 580166 218056 580172 218068
rect 551612 218028 580172 218056
rect 551612 218016 551618 218028
rect 580166 218016 580172 218028
rect 580224 218016 580230 218068
rect 111794 217948 111800 218000
rect 111852 217988 111858 218000
rect 114186 217988 114192 218000
rect 111852 217960 114192 217988
rect 111852 217948 111858 217960
rect 114186 217948 114192 217960
rect 114244 217948 114250 218000
rect 223298 217948 223304 218000
rect 223356 217988 223362 218000
rect 256694 217988 256700 218000
rect 223356 217960 256700 217988
rect 223356 217948 223362 217960
rect 256694 217948 256700 217960
rect 256752 217948 256758 218000
rect 112622 217268 112628 217320
rect 112680 217308 112686 217320
rect 149790 217308 149796 217320
rect 112680 217280 149796 217308
rect 112680 217268 112686 217280
rect 149790 217268 149796 217280
rect 149848 217268 149854 217320
rect 111794 216588 111800 216640
rect 111852 216628 111858 216640
rect 138934 216628 138940 216640
rect 111852 216600 138940 216628
rect 111852 216588 111858 216600
rect 138934 216588 138940 216600
rect 138992 216588 138998 216640
rect 112714 215908 112720 215960
rect 112772 215948 112778 215960
rect 129182 215948 129188 215960
rect 112772 215920 129188 215948
rect 112772 215908 112778 215920
rect 129182 215908 129188 215920
rect 129240 215908 129246 215960
rect 111794 215228 111800 215280
rect 111852 215268 111858 215280
rect 144362 215268 144368 215280
rect 111852 215240 144368 215268
rect 111852 215228 111858 215240
rect 144362 215228 144368 215240
rect 144420 215228 144426 215280
rect 252002 215228 252008 215280
rect 252060 215268 252066 215280
rect 256694 215268 256700 215280
rect 252060 215240 256700 215268
rect 252060 215228 252066 215240
rect 256694 215228 256700 215240
rect 256752 215228 256758 215280
rect 111886 215160 111892 215212
rect 111944 215200 111950 215212
rect 130470 215200 130476 215212
rect 111944 215172 130476 215200
rect 111944 215160 111950 215172
rect 130470 215160 130476 215172
rect 130528 215160 130534 215212
rect 3326 213936 3332 213988
rect 3384 213976 3390 213988
rect 30282 213976 30288 213988
rect 3384 213948 30288 213976
rect 3384 213936 3390 213948
rect 30282 213936 30288 213948
rect 30340 213936 30346 213988
rect 111794 213868 111800 213920
rect 111852 213908 111858 213920
rect 127710 213908 127716 213920
rect 111852 213880 127716 213908
rect 111852 213868 111858 213880
rect 127710 213868 127716 213880
rect 127768 213868 127774 213920
rect 221826 213868 221832 213920
rect 221884 213908 221890 213920
rect 256694 213908 256700 213920
rect 221884 213880 256700 213908
rect 221884 213868 221890 213880
rect 256694 213868 256700 213880
rect 256752 213868 256758 213920
rect 111886 213800 111892 213852
rect 111944 213840 111950 213852
rect 126422 213840 126428 213852
rect 111944 213812 126428 213840
rect 111944 213800 111950 213812
rect 126422 213800 126428 213812
rect 126480 213800 126486 213852
rect 111794 212440 111800 212492
rect 111852 212480 111858 212492
rect 124950 212480 124956 212492
rect 111852 212452 124956 212480
rect 111852 212440 111858 212452
rect 124950 212440 124956 212452
rect 125008 212440 125014 212492
rect 111886 212372 111892 212424
rect 111944 212412 111950 212424
rect 123570 212412 123576 212424
rect 111944 212384 123576 212412
rect 111944 212372 111950 212384
rect 123570 212372 123576 212384
rect 123628 212372 123634 212424
rect 111794 211080 111800 211132
rect 111852 211120 111858 211132
rect 141694 211120 141700 211132
rect 111852 211092 141700 211120
rect 111852 211080 111858 211092
rect 141694 211080 141700 211092
rect 141752 211080 141758 211132
rect 239674 211080 239680 211132
rect 239732 211120 239738 211132
rect 256694 211120 256700 211132
rect 239732 211092 256700 211120
rect 239732 211080 239738 211092
rect 256694 211080 256700 211092
rect 256752 211080 256758 211132
rect 111886 211012 111892 211064
rect 111944 211052 111950 211064
rect 117958 211052 117964 211064
rect 111944 211024 117964 211052
rect 111944 211012 111950 211024
rect 117958 211012 117964 211024
rect 118016 211012 118022 211064
rect 111794 209720 111800 209772
rect 111852 209760 111858 209772
rect 155678 209760 155684 209772
rect 111852 209732 155684 209760
rect 111852 209720 111858 209732
rect 155678 209720 155684 209732
rect 155736 209720 155742 209772
rect 111794 209040 111800 209092
rect 111852 209080 111858 209092
rect 148502 209080 148508 209092
rect 111852 209052 148508 209080
rect 111852 209040 111858 209052
rect 148502 209040 148508 209052
rect 148560 209040 148566 209092
rect 112622 207748 112628 207800
rect 112680 207788 112686 207800
rect 120902 207788 120908 207800
rect 112680 207760 120908 207788
rect 112680 207748 112686 207760
rect 120902 207748 120908 207760
rect 120960 207748 120966 207800
rect 111978 207680 111984 207732
rect 112036 207720 112042 207732
rect 127618 207720 127624 207732
rect 112036 207692 127624 207720
rect 112036 207680 112042 207692
rect 127618 207680 127624 207692
rect 127676 207680 127682 207732
rect 112070 207612 112076 207664
rect 112128 207652 112134 207664
rect 152642 207652 152648 207664
rect 112128 207624 152648 207652
rect 112128 207612 112134 207624
rect 152642 207612 152648 207624
rect 152700 207612 152706 207664
rect 111794 206932 111800 206984
rect 111852 206972 111858 206984
rect 143074 206972 143080 206984
rect 111852 206944 143080 206972
rect 111852 206932 111858 206944
rect 143074 206932 143080 206944
rect 143132 206932 143138 206984
rect 254854 206932 254860 206984
rect 254912 206972 254918 206984
rect 256694 206972 256700 206984
rect 254912 206944 256700 206972
rect 254912 206932 254918 206944
rect 256694 206932 256700 206944
rect 256752 206932 256758 206984
rect 111886 206864 111892 206916
rect 111944 206904 111950 206916
rect 130378 206904 130384 206916
rect 111944 206876 130384 206904
rect 111944 206864 111950 206876
rect 130378 206864 130384 206876
rect 130436 206864 130442 206916
rect 111794 205572 111800 205624
rect 111852 205612 111858 205624
rect 126330 205612 126336 205624
rect 111852 205584 126336 205612
rect 111852 205572 111858 205584
rect 126330 205572 126336 205584
rect 126388 205572 126394 205624
rect 225874 205572 225880 205624
rect 225932 205612 225938 205624
rect 256694 205612 256700 205624
rect 225932 205584 256700 205612
rect 225932 205572 225938 205584
rect 256694 205572 256700 205584
rect 256752 205572 256758 205624
rect 111886 205504 111892 205556
rect 111944 205544 111950 205556
rect 124858 205544 124864 205556
rect 111944 205516 124864 205544
rect 111944 205504 111950 205516
rect 124858 205504 124864 205516
rect 124916 205504 124922 205556
rect 111794 204212 111800 204264
rect 111852 204252 111858 204264
rect 123662 204252 123668 204264
rect 111852 204224 123668 204252
rect 111852 204212 111858 204224
rect 123662 204212 123668 204224
rect 123720 204212 123726 204264
rect 111886 204008 111892 204060
rect 111944 204048 111950 204060
rect 114094 204048 114100 204060
rect 111944 204020 114100 204048
rect 111944 204008 111950 204020
rect 114094 204008 114100 204020
rect 114152 204008 114158 204060
rect 111794 202784 111800 202836
rect 111852 202824 111858 202836
rect 119522 202824 119528 202836
rect 111852 202796 119528 202824
rect 111852 202784 111858 202796
rect 119522 202784 119528 202796
rect 119580 202784 119586 202836
rect 248046 202784 248052 202836
rect 248104 202824 248110 202836
rect 256694 202824 256700 202836
rect 248104 202796 256700 202824
rect 248104 202784 248110 202796
rect 256694 202784 256700 202796
rect 256752 202784 256758 202836
rect 111886 202716 111892 202768
rect 111944 202756 111950 202768
rect 116762 202756 116768 202768
rect 111944 202728 116768 202756
rect 111944 202716 111950 202728
rect 116762 202716 116768 202728
rect 116820 202716 116826 202768
rect 112254 202104 112260 202156
rect 112312 202144 112318 202156
rect 153838 202144 153844 202156
rect 112312 202116 153844 202144
rect 112312 202104 112318 202116
rect 153838 202104 153844 202116
rect 153896 202104 153902 202156
rect 3234 201492 3240 201544
rect 3292 201532 3298 201544
rect 29546 201532 29552 201544
rect 3292 201504 29552 201532
rect 3292 201492 3298 201504
rect 29546 201492 29552 201504
rect 29604 201492 29610 201544
rect 230198 201424 230204 201476
rect 230256 201464 230262 201476
rect 256694 201464 256700 201476
rect 230256 201436 256700 201464
rect 230256 201424 230262 201436
rect 256694 201424 256700 201436
rect 256752 201424 256758 201476
rect 111794 201356 111800 201408
rect 111852 201396 111858 201408
rect 115290 201396 115296 201408
rect 111852 201368 115296 201396
rect 111852 201356 111858 201368
rect 115290 201356 115296 201368
rect 115348 201356 115354 201408
rect 112990 200744 112996 200796
rect 113048 200784 113054 200796
rect 138842 200784 138848 200796
rect 113048 200756 138848 200784
rect 113048 200744 113054 200756
rect 138842 200744 138848 200756
rect 138900 200744 138906 200796
rect 111886 200064 111892 200116
rect 111944 200104 111950 200116
rect 141602 200104 141608 200116
rect 111944 200076 141608 200104
rect 111944 200064 111950 200076
rect 141602 200064 141608 200076
rect 141660 200064 141666 200116
rect 111794 199996 111800 200048
rect 111852 200036 111858 200048
rect 140314 200036 140320 200048
rect 111852 200008 140320 200036
rect 111852 199996 111858 200008
rect 140314 199996 140320 200008
rect 140372 199996 140378 200048
rect 111794 198636 111800 198688
rect 111852 198676 111858 198688
rect 114002 198676 114008 198688
rect 111852 198648 114008 198676
rect 111852 198636 111858 198648
rect 114002 198636 114008 198648
rect 114060 198636 114066 198688
rect 227346 198636 227352 198688
rect 227404 198676 227410 198688
rect 256694 198676 256700 198688
rect 227404 198648 256700 198676
rect 227404 198636 227410 198648
rect 256694 198636 256700 198648
rect 256752 198636 256758 198688
rect 111794 197276 111800 197328
rect 111852 197316 111858 197328
rect 126238 197316 126244 197328
rect 111852 197288 126244 197316
rect 111852 197276 111858 197288
rect 126238 197276 126244 197288
rect 126296 197276 126302 197328
rect 243906 197276 243912 197328
rect 243964 197316 243970 197328
rect 256694 197316 256700 197328
rect 243964 197288 256700 197316
rect 243964 197276 243970 197288
rect 256694 197276 256700 197288
rect 256752 197276 256758 197328
rect 111794 195916 111800 195968
rect 111852 195956 111858 195968
rect 138750 195956 138756 195968
rect 111852 195928 138756 195956
rect 111852 195916 111858 195928
rect 138750 195916 138756 195928
rect 138808 195916 138814 195968
rect 111886 195848 111892 195900
rect 111944 195888 111950 195900
rect 137370 195888 137376 195900
rect 111944 195860 137376 195888
rect 111944 195848 111950 195860
rect 137370 195848 137376 195860
rect 137428 195848 137434 195900
rect 112530 195236 112536 195288
rect 112588 195276 112594 195288
rect 112990 195276 112996 195288
rect 112588 195248 112996 195276
rect 112588 195236 112594 195248
rect 112990 195236 112996 195248
rect 113048 195236 113054 195288
rect 111794 194488 111800 194540
rect 111852 194528 111858 194540
rect 120810 194528 120816 194540
rect 111852 194500 120816 194528
rect 111852 194488 111858 194500
rect 120810 194488 120816 194500
rect 120868 194488 120874 194540
rect 223206 194488 223212 194540
rect 223264 194528 223270 194540
rect 256694 194528 256700 194540
rect 223264 194500 256700 194528
rect 223264 194488 223270 194500
rect 256694 194488 256700 194500
rect 256752 194488 256758 194540
rect 111886 194420 111892 194472
rect 111944 194460 111950 194472
rect 119430 194460 119436 194472
rect 111944 194432 119436 194460
rect 111944 194420 111950 194432
rect 119430 194420 119436 194432
rect 119488 194420 119494 194472
rect 112898 193808 112904 193860
rect 112956 193848 112962 193860
rect 149698 193848 149704 193860
rect 112956 193820 149704 193848
rect 112956 193808 112962 193820
rect 149698 193808 149704 193820
rect 149756 193808 149762 193860
rect 111886 193128 111892 193180
rect 111944 193168 111950 193180
rect 155586 193168 155592 193180
rect 111944 193140 155592 193168
rect 111944 193128 111950 193140
rect 155586 193128 155592 193140
rect 155644 193128 155650 193180
rect 249426 193128 249432 193180
rect 249484 193168 249490 193180
rect 256694 193168 256700 193180
rect 249484 193140 256700 193168
rect 249484 193128 249490 193140
rect 256694 193128 256700 193140
rect 256752 193128 256758 193180
rect 111794 193060 111800 193112
rect 111852 193100 111858 193112
rect 140222 193100 140228 193112
rect 111852 193072 140228 193100
rect 111852 193060 111858 193072
rect 140222 193060 140228 193072
rect 140280 193060 140286 193112
rect 111794 191700 111800 191752
rect 111852 191740 111858 191752
rect 133230 191740 133236 191752
rect 111852 191712 133236 191740
rect 111852 191700 111858 191712
rect 133230 191700 133236 191712
rect 133288 191700 133294 191752
rect 111794 191156 111800 191208
rect 111852 191196 111858 191208
rect 113910 191196 113916 191208
rect 111852 191168 113916 191196
rect 111852 191156 111858 191168
rect 113910 191156 113916 191168
rect 113968 191156 113974 191208
rect 111886 190408 111892 190460
rect 111944 190448 111950 190460
rect 142982 190448 142988 190460
rect 111944 190420 142988 190448
rect 111944 190408 111950 190420
rect 142982 190408 142988 190420
rect 143040 190408 143046 190460
rect 239582 190408 239588 190460
rect 239640 190448 239646 190460
rect 256694 190448 256700 190460
rect 239640 190420 256700 190448
rect 239640 190408 239646 190420
rect 256694 190408 256700 190420
rect 256752 190408 256758 190460
rect 111794 190340 111800 190392
rect 111852 190380 111858 190392
rect 131850 190380 131856 190392
rect 111852 190352 131856 190380
rect 111852 190340 111858 190352
rect 131850 190340 131856 190352
rect 131908 190340 131914 190392
rect 111886 188980 111892 189032
rect 111944 189020 111950 189032
rect 148410 189020 148416 189032
rect 111944 188992 148416 189020
rect 111944 188980 111950 188992
rect 148410 188980 148416 188992
rect 148468 188980 148474 189032
rect 230106 188980 230112 189032
rect 230164 189020 230170 189032
rect 256694 189020 256700 189032
rect 230164 188992 256700 189020
rect 230164 188980 230170 188992
rect 256694 188980 256700 188992
rect 256752 188980 256758 189032
rect 111794 188912 111800 188964
rect 111852 188952 111858 188964
rect 141510 188952 141516 188964
rect 111852 188924 141516 188952
rect 111852 188912 111858 188924
rect 141510 188912 141516 188924
rect 141568 188912 141574 188964
rect 111886 187620 111892 187672
rect 111944 187660 111950 187672
rect 144270 187660 144276 187672
rect 111944 187632 144276 187660
rect 111944 187620 111950 187632
rect 144270 187620 144276 187632
rect 144328 187620 144334 187672
rect 111794 187552 111800 187604
rect 111852 187592 111858 187604
rect 123478 187592 123484 187604
rect 111852 187564 123484 187592
rect 111852 187552 111858 187564
rect 123478 187552 123484 187564
rect 123536 187552 123542 187604
rect 111794 186260 111800 186312
rect 111852 186300 111858 186312
rect 147030 186300 147036 186312
rect 111852 186272 147036 186300
rect 111852 186260 111858 186272
rect 147030 186260 147036 186272
rect 147088 186260 147094 186312
rect 227254 186260 227260 186312
rect 227312 186300 227318 186312
rect 256694 186300 256700 186312
rect 227312 186272 256700 186300
rect 227312 186260 227318 186272
rect 256694 186260 256700 186272
rect 256752 186260 256758 186312
rect 111886 184832 111892 184884
rect 111944 184872 111950 184884
rect 116670 184872 116676 184884
rect 111944 184844 116676 184872
rect 111944 184832 111950 184844
rect 116670 184832 116676 184844
rect 116728 184832 116734 184884
rect 224494 184832 224500 184884
rect 224552 184872 224558 184884
rect 256694 184872 256700 184884
rect 224552 184844 256700 184872
rect 224552 184832 224558 184844
rect 256694 184832 256700 184844
rect 256752 184832 256758 184884
rect 111794 184764 111800 184816
rect 111852 184804 111858 184816
rect 115198 184804 115204 184816
rect 111852 184776 115204 184804
rect 111852 184764 111858 184776
rect 115198 184764 115204 184776
rect 115256 184764 115262 184816
rect 112806 184152 112812 184204
rect 112864 184192 112870 184204
rect 140130 184192 140136 184204
rect 112864 184164 140136 184192
rect 112864 184152 112870 184164
rect 140130 184152 140136 184164
rect 140188 184152 140194 184204
rect 111794 183472 111800 183524
rect 111852 183512 111858 183524
rect 137278 183512 137284 183524
rect 111852 183484 137284 183512
rect 111852 183472 111858 183484
rect 137278 183472 137284 183484
rect 137336 183472 137342 183524
rect 111794 182112 111800 182164
rect 111852 182152 111858 182164
rect 155494 182152 155500 182164
rect 111852 182124 155500 182152
rect 111852 182112 111858 182124
rect 155494 182112 155500 182124
rect 155552 182112 155558 182164
rect 235442 182112 235448 182164
rect 235500 182152 235506 182164
rect 256694 182152 256700 182164
rect 235500 182124 256700 182152
rect 235500 182112 235506 182124
rect 256694 182112 256700 182124
rect 256752 182112 256758 182164
rect 111794 181772 111800 181824
rect 111852 181812 111858 181824
rect 113818 181812 113824 181824
rect 111852 181784 113824 181812
rect 111852 181772 111858 181784
rect 113818 181772 113824 181784
rect 113876 181772 113882 181824
rect 111886 180752 111892 180804
rect 111944 180792 111950 180804
rect 128998 180792 129004 180804
rect 111944 180764 129004 180792
rect 111944 180752 111950 180764
rect 128998 180752 129004 180764
rect 129056 180752 129062 180804
rect 225782 180752 225788 180804
rect 225840 180792 225846 180804
rect 256694 180792 256700 180804
rect 225840 180764 256700 180792
rect 225840 180752 225846 180764
rect 256694 180752 256700 180764
rect 256752 180752 256758 180804
rect 111794 180684 111800 180736
rect 111852 180724 111858 180736
rect 129090 180724 129096 180736
rect 111852 180696 129096 180724
rect 111852 180684 111858 180696
rect 129090 180684 129096 180696
rect 129148 180684 129154 180736
rect 111886 179324 111892 179376
rect 111944 179364 111950 179376
rect 155402 179364 155408 179376
rect 111944 179336 155408 179364
rect 111944 179324 111950 179336
rect 155402 179324 155408 179336
rect 155460 179324 155466 179376
rect 111794 179256 111800 179308
rect 111852 179296 111858 179308
rect 145558 179296 145564 179308
rect 111852 179268 145564 179296
rect 111852 179256 111858 179268
rect 145558 179256 145564 179268
rect 145616 179256 145622 179308
rect 552658 178032 552664 178084
rect 552716 178072 552722 178084
rect 580166 178072 580172 178084
rect 552716 178044 580172 178072
rect 552716 178032 552722 178044
rect 580166 178032 580172 178044
rect 580224 178032 580230 178084
rect 245102 177964 245108 178016
rect 245160 178004 245166 178016
rect 256694 178004 256700 178016
rect 245160 177976 256700 178004
rect 245160 177964 245166 177976
rect 256694 177964 256700 177976
rect 256752 177964 256758 178016
rect 111978 177284 111984 177336
rect 112036 177324 112042 177336
rect 131758 177324 131764 177336
rect 112036 177296 131764 177324
rect 112036 177284 112042 177296
rect 131758 177284 131764 177296
rect 131816 177284 131822 177336
rect 111794 176604 111800 176656
rect 111852 176644 111858 176656
rect 151170 176644 151176 176656
rect 111852 176616 151176 176644
rect 111852 176604 111858 176616
rect 151170 176604 151176 176616
rect 151228 176604 151234 176656
rect 230014 176604 230020 176656
rect 230072 176644 230078 176656
rect 256694 176644 256700 176656
rect 230072 176616 256700 176644
rect 230072 176604 230078 176616
rect 256694 176604 256700 176616
rect 256752 176604 256758 176656
rect 111886 176536 111892 176588
rect 111944 176576 111950 176588
rect 122098 176576 122104 176588
rect 111944 176548 122104 176576
rect 111944 176536 111950 176548
rect 122098 176536 122104 176548
rect 122156 176536 122162 176588
rect 111794 173816 111800 173868
rect 111852 173856 111858 173868
rect 120718 173856 120724 173868
rect 111852 173828 120724 173856
rect 111852 173816 111858 173828
rect 120718 173816 120724 173828
rect 120776 173816 120782 173868
rect 111886 173748 111892 173800
rect 111944 173788 111950 173800
rect 119338 173788 119344 173800
rect 111944 173760 119344 173788
rect 111944 173748 111950 173760
rect 119338 173748 119344 173760
rect 119396 173748 119402 173800
rect 111794 172456 111800 172508
rect 111852 172496 111858 172508
rect 155218 172496 155224 172508
rect 111852 172468 155224 172496
rect 111852 172456 111858 172468
rect 155218 172456 155224 172468
rect 155276 172456 155282 172508
rect 246758 172456 246764 172508
rect 246816 172496 246822 172508
rect 256694 172496 256700 172508
rect 246816 172468 256700 172496
rect 246816 172456 246822 172468
rect 256694 172456 256700 172468
rect 256752 172456 256758 172508
rect 111886 171028 111892 171080
rect 111944 171068 111950 171080
rect 155310 171068 155316 171080
rect 111944 171040 155316 171068
rect 111944 171028 111950 171040
rect 155310 171028 155316 171040
rect 155368 171028 155374 171080
rect 234246 171028 234252 171080
rect 234304 171068 234310 171080
rect 256694 171068 256700 171080
rect 234304 171040 256700 171068
rect 234304 171028 234310 171040
rect 256694 171028 256700 171040
rect 256752 171028 256758 171080
rect 111794 170960 111800 171012
rect 111852 171000 111858 171012
rect 116578 171000 116584 171012
rect 111852 170972 116584 171000
rect 111852 170960 111858 170972
rect 116578 170960 116584 170972
rect 116636 170960 116642 171012
rect 224402 168308 224408 168360
rect 224460 168348 224466 168360
rect 256694 168348 256700 168360
rect 224460 168320 256700 168348
rect 224460 168308 224466 168320
rect 256694 168308 256700 168320
rect 256752 168308 256758 168360
rect 242250 166948 242256 167000
rect 242308 166988 242314 167000
rect 256694 166988 256700 167000
rect 242308 166960 256700 166988
rect 242308 166948 242314 166960
rect 256694 166948 256700 166960
rect 256752 166948 256758 167000
rect 225690 164160 225696 164212
rect 225748 164200 225754 164212
rect 256694 164200 256700 164212
rect 225748 164172 256700 164200
rect 225748 164160 225754 164172
rect 256694 164160 256700 164172
rect 256752 164160 256758 164212
rect 238202 162800 238208 162852
rect 238260 162840 238266 162852
rect 256694 162840 256700 162852
rect 238260 162812 256700 162840
rect 238260 162800 238266 162812
rect 256694 162800 256700 162812
rect 256752 162800 256758 162852
rect 3418 160760 3424 160812
rect 3476 160800 3482 160812
rect 134610 160800 134616 160812
rect 3476 160772 134616 160800
rect 3476 160760 3482 160772
rect 134610 160760 134616 160772
rect 134668 160760 134674 160812
rect 3326 160692 3332 160744
rect 3384 160732 3390 160744
rect 156874 160732 156880 160744
rect 3384 160704 156880 160732
rect 3384 160692 3390 160704
rect 156874 160692 156880 160704
rect 156932 160692 156938 160744
rect 232682 160012 232688 160064
rect 232740 160052 232746 160064
rect 256694 160052 256700 160064
rect 232740 160024 256700 160052
rect 232740 160012 232746 160024
rect 256694 160012 256700 160024
rect 256752 160012 256758 160064
rect 3602 159332 3608 159384
rect 3660 159372 3666 159384
rect 158346 159372 158352 159384
rect 3660 159344 158352 159372
rect 3660 159332 3666 159344
rect 158346 159332 158352 159344
rect 158404 159332 158410 159384
rect 3510 157972 3516 158024
rect 3568 158012 3574 158024
rect 155218 158012 155224 158024
rect 3568 157984 155224 158012
rect 3568 157972 3574 157984
rect 155218 157972 155224 157984
rect 155276 157972 155282 158024
rect 241146 157972 241152 158024
rect 241204 158012 241210 158024
rect 257522 158012 257528 158024
rect 241204 157984 257528 158012
rect 241204 157972 241210 157984
rect 257522 157972 257528 157984
rect 257580 157972 257586 158024
rect 247954 155864 247960 155916
rect 248012 155904 248018 155916
rect 256694 155904 256700 155916
rect 248012 155876 256700 155904
rect 248012 155864 248018 155876
rect 256694 155864 256700 155876
rect 256752 155864 256758 155916
rect 238110 154504 238116 154556
rect 238168 154544 238174 154556
rect 256694 154544 256700 154556
rect 238168 154516 256700 154544
rect 238168 154504 238174 154516
rect 256694 154504 256700 154516
rect 256752 154504 256758 154556
rect 550082 151784 550088 151836
rect 550140 151824 550146 151836
rect 579982 151824 579988 151836
rect 550140 151796 579988 151824
rect 550140 151784 550146 151796
rect 579982 151784 579988 151796
rect 580040 151784 580046 151836
rect 246666 151716 246672 151768
rect 246724 151756 246730 151768
rect 256694 151756 256700 151768
rect 246724 151728 256700 151756
rect 246724 151716 246730 151728
rect 256694 151716 256700 151728
rect 256752 151716 256758 151768
rect 245010 150356 245016 150408
rect 245068 150396 245074 150408
rect 256694 150396 256700 150408
rect 245068 150368 256700 150396
rect 245068 150356 245074 150368
rect 256694 150356 256700 150368
rect 256752 150356 256758 150408
rect 3418 149064 3424 149116
rect 3476 149104 3482 149116
rect 156966 149104 156972 149116
rect 3476 149076 156972 149104
rect 3476 149064 3482 149076
rect 156966 149064 156972 149076
rect 157024 149064 157030 149116
rect 224310 147568 224316 147620
rect 224368 147608 224374 147620
rect 256694 147608 256700 147620
rect 224368 147580 256700 147608
rect 224368 147568 224374 147580
rect 256694 147568 256700 147580
rect 256752 147568 256758 147620
rect 243814 146208 243820 146260
rect 243872 146248 243878 146260
rect 256694 146248 256700 146260
rect 243872 146220 256700 146248
rect 243872 146208 243878 146220
rect 256694 146208 256700 146220
rect 256752 146208 256758 146260
rect 250622 143488 250628 143540
rect 250680 143528 250686 143540
rect 256694 143528 256700 143540
rect 250680 143500 256700 143528
rect 250680 143488 250686 143500
rect 256694 143488 256700 143500
rect 256752 143488 256758 143540
rect 231394 142060 231400 142112
rect 231452 142100 231458 142112
rect 256694 142100 256700 142112
rect 231452 142072 256700 142100
rect 231452 142060 231458 142072
rect 256694 142060 256700 142072
rect 256752 142060 256758 142112
rect 194594 140700 194600 140752
rect 194652 140740 194658 140752
rect 195514 140740 195520 140752
rect 194652 140712 195520 140740
rect 194652 140700 194658 140712
rect 195514 140700 195520 140712
rect 195572 140700 195578 140752
rect 186314 140632 186320 140684
rect 186372 140672 186378 140684
rect 187234 140672 187240 140684
rect 186372 140644 187240 140672
rect 186372 140632 186378 140644
rect 187234 140632 187240 140644
rect 187292 140632 187298 140684
rect 178034 140428 178040 140480
rect 178092 140468 178098 140480
rect 178954 140468 178960 140480
rect 178092 140440 178960 140468
rect 178092 140428 178098 140440
rect 178954 140428 178960 140440
rect 179012 140428 179018 140480
rect 236730 140020 236736 140072
rect 236788 140060 236794 140072
rect 257430 140060 257436 140072
rect 236788 140032 257436 140060
rect 236788 140020 236794 140032
rect 257430 140020 257436 140032
rect 257488 140020 257494 140072
rect 215294 139884 215300 139936
rect 215352 139924 215358 139936
rect 216214 139924 216220 139936
rect 215352 139896 216220 139924
rect 215352 139884 215358 139896
rect 216214 139884 216220 139896
rect 216272 139884 216278 139936
rect 173894 139408 173900 139460
rect 173952 139448 173958 139460
rect 174814 139448 174820 139460
rect 173952 139420 174820 139448
rect 173952 139408 173958 139420
rect 174814 139408 174820 139420
rect 174872 139408 174878 139460
rect 239490 139340 239496 139392
rect 239548 139380 239554 139392
rect 256694 139380 256700 139392
rect 239548 139352 256700 139380
rect 239548 139340 239554 139352
rect 256694 139340 256700 139352
rect 256752 139340 256758 139392
rect 551646 137980 551652 138032
rect 551704 138020 551710 138032
rect 580166 138020 580172 138032
rect 551704 137992 580172 138020
rect 551704 137980 551710 137992
rect 580166 137980 580172 137992
rect 580224 137980 580230 138032
rect 168374 137300 168380 137352
rect 168432 137340 168438 137352
rect 169018 137340 169024 137352
rect 168432 137312 169024 137340
rect 168432 137300 168438 137312
rect 169018 137300 169024 137312
rect 169076 137300 169082 137352
rect 169754 137300 169760 137352
rect 169812 137340 169818 137352
rect 170674 137340 170680 137352
rect 169812 137312 170680 137340
rect 169812 137300 169818 137312
rect 170674 137300 170680 137312
rect 170732 137300 170738 137352
rect 176654 137300 176660 137352
rect 176712 137340 176718 137352
rect 177298 137340 177304 137352
rect 176712 137312 177304 137340
rect 176712 137300 176718 137312
rect 177298 137300 177304 137312
rect 177356 137300 177362 137352
rect 190454 137300 190460 137352
rect 190512 137340 190518 137352
rect 191374 137340 191380 137352
rect 190512 137312 191380 137340
rect 190512 137300 190518 137312
rect 191374 137300 191380 137312
rect 191432 137300 191438 137352
rect 202874 137300 202880 137352
rect 202932 137340 202938 137352
rect 203794 137340 203800 137352
rect 202932 137312 203800 137340
rect 202932 137300 202938 137312
rect 203794 137300 203800 137312
rect 203852 137300 203858 137352
rect 3418 136620 3424 136672
rect 3476 136660 3482 136672
rect 134702 136660 134708 136672
rect 3476 136632 134708 136660
rect 3476 136620 3482 136632
rect 134702 136620 134708 136632
rect 134760 136620 134766 136672
rect 224218 135192 224224 135244
rect 224276 135232 224282 135244
rect 256694 135232 256700 135244
rect 224276 135204 256700 135232
rect 224276 135192 224282 135204
rect 256694 135192 256700 135204
rect 256752 135192 256758 135244
rect 161382 133900 161388 133952
rect 161440 133940 161446 133952
rect 161658 133940 161664 133952
rect 161440 133912 161664 133940
rect 161440 133900 161446 133912
rect 161658 133900 161664 133912
rect 161716 133900 161722 133952
rect 30098 133832 30104 133884
rect 30156 133872 30162 133884
rect 151262 133872 151268 133884
rect 30156 133844 151268 133872
rect 30156 133832 30162 133844
rect 151262 133832 151268 133844
rect 151320 133832 151326 133884
rect 241054 133832 241060 133884
rect 241112 133872 241118 133884
rect 256694 133872 256700 133884
rect 241112 133844 256700 133872
rect 241112 133832 241118 133844
rect 256694 133832 256700 133844
rect 256752 133832 256758 133884
rect 29914 133764 29920 133816
rect 29972 133804 29978 133816
rect 151170 133804 151176 133816
rect 29972 133776 151176 133804
rect 29972 133764 29978 133776
rect 151170 133764 151176 133776
rect 151228 133764 151234 133816
rect 29546 133696 29552 133748
rect 29604 133736 29610 133748
rect 151354 133736 151360 133748
rect 29604 133708 151360 133736
rect 29604 133696 29610 133708
rect 151354 133696 151360 133708
rect 151412 133696 151418 133748
rect 30282 133628 30288 133680
rect 30340 133668 30346 133680
rect 154022 133668 154028 133680
rect 30340 133640 154028 133668
rect 30340 133628 30346 133640
rect 154022 133628 154028 133640
rect 154080 133628 154086 133680
rect 30190 133560 30196 133612
rect 30248 133600 30254 133612
rect 154114 133600 154120 133612
rect 30248 133572 154120 133600
rect 30248 133560 30254 133572
rect 154114 133560 154120 133572
rect 154172 133560 154178 133612
rect 29730 133492 29736 133544
rect 29788 133532 29794 133544
rect 153838 133532 153844 133544
rect 29788 133504 153844 133532
rect 29788 133492 29794 133504
rect 153838 133492 153844 133504
rect 153896 133492 153902 133544
rect 30006 133424 30012 133476
rect 30064 133464 30070 133476
rect 154206 133464 154212 133476
rect 30064 133436 154212 133464
rect 30064 133424 30070 133436
rect 154206 133424 154212 133436
rect 154264 133424 154270 133476
rect 26878 133356 26884 133408
rect 26936 133396 26942 133408
rect 151446 133396 151452 133408
rect 26936 133368 151452 133396
rect 26936 133356 26942 133368
rect 151446 133356 151452 133368
rect 151504 133356 151510 133408
rect 29822 133288 29828 133340
rect 29880 133328 29886 133340
rect 157150 133328 157156 133340
rect 29880 133300 157156 133328
rect 29880 133288 29886 133300
rect 157150 133288 157156 133300
rect 157208 133288 157214 133340
rect 29638 133220 29644 133272
rect 29696 133260 29702 133272
rect 157058 133260 157064 133272
rect 29696 133232 157064 133260
rect 29696 133220 29702 133232
rect 157058 133220 157064 133232
rect 157116 133220 157122 133272
rect 6914 133152 6920 133204
rect 6972 133192 6978 133204
rect 153930 133192 153936 133204
rect 6972 133164 153936 133192
rect 6972 133152 6978 133164
rect 153930 133152 153936 133164
rect 153988 133152 153994 133204
rect 136542 130364 136548 130416
rect 136600 130404 136606 130416
rect 154942 130404 154948 130416
rect 136600 130376 154948 130404
rect 136600 130364 136606 130376
rect 154942 130364 154948 130376
rect 155000 130364 155006 130416
rect 234154 129684 234160 129736
rect 234212 129724 234218 129736
rect 256694 129724 256700 129736
rect 234212 129696 256700 129724
rect 234212 129684 234218 129696
rect 256694 129684 256700 129696
rect 256752 129684 256758 129736
rect 136542 127576 136548 127628
rect 136600 127616 136606 127628
rect 154942 127616 154948 127628
rect 136600 127588 154948 127616
rect 136600 127576 136606 127588
rect 154942 127576 154948 127588
rect 155000 127576 155006 127628
rect 232590 126896 232596 126948
rect 232648 126936 232654 126948
rect 256694 126936 256700 126948
rect 232648 126908 256700 126936
rect 232648 126896 232654 126908
rect 256694 126896 256700 126908
rect 256752 126896 256758 126948
rect 154942 125644 154948 125656
rect 151786 125616 154948 125644
rect 136542 125536 136548 125588
rect 136600 125576 136606 125588
rect 151786 125576 151814 125616
rect 154942 125604 154948 125616
rect 155000 125604 155006 125656
rect 136600 125548 151814 125576
rect 136600 125536 136606 125548
rect 233970 125536 233976 125588
rect 234028 125576 234034 125588
rect 256694 125576 256700 125588
rect 234028 125548 256700 125576
rect 234028 125536 234034 125548
rect 256694 125536 256700 125548
rect 256752 125536 256758 125588
rect 136174 124108 136180 124160
rect 136232 124148 136238 124160
rect 154482 124148 154488 124160
rect 136232 124120 154488 124148
rect 136232 124108 136238 124120
rect 154482 124108 154488 124120
rect 154540 124108 154546 124160
rect 154942 121496 154948 121508
rect 151786 121468 154948 121496
rect 135254 121388 135260 121440
rect 135312 121428 135318 121440
rect 151786 121428 151814 121468
rect 154942 121456 154948 121468
rect 155000 121456 155006 121508
rect 135312 121400 151814 121428
rect 135312 121388 135318 121400
rect 236638 121388 236644 121440
rect 236696 121428 236702 121440
rect 256694 121428 256700 121440
rect 236696 121400 256700 121428
rect 236696 121388 236702 121400
rect 256694 121388 256700 121400
rect 256752 121388 256758 121440
rect 149054 120096 149060 120148
rect 149112 120136 149118 120148
rect 154574 120136 154580 120148
rect 149112 120108 154580 120136
rect 149112 120096 149118 120108
rect 154574 120096 154580 120108
rect 154632 120096 154638 120148
rect 251910 120028 251916 120080
rect 251968 120068 251974 120080
rect 256694 120068 256700 120080
rect 251968 120040 256700 120068
rect 251968 120028 251974 120040
rect 256694 120028 256700 120040
rect 256752 120028 256758 120080
rect 220446 119824 220452 119876
rect 220504 119864 220510 119876
rect 224218 119864 224224 119876
rect 220504 119836 224224 119864
rect 220504 119824 220510 119836
rect 224218 119824 224224 119836
rect 224276 119824 224282 119876
rect 135438 118600 135444 118652
rect 135496 118640 135502 118652
rect 149054 118640 149060 118652
rect 135496 118612 149060 118640
rect 135496 118600 135502 118612
rect 149054 118600 149060 118612
rect 149112 118600 149118 118652
rect 149054 117308 149060 117360
rect 149112 117348 149118 117360
rect 154574 117348 154580 117360
rect 149112 117320 154580 117348
rect 149112 117308 149118 117320
rect 154574 117308 154580 117320
rect 154632 117308 154638 117360
rect 231302 117240 231308 117292
rect 231360 117280 231366 117292
rect 256694 117280 256700 117292
rect 231360 117252 256700 117280
rect 231360 117240 231366 117252
rect 256694 117240 256700 117252
rect 256752 117240 256758 117292
rect 136542 115880 136548 115932
rect 136600 115920 136606 115932
rect 149054 115920 149060 115932
rect 136600 115892 149060 115920
rect 136600 115880 136606 115892
rect 149054 115880 149060 115892
rect 149112 115880 149118 115932
rect 223114 115880 223120 115932
rect 223172 115920 223178 115932
rect 256694 115920 256700 115932
rect 223172 115892 256700 115920
rect 223172 115880 223178 115892
rect 256694 115880 256700 115892
rect 256752 115880 256758 115932
rect 136542 113092 136548 113144
rect 136600 113132 136606 113144
rect 155402 113132 155408 113144
rect 136600 113104 155408 113132
rect 136600 113092 136606 113104
rect 155402 113092 155408 113104
rect 155460 113092 155466 113144
rect 254762 112888 254768 112940
rect 254820 112928 254826 112940
rect 256694 112928 256700 112940
rect 254820 112900 256700 112928
rect 254820 112888 254826 112900
rect 256694 112888 256700 112900
rect 256752 112888 256758 112940
rect 550174 111800 550180 111852
rect 550232 111840 550238 111852
rect 580166 111840 580172 111852
rect 550232 111812 580172 111840
rect 550232 111800 550238 111812
rect 580166 111800 580172 111812
rect 580224 111800 580230 111852
rect 247862 111732 247868 111784
rect 247920 111772 247926 111784
rect 256694 111772 256700 111784
rect 247920 111744 256700 111772
rect 247920 111732 247926 111744
rect 256694 111732 256700 111744
rect 256752 111732 256758 111784
rect 3418 110440 3424 110492
rect 3476 110480 3482 110492
rect 22738 110480 22744 110492
rect 3476 110452 22744 110480
rect 3476 110440 3482 110452
rect 22738 110440 22744 110452
rect 22796 110440 22802 110492
rect 136542 110372 136548 110424
rect 136600 110412 136606 110424
rect 154758 110412 154764 110424
rect 136600 110384 154764 110412
rect 136600 110372 136606 110384
rect 154758 110372 154764 110384
rect 154816 110372 154822 110424
rect 223022 108944 223028 108996
rect 223080 108984 223086 108996
rect 256694 108984 256700 108996
rect 223080 108956 256700 108984
rect 223080 108944 223086 108956
rect 256694 108944 256700 108956
rect 256752 108944 256758 108996
rect 136542 107584 136548 107636
rect 136600 107624 136606 107636
rect 154942 107624 154948 107636
rect 136600 107596 154948 107624
rect 136600 107584 136606 107596
rect 154942 107584 154948 107596
rect 155000 107584 155006 107636
rect 246574 107584 246580 107636
rect 246632 107624 246638 107636
rect 256694 107624 256700 107636
rect 246632 107596 256700 107624
rect 246632 107584 246638 107596
rect 256694 107584 256700 107596
rect 256752 107584 256758 107636
rect 136726 104864 136732 104916
rect 136784 104904 136790 104916
rect 154574 104904 154580 104916
rect 136784 104876 154580 104904
rect 136784 104864 136790 104876
rect 154574 104864 154580 104876
rect 154632 104864 154638 104916
rect 136542 104796 136548 104848
rect 136600 104836 136606 104848
rect 154850 104836 154856 104848
rect 136600 104808 154856 104836
rect 136600 104796 136606 104808
rect 154850 104796 154856 104808
rect 154908 104796 154914 104848
rect 220354 104796 220360 104848
rect 220412 104836 220418 104848
rect 256694 104836 256700 104848
rect 220412 104808 256700 104836
rect 220412 104796 220418 104808
rect 256694 104796 256700 104808
rect 256752 104796 256758 104848
rect 136174 103436 136180 103488
rect 136232 103476 136238 103488
rect 155494 103476 155500 103488
rect 136232 103448 155500 103476
rect 136232 103436 136238 103448
rect 155494 103436 155500 103448
rect 155552 103436 155558 103488
rect 231210 103436 231216 103488
rect 231268 103476 231274 103488
rect 256694 103476 256700 103488
rect 231268 103448 256700 103476
rect 231268 103436 231274 103448
rect 256694 103436 256700 103448
rect 256752 103436 256758 103488
rect 139394 102144 139400 102196
rect 139452 102184 139458 102196
rect 154574 102184 154580 102196
rect 139452 102156 154580 102184
rect 139452 102144 139458 102156
rect 154574 102144 154580 102156
rect 154632 102144 154638 102196
rect 138842 100716 138848 100768
rect 138900 100756 138906 100768
rect 154942 100756 154948 100768
rect 138900 100728 154948 100756
rect 138900 100716 138906 100728
rect 154942 100716 154948 100728
rect 155000 100716 155006 100768
rect 136174 100648 136180 100700
rect 136232 100688 136238 100700
rect 155310 100688 155316 100700
rect 136232 100660 155316 100688
rect 136232 100648 136238 100660
rect 155310 100648 155316 100660
rect 155368 100648 155374 100700
rect 228542 100648 228548 100700
rect 228600 100688 228606 100700
rect 256694 100688 256700 100700
rect 228600 100660 256700 100688
rect 228600 100648 228606 100660
rect 256694 100648 256700 100660
rect 256752 100648 256758 100700
rect 147030 99356 147036 99408
rect 147088 99396 147094 99408
rect 154942 99396 154948 99408
rect 147088 99368 154948 99396
rect 147088 99356 147094 99368
rect 154942 99356 154948 99368
rect 155000 99356 155006 99408
rect 3418 96636 3424 96688
rect 3476 96676 3482 96688
rect 24118 96676 24124 96688
rect 3476 96648 24124 96676
rect 3476 96636 3482 96648
rect 24118 96636 24124 96648
rect 24176 96636 24182 96688
rect 225598 96568 225604 96620
rect 225656 96608 225662 96620
rect 256694 96608 256700 96620
rect 225656 96580 256700 96608
rect 225656 96568 225662 96580
rect 256694 96568 256700 96580
rect 256752 96568 256758 96620
rect 136542 96228 136548 96280
rect 136600 96268 136606 96280
rect 139394 96268 139400 96280
rect 136600 96240 139400 96268
rect 136600 96228 136606 96240
rect 139394 96228 139400 96240
rect 139452 96228 139458 96280
rect 142154 95208 142160 95260
rect 142212 95248 142218 95260
rect 154942 95248 154948 95260
rect 142212 95220 154948 95248
rect 142212 95208 142218 95220
rect 154942 95208 154948 95220
rect 155000 95208 155006 95260
rect 222930 95140 222936 95192
rect 222988 95180 222994 95192
rect 256694 95180 256700 95192
rect 222988 95152 256700 95180
rect 222988 95140 222994 95152
rect 256694 95140 256700 95152
rect 256752 95140 256758 95192
rect 137278 94460 137284 94512
rect 137336 94500 137342 94512
rect 154850 94500 154856 94512
rect 137336 94472 154856 94500
rect 137336 94460 137342 94472
rect 154850 94460 154856 94472
rect 154908 94460 154914 94512
rect 140130 92488 140136 92540
rect 140188 92528 140194 92540
rect 154574 92528 154580 92540
rect 140188 92500 154580 92528
rect 140188 92488 140194 92500
rect 154574 92488 154580 92500
rect 154632 92488 154638 92540
rect 136082 92420 136088 92472
rect 136140 92460 136146 92472
rect 138842 92460 138848 92472
rect 136140 92432 138848 92460
rect 136140 92420 136146 92432
rect 138842 92420 138848 92432
rect 138900 92420 138906 92472
rect 254670 92420 254676 92472
rect 254728 92460 254734 92472
rect 256694 92460 256700 92472
rect 254728 92432 256700 92460
rect 254728 92420 254734 92432
rect 256694 92420 256700 92432
rect 256752 92420 256758 92472
rect 138750 91060 138756 91112
rect 138808 91100 138814 91112
rect 154942 91100 154948 91112
rect 138808 91072 154948 91100
rect 138808 91060 138814 91072
rect 154942 91060 154948 91072
rect 155000 91060 155006 91112
rect 224218 90992 224224 91044
rect 224276 91032 224282 91044
rect 256694 91032 256700 91044
rect 224276 91004 256700 91032
rect 224276 90992 224282 91004
rect 256694 90992 256700 91004
rect 256752 90992 256758 91044
rect 141602 89700 141608 89752
rect 141660 89740 141666 89752
rect 154942 89740 154948 89752
rect 141660 89712 154948 89740
rect 141660 89700 141666 89712
rect 154942 89700 154948 89712
rect 155000 89700 155006 89752
rect 136542 89632 136548 89684
rect 136600 89672 136606 89684
rect 147030 89672 147036 89684
rect 136600 89644 147036 89672
rect 136600 89632 136606 89644
rect 147030 89632 147036 89644
rect 147088 89632 147094 89684
rect 249334 88272 249340 88324
rect 249392 88312 249398 88324
rect 256694 88312 256700 88324
rect 249392 88284 256700 88312
rect 249392 88272 249398 88284
rect 256694 88272 256700 88284
rect 256752 88272 256758 88324
rect 135806 87320 135812 87372
rect 135864 87360 135870 87372
rect 142154 87360 142160 87372
rect 135864 87332 142160 87360
rect 135864 87320 135870 87332
rect 142154 87320 142160 87332
rect 142212 87320 142218 87372
rect 144270 86980 144276 87032
rect 144328 87020 144334 87032
rect 154942 87020 154948 87032
rect 144328 86992 154948 87020
rect 144328 86980 144334 86992
rect 154942 86980 154948 86992
rect 155000 86980 155006 87032
rect 243722 86912 243728 86964
rect 243780 86952 243786 86964
rect 256694 86952 256700 86964
rect 243780 86924 256700 86952
rect 243780 86912 243786 86924
rect 256694 86912 256700 86924
rect 256752 86912 256758 86964
rect 135254 86844 135260 86896
rect 135312 86884 135318 86896
rect 137278 86884 137284 86896
rect 135312 86856 137284 86884
rect 135312 86844 135318 86856
rect 137278 86844 137284 86856
rect 137336 86844 137342 86896
rect 137370 85552 137376 85604
rect 137428 85592 137434 85604
rect 154942 85592 154948 85604
rect 137428 85564 154948 85592
rect 137428 85552 137434 85564
rect 154942 85552 154948 85564
rect 155000 85552 155006 85604
rect 151630 84192 151636 84244
rect 151688 84232 151694 84244
rect 154942 84232 154948 84244
rect 151688 84204 154948 84232
rect 151688 84192 151694 84204
rect 154942 84192 154948 84204
rect 155000 84192 155006 84244
rect 228450 84124 228456 84176
rect 228508 84164 228514 84176
rect 256694 84164 256700 84176
rect 228508 84136 256700 84164
rect 228508 84124 228514 84136
rect 256694 84124 256700 84136
rect 256752 84124 256758 84176
rect 227162 82764 227168 82816
rect 227220 82804 227226 82816
rect 256694 82804 256700 82816
rect 227220 82776 256700 82804
rect 227220 82764 227226 82776
rect 256694 82764 256700 82776
rect 256752 82764 256758 82816
rect 136542 82220 136548 82272
rect 136600 82260 136606 82272
rect 140130 82260 140136 82272
rect 136600 82232 140136 82260
rect 136600 82220 136606 82232
rect 140130 82220 140136 82232
rect 140188 82220 140194 82272
rect 138842 81404 138848 81456
rect 138900 81444 138906 81456
rect 154942 81444 154948 81456
rect 138900 81416 154948 81444
rect 138900 81404 138906 81416
rect 154942 81404 154948 81416
rect 155000 81404 155006 81456
rect 140222 80044 140228 80096
rect 140280 80084 140286 80096
rect 154758 80084 154764 80096
rect 140280 80056 154764 80084
rect 140280 80044 140286 80056
rect 154758 80044 154764 80056
rect 154816 80044 154822 80096
rect 249150 79976 249156 80028
rect 249208 80016 249214 80028
rect 256694 80016 256700 80028
rect 249208 79988 256700 80016
rect 249208 79976 249214 79988
rect 256694 79976 256700 79988
rect 256752 79976 256758 80028
rect 136082 79704 136088 79756
rect 136140 79744 136146 79756
rect 138750 79744 138756 79756
rect 136140 79716 138756 79744
rect 136140 79704 136146 79716
rect 138750 79704 138756 79716
rect 138808 79704 138814 79756
rect 250530 78616 250536 78668
rect 250588 78656 250594 78668
rect 256694 78656 256700 78668
rect 250588 78628 256700 78656
rect 250588 78616 250594 78628
rect 256694 78616 256700 78628
rect 256752 78616 256758 78668
rect 147030 77256 147036 77308
rect 147088 77296 147094 77308
rect 154942 77296 154948 77308
rect 147088 77268 154948 77296
rect 147088 77256 147094 77268
rect 154942 77256 154948 77268
rect 155000 77256 155006 77308
rect 220262 77188 220268 77240
rect 220320 77228 220326 77240
rect 224862 77228 224868 77240
rect 220320 77200 224868 77228
rect 220320 77188 220326 77200
rect 224862 77188 224868 77200
rect 224920 77188 224926 77240
rect 235350 77188 235356 77240
rect 235408 77228 235414 77240
rect 256694 77228 256700 77240
rect 235408 77200 256700 77228
rect 235408 77188 235414 77200
rect 256694 77188 256700 77200
rect 256752 77188 256758 77240
rect 136542 77052 136548 77104
rect 136600 77092 136606 77104
rect 141602 77092 141608 77104
rect 136600 77064 141608 77092
rect 136600 77052 136606 77064
rect 141602 77052 141608 77064
rect 141660 77052 141666 77104
rect 141510 75896 141516 75948
rect 141568 75936 141574 75948
rect 154942 75936 154948 75948
rect 141568 75908 154948 75936
rect 141568 75896 141574 75908
rect 154942 75896 154948 75908
rect 155000 75896 155006 75948
rect 137278 74536 137284 74588
rect 137336 74576 137342 74588
rect 154942 74576 154948 74588
rect 137336 74548 154948 74576
rect 137336 74536 137342 74548
rect 154942 74536 154948 74548
rect 155000 74536 155006 74588
rect 244918 74468 244924 74520
rect 244976 74508 244982 74520
rect 256694 74508 256700 74520
rect 244976 74480 256700 74508
rect 244976 74468 244982 74480
rect 256694 74468 256700 74480
rect 256752 74468 256758 74520
rect 136542 73720 136548 73772
rect 136600 73760 136606 73772
rect 144270 73760 144276 73772
rect 136600 73732 144276 73760
rect 136600 73720 136606 73732
rect 144270 73720 144276 73732
rect 144328 73720 144334 73772
rect 224862 73108 224868 73160
rect 224920 73148 224926 73160
rect 256694 73148 256700 73160
rect 224920 73120 256700 73148
rect 224920 73108 224926 73120
rect 256694 73108 256700 73120
rect 256752 73108 256758 73160
rect 135714 72428 135720 72480
rect 135772 72468 135778 72480
rect 151630 72468 151636 72480
rect 135772 72440 151636 72468
rect 135772 72428 135778 72440
rect 151630 72428 151636 72440
rect 151688 72428 151694 72480
rect 151538 71748 151544 71800
rect 151596 71788 151602 71800
rect 154574 71788 154580 71800
rect 151596 71760 154580 71788
rect 151596 71748 151602 71760
rect 154574 71748 154580 71760
rect 154632 71748 154638 71800
rect 135346 71612 135352 71664
rect 135404 71652 135410 71664
rect 137370 71652 137376 71664
rect 135404 71624 137376 71652
rect 135404 71612 135410 71624
rect 137370 71612 137376 71624
rect 137428 71612 137434 71664
rect 247770 70320 247776 70372
rect 247828 70360 247834 70372
rect 256694 70360 256700 70372
rect 247828 70332 256700 70360
rect 247828 70320 247834 70332
rect 256694 70320 256700 70332
rect 256752 70320 256758 70372
rect 143074 69028 143080 69080
rect 143132 69068 143138 69080
rect 154574 69068 154580 69080
rect 143132 69040 154580 69068
rect 143132 69028 143138 69040
rect 154574 69028 154580 69040
rect 154632 69028 154638 69080
rect 229830 68960 229836 69012
rect 229888 69000 229894 69012
rect 256694 69000 256700 69012
rect 229888 68972 256700 69000
rect 229888 68960 229894 68972
rect 256694 68960 256700 68972
rect 256752 68960 256758 69012
rect 137370 68280 137376 68332
rect 137428 68320 137434 68332
rect 154942 68320 154948 68332
rect 137428 68292 154948 68320
rect 137428 68280 137434 68292
rect 154942 68280 154948 68292
rect 155000 68280 155006 68332
rect 138750 66240 138756 66292
rect 138808 66280 138814 66292
rect 154942 66280 154948 66292
rect 138808 66252 154948 66280
rect 138808 66240 138814 66252
rect 154942 66240 154948 66252
rect 155000 66240 155006 66292
rect 136082 66172 136088 66224
rect 136140 66212 136146 66224
rect 138842 66212 138848 66224
rect 136140 66184 138848 66212
rect 136140 66172 136146 66184
rect 138842 66172 138848 66184
rect 138900 66172 138906 66224
rect 140130 64880 140136 64932
rect 140188 64920 140194 64932
rect 154574 64920 154580 64932
rect 140188 64892 154580 64920
rect 140188 64880 140194 64892
rect 154574 64880 154580 64892
rect 154632 64880 154638 64932
rect 250438 64404 250444 64456
rect 250496 64444 250502 64456
rect 256694 64444 256700 64456
rect 250496 64416 256700 64444
rect 250496 64404 250502 64416
rect 256694 64404 256700 64416
rect 256752 64404 256758 64456
rect 136542 64132 136548 64184
rect 136600 64172 136606 64184
rect 140222 64172 140228 64184
rect 136600 64144 140228 64172
rect 136600 64132 136606 64144
rect 140222 64132 140228 64144
rect 140280 64132 140286 64184
rect 138842 62092 138848 62144
rect 138900 62132 138906 62144
rect 154574 62132 154580 62144
rect 138900 62104 154580 62132
rect 138900 62092 138906 62104
rect 154574 62092 154580 62104
rect 154632 62092 154638 62144
rect 135622 62024 135628 62076
rect 135680 62064 135686 62076
rect 147030 62064 147036 62076
rect 135680 62036 147036 62064
rect 135680 62024 135686 62036
rect 147030 62024 147036 62036
rect 147088 62024 147094 62076
rect 235258 62024 235264 62076
rect 235316 62064 235322 62076
rect 256694 62064 256700 62076
rect 235316 62036 256700 62064
rect 235316 62024 235322 62036
rect 256694 62024 256700 62036
rect 256752 62024 256758 62076
rect 144270 60732 144276 60784
rect 144328 60772 144334 60784
rect 154942 60772 154948 60784
rect 144328 60744 154948 60772
rect 144328 60732 144334 60744
rect 154942 60732 154948 60744
rect 155000 60732 155006 60784
rect 227070 60664 227076 60716
rect 227128 60704 227134 60716
rect 256694 60704 256700 60716
rect 227128 60676 256700 60704
rect 227128 60664 227134 60676
rect 256694 60664 256700 60676
rect 256752 60664 256758 60716
rect 147030 59372 147036 59424
rect 147088 59412 147094 59424
rect 154942 59412 154948 59424
rect 147088 59384 154948 59412
rect 147088 59372 147094 59384
rect 154942 59372 154948 59384
rect 155000 59372 155006 59424
rect 551738 59372 551744 59424
rect 551796 59412 551802 59424
rect 580074 59412 580080 59424
rect 551796 59384 580080 59412
rect 551796 59372 551802 59384
rect 580074 59372 580080 59384
rect 580132 59372 580138 59424
rect 136542 58964 136548 59016
rect 136600 59004 136606 59016
rect 141510 59004 141516 59016
rect 136600 58976 141516 59004
rect 136600 58964 136606 58976
rect 141510 58964 141516 58976
rect 141568 58964 141574 59016
rect 222838 57876 222844 57928
rect 222896 57916 222902 57928
rect 256694 57916 256700 57928
rect 222896 57888 256700 57916
rect 222896 57876 222902 57888
rect 256694 57876 256700 57888
rect 256752 57876 256758 57928
rect 141510 56584 141516 56636
rect 141568 56624 141574 56636
rect 154942 56624 154948 56636
rect 141568 56596 154948 56624
rect 141568 56584 141574 56596
rect 154942 56584 154948 56596
rect 155000 56584 155006 56636
rect 221734 56516 221740 56568
rect 221792 56556 221798 56568
rect 256694 56556 256700 56568
rect 221792 56528 256700 56556
rect 221792 56516 221798 56528
rect 256694 56516 256700 56528
rect 256752 56516 256758 56568
rect 135254 56380 135260 56432
rect 135312 56420 135318 56432
rect 137278 56420 137284 56432
rect 135312 56392 137284 56420
rect 135312 56380 135318 56392
rect 137278 56380 137284 56392
rect 137336 56380 137342 56432
rect 142982 55224 142988 55276
rect 143040 55264 143046 55276
rect 154942 55264 154948 55276
rect 143040 55236 154948 55264
rect 143040 55224 143046 55236
rect 154942 55224 154948 55236
rect 155000 55224 155006 55276
rect 242158 54476 242164 54528
rect 242216 54516 242222 54528
rect 256694 54516 256700 54528
rect 242216 54488 256700 54516
rect 242216 54476 242222 54488
rect 256694 54476 256700 54488
rect 256752 54476 256758 54528
rect 136542 53728 136548 53780
rect 136600 53768 136606 53780
rect 151538 53768 151544 53780
rect 136600 53740 151544 53768
rect 136600 53728 136606 53740
rect 151538 53728 151544 53740
rect 151596 53728 151602 53780
rect 142798 52776 142804 52828
rect 142856 52816 142862 52828
rect 142856 52788 175918 52816
rect 142856 52776 142862 52788
rect 175890 52692 175918 52788
rect 190426 52788 212534 52816
rect 175982 52720 177390 52748
rect 158438 52640 158444 52692
rect 158496 52680 158502 52692
rect 175596 52680 175602 52692
rect 158496 52652 175602 52680
rect 158496 52640 158502 52652
rect 175596 52640 175602 52652
rect 175654 52640 175660 52692
rect 175872 52640 175878 52692
rect 175930 52640 175936 52692
rect 157058 52572 157064 52624
rect 157116 52612 157122 52624
rect 175982 52612 176010 52720
rect 177252 52680 177258 52692
rect 157116 52584 176010 52612
rect 176994 52652 177258 52680
rect 157116 52572 157122 52584
rect 157150 52504 157156 52556
rect 157208 52544 157214 52556
rect 176994 52544 177022 52652
rect 177252 52640 177258 52652
rect 177310 52640 177316 52692
rect 177362 52612 177390 52720
rect 157208 52516 177022 52544
rect 177086 52584 177390 52612
rect 178466 52584 183554 52612
rect 157208 52504 157214 52516
rect 148410 52436 148416 52488
rect 148468 52476 148474 52488
rect 154942 52476 154948 52488
rect 148468 52448 154948 52476
rect 148468 52436 148474 52448
rect 154942 52436 154948 52448
rect 155000 52436 155006 52488
rect 177086 52476 177114 52584
rect 176994 52448 177114 52476
rect 176994 52420 177022 52448
rect 159910 52368 159916 52420
rect 159968 52408 159974 52420
rect 159968 52380 168374 52408
rect 159968 52368 159974 52380
rect 154546 52244 158714 52272
rect 154546 52136 154574 52244
rect 150406 52108 154574 52136
rect 158686 52136 158714 52244
rect 168346 52204 168374 52380
rect 173866 52380 176654 52408
rect 173866 52340 173894 52380
rect 172486 52312 173894 52340
rect 176626 52340 176654 52380
rect 176976 52368 176982 52420
rect 177034 52368 177040 52420
rect 176626 52312 178034 52340
rect 169726 52244 171134 52272
rect 169726 52204 169754 52244
rect 168346 52176 169754 52204
rect 171106 52204 171134 52244
rect 172486 52204 172514 52312
rect 178006 52272 178034 52312
rect 178006 52244 178402 52272
rect 171106 52176 172514 52204
rect 158686 52108 169754 52136
rect 136634 51960 136640 52012
rect 136692 52000 136698 52012
rect 150406 52000 150434 52108
rect 156598 52028 156604 52080
rect 156656 52068 156662 52080
rect 159818 52068 159824 52080
rect 156656 52040 159824 52068
rect 156656 52028 156662 52040
rect 159818 52028 159824 52040
rect 159876 52028 159882 52080
rect 169726 52068 169754 52108
rect 169726 52040 175734 52068
rect 159910 52000 159916 52012
rect 136692 51972 150434 52000
rect 154546 51972 159916 52000
rect 136692 51960 136698 51972
rect 154206 51892 154212 51944
rect 154264 51932 154270 51944
rect 154546 51932 154574 51972
rect 159910 51960 159916 51972
rect 159968 51960 159974 52012
rect 172026 51972 175044 52000
rect 172026 51944 172054 51972
rect 154264 51904 154574 51932
rect 154264 51892 154270 51904
rect 161428 51892 161434 51944
rect 161486 51892 161492 51944
rect 161796 51892 161802 51944
rect 161854 51892 161860 51944
rect 161888 51892 161894 51944
rect 161946 51892 161952 51944
rect 162992 51892 162998 51944
rect 163050 51892 163056 51944
rect 163728 51932 163734 51944
rect 163102 51904 163734 51932
rect 161060 51824 161066 51876
rect 161118 51824 161124 51876
rect 154114 51756 154120 51808
rect 154172 51796 154178 51808
rect 154172 51768 158484 51796
rect 154172 51756 154178 51768
rect 153194 51688 153200 51740
rect 153252 51728 153258 51740
rect 158456 51728 158484 51768
rect 160692 51756 160698 51808
rect 160750 51796 160756 51808
rect 161078 51796 161106 51824
rect 161446 51796 161474 51892
rect 161612 51824 161618 51876
rect 161670 51824 161676 51876
rect 160750 51768 160968 51796
rect 160750 51756 160756 51768
rect 153252 51700 157334 51728
rect 158456 51700 160692 51728
rect 153252 51688 153258 51700
rect 157306 51660 157334 51700
rect 159358 51660 159364 51672
rect 157306 51632 159364 51660
rect 159358 51620 159364 51632
rect 159416 51620 159422 51672
rect 151446 51552 151452 51604
rect 151504 51592 151510 51604
rect 151504 51564 160554 51592
rect 151504 51552 151510 51564
rect 151078 51484 151084 51536
rect 151136 51524 151142 51536
rect 159266 51524 159272 51536
rect 151136 51496 159272 51524
rect 151136 51484 151142 51496
rect 159266 51484 159272 51496
rect 159324 51484 159330 51536
rect 135990 51416 135996 51468
rect 136048 51456 136054 51468
rect 136048 51428 160232 51456
rect 136048 51416 136054 51428
rect 135898 51348 135904 51400
rect 135956 51388 135962 51400
rect 159450 51388 159456 51400
rect 135956 51360 159456 51388
rect 135956 51348 135962 51360
rect 159450 51348 159456 51360
rect 159508 51348 159514 51400
rect 160204 51332 160232 51428
rect 134702 51280 134708 51332
rect 134760 51320 134766 51332
rect 134760 51292 157334 51320
rect 134760 51280 134766 51292
rect 157306 51252 157334 51292
rect 160186 51280 160192 51332
rect 160244 51280 160250 51332
rect 160526 51320 160554 51564
rect 160664 51388 160692 51700
rect 160940 51672 160968 51768
rect 161032 51768 161106 51796
rect 161308 51768 161474 51796
rect 160922 51620 160928 51672
rect 160980 51620 160986 51672
rect 161032 51660 161060 51768
rect 161106 51660 161112 51672
rect 161032 51632 161112 51660
rect 161106 51620 161112 51632
rect 161164 51620 161170 51672
rect 161308 51536 161336 51768
rect 161630 51728 161658 51824
rect 161814 51740 161842 51892
rect 161492 51700 161658 51728
rect 161290 51484 161296 51536
rect 161348 51484 161354 51536
rect 161492 51524 161520 51700
rect 161750 51688 161756 51740
rect 161808 51700 161842 51740
rect 161808 51688 161814 51700
rect 161906 51672 161934 51892
rect 163010 51808 163038 51892
rect 162992 51756 162998 51808
rect 163050 51756 163056 51808
rect 161842 51620 161848 51672
rect 161900 51632 161934 51672
rect 161900 51620 161906 51632
rect 161934 51552 161940 51604
rect 161992 51592 161998 51604
rect 163102 51592 163130 51904
rect 163728 51892 163734 51904
rect 163786 51892 163792 51944
rect 164004 51892 164010 51944
rect 164062 51892 164068 51944
rect 164188 51892 164194 51944
rect 164246 51892 164252 51944
rect 164372 51892 164378 51944
rect 164430 51892 164436 51944
rect 164556 51892 164562 51944
rect 164614 51892 164620 51944
rect 164924 51932 164930 51944
rect 164666 51904 164930 51932
rect 163360 51824 163366 51876
rect 163418 51824 163424 51876
rect 163378 51740 163406 51824
rect 163544 51756 163550 51808
rect 163602 51756 163608 51808
rect 163378 51700 163412 51740
rect 163406 51688 163412 51700
rect 163464 51688 163470 51740
rect 161992 51564 163130 51592
rect 161992 51552 161998 51564
rect 163562 51536 163590 51756
rect 164022 51536 164050 51892
rect 164206 51672 164234 51892
rect 164280 51824 164286 51876
rect 164338 51824 164344 51876
rect 164142 51620 164148 51672
rect 164200 51632 164234 51672
rect 164200 51620 164206 51632
rect 164298 51604 164326 51824
rect 164390 51740 164418 51892
rect 164574 51808 164602 51892
rect 164510 51756 164516 51808
rect 164568 51768 164602 51808
rect 164568 51756 164574 51768
rect 164390 51700 164424 51740
rect 164418 51688 164424 51700
rect 164476 51688 164482 51740
rect 164666 51672 164694 51904
rect 164924 51892 164930 51904
rect 164982 51892 164988 51944
rect 165016 51892 165022 51944
rect 165074 51892 165080 51944
rect 165108 51892 165114 51944
rect 165166 51892 165172 51944
rect 165476 51932 165482 51944
rect 165264 51904 165482 51932
rect 164832 51824 164838 51876
rect 164890 51824 164896 51876
rect 164602 51620 164608 51672
rect 164660 51632 164694 51672
rect 164660 51620 164666 51632
rect 164234 51552 164240 51604
rect 164292 51564 164326 51604
rect 164292 51552 164298 51564
rect 161750 51524 161756 51536
rect 161492 51496 161756 51524
rect 161750 51484 161756 51496
rect 161808 51484 161814 51536
rect 163562 51496 163596 51536
rect 163590 51484 163596 51496
rect 163648 51484 163654 51536
rect 163958 51484 163964 51536
rect 164016 51496 164050 51536
rect 164850 51524 164878 51824
rect 165034 51808 165062 51892
rect 164970 51756 164976 51808
rect 165028 51768 165062 51808
rect 165028 51756 165034 51768
rect 165126 51740 165154 51892
rect 165062 51688 165068 51740
rect 165120 51700 165154 51740
rect 165120 51688 165126 51700
rect 165264 51592 165292 51904
rect 165476 51892 165482 51904
rect 165534 51892 165540 51944
rect 165660 51892 165666 51944
rect 165718 51892 165724 51944
rect 165752 51892 165758 51944
rect 165810 51892 165816 51944
rect 165936 51892 165942 51944
rect 165994 51892 166000 51944
rect 166028 51892 166034 51944
rect 166086 51892 166092 51944
rect 166212 51892 166218 51944
rect 166270 51892 166276 51944
rect 166304 51892 166310 51944
rect 166362 51892 166368 51944
rect 167132 51892 167138 51944
rect 167190 51892 167196 51944
rect 167316 51892 167322 51944
rect 167374 51892 167380 51944
rect 167408 51892 167414 51944
rect 167466 51892 167472 51944
rect 167868 51892 167874 51944
rect 167926 51892 167932 51944
rect 168052 51892 168058 51944
rect 168110 51892 168116 51944
rect 168144 51892 168150 51944
rect 168202 51892 168208 51944
rect 169156 51892 169162 51944
rect 169214 51892 169220 51944
rect 169340 51892 169346 51944
rect 169398 51892 169404 51944
rect 169616 51892 169622 51944
rect 169674 51892 169680 51944
rect 170720 51932 170726 51944
rect 170278 51904 170726 51932
rect 165522 51756 165528 51808
rect 165580 51796 165586 51808
rect 165678 51796 165706 51892
rect 165580 51768 165706 51796
rect 165580 51756 165586 51768
rect 165770 51672 165798 51892
rect 165954 51796 165982 51892
rect 165908 51768 165982 51796
rect 165908 51740 165936 51768
rect 166046 51740 166074 51892
rect 166230 51796 166258 51892
rect 166184 51768 166258 51796
rect 166184 51740 166212 51768
rect 166322 51740 166350 51892
rect 166396 51824 166402 51876
rect 166454 51824 166460 51876
rect 166580 51824 166586 51876
rect 166638 51824 166644 51876
rect 167040 51864 167046 51876
rect 167012 51824 167046 51864
rect 167098 51824 167104 51876
rect 165890 51688 165896 51740
rect 165948 51688 165954 51740
rect 165982 51688 165988 51740
rect 166040 51700 166074 51740
rect 166040 51688 166046 51700
rect 166166 51688 166172 51740
rect 166224 51688 166230 51740
rect 166258 51688 166264 51740
rect 166316 51700 166350 51740
rect 166316 51688 166322 51700
rect 166414 51672 166442 51824
rect 166488 51756 166494 51808
rect 166546 51756 166552 51808
rect 165706 51620 165712 51672
rect 165764 51632 165798 51672
rect 165764 51620 165770 51632
rect 166350 51620 166356 51672
rect 166408 51632 166442 51672
rect 166408 51620 166414 51632
rect 165172 51564 165292 51592
rect 165062 51524 165068 51536
rect 164850 51496 165068 51524
rect 164016 51484 164022 51496
rect 165062 51484 165068 51496
rect 165120 51484 165126 51536
rect 165172 51456 165200 51564
rect 166074 51552 166080 51604
rect 166132 51592 166138 51604
rect 166506 51592 166534 51756
rect 166132 51564 166534 51592
rect 166132 51552 166138 51564
rect 165614 51456 165620 51468
rect 165172 51428 165620 51456
rect 165614 51416 165620 51428
rect 165672 51416 165678 51468
rect 166442 51416 166448 51468
rect 166500 51456 166506 51468
rect 166598 51456 166626 51824
rect 167012 51740 167040 51824
rect 167150 51796 167178 51892
rect 167224 51824 167230 51876
rect 167282 51824 167288 51876
rect 167104 51768 167178 51796
rect 166994 51688 167000 51740
rect 167052 51688 167058 51740
rect 167104 51672 167132 51768
rect 167242 51740 167270 51824
rect 167178 51688 167184 51740
rect 167236 51700 167270 51740
rect 167236 51688 167242 51700
rect 167334 51672 167362 51892
rect 167426 51808 167454 51892
rect 167500 51824 167506 51876
rect 167558 51824 167564 51876
rect 167408 51756 167414 51808
rect 167466 51756 167472 51808
rect 167518 51672 167546 51824
rect 167086 51620 167092 51672
rect 167144 51620 167150 51672
rect 167334 51632 167368 51672
rect 167362 51620 167368 51632
rect 167420 51620 167426 51672
rect 167454 51620 167460 51672
rect 167512 51632 167546 51672
rect 167512 51620 167518 51632
rect 167886 51604 167914 51892
rect 168070 51740 168098 51892
rect 168006 51688 168012 51740
rect 168064 51700 168098 51740
rect 168064 51688 168070 51700
rect 168162 51672 168190 51892
rect 168236 51824 168242 51876
rect 168294 51824 168300 51876
rect 168880 51824 168886 51876
rect 168938 51824 168944 51876
rect 168098 51620 168104 51672
rect 168156 51632 168190 51672
rect 168156 51620 168162 51632
rect 168254 51604 168282 51824
rect 168696 51756 168702 51808
rect 168754 51756 168760 51808
rect 168714 51672 168742 51756
rect 168898 51740 168926 51824
rect 168834 51688 168840 51740
rect 168892 51700 168926 51740
rect 168892 51688 168898 51700
rect 168714 51632 168748 51672
rect 168742 51620 168748 51632
rect 168800 51620 168806 51672
rect 167822 51552 167828 51604
rect 167880 51564 167914 51604
rect 167880 51552 167886 51564
rect 168190 51552 168196 51604
rect 168248 51564 168282 51604
rect 168248 51552 168254 51564
rect 168374 51552 168380 51604
rect 168432 51592 168438 51604
rect 169174 51592 169202 51892
rect 169358 51672 169386 51892
rect 169634 51672 169662 51892
rect 169892 51824 169898 51876
rect 169950 51864 169956 51876
rect 169950 51836 170168 51864
rect 169950 51824 169956 51836
rect 170140 51672 170168 51836
rect 169294 51620 169300 51672
rect 169352 51632 169386 51672
rect 169352 51620 169358 51632
rect 169570 51620 169576 51672
rect 169628 51632 169662 51672
rect 169628 51620 169634 51632
rect 170122 51620 170128 51672
rect 170180 51620 170186 51672
rect 168432 51564 169202 51592
rect 168432 51552 168438 51564
rect 170278 51536 170306 51904
rect 170720 51892 170726 51904
rect 170778 51892 170784 51944
rect 172008 51892 172014 51944
rect 172066 51892 172072 51944
rect 174676 51892 174682 51944
rect 174734 51892 174740 51944
rect 170352 51824 170358 51876
rect 170410 51864 170416 51876
rect 170410 51836 170536 51864
rect 170410 51824 170416 51836
rect 170508 51604 170536 51836
rect 170904 51824 170910 51876
rect 170962 51824 170968 51876
rect 170996 51824 171002 51876
rect 171054 51824 171060 51876
rect 172284 51824 172290 51876
rect 172342 51824 172348 51876
rect 173296 51864 173302 51876
rect 173176 51836 173302 51864
rect 170582 51688 170588 51740
rect 170640 51688 170646 51740
rect 170490 51552 170496 51604
rect 170548 51552 170554 51604
rect 166902 51484 166908 51536
rect 166960 51524 166966 51536
rect 170122 51524 170128 51536
rect 166960 51496 170128 51524
rect 166960 51484 166966 51496
rect 170122 51484 170128 51496
rect 170180 51484 170186 51536
rect 170278 51496 170312 51536
rect 170306 51484 170312 51496
rect 170364 51484 170370 51536
rect 170600 51524 170628 51688
rect 170922 51672 170950 51824
rect 170858 51620 170864 51672
rect 170916 51632 170950 51672
rect 171014 51660 171042 51824
rect 171962 51660 171968 51672
rect 171014 51632 171968 51660
rect 170916 51620 170922 51632
rect 171962 51620 171968 51632
rect 172020 51620 172026 51672
rect 172146 51620 172152 51672
rect 172204 51660 172210 51672
rect 172302 51660 172330 51824
rect 172928 51756 172934 51808
rect 172986 51756 172992 51808
rect 173020 51756 173026 51808
rect 173078 51756 173084 51808
rect 172204 51632 172330 51660
rect 172946 51672 172974 51756
rect 173038 51728 173066 51756
rect 173038 51700 173112 51728
rect 173084 51672 173112 51700
rect 173176 51672 173204 51836
rect 173296 51824 173302 51836
rect 173354 51824 173360 51876
rect 173388 51756 173394 51808
rect 173446 51756 173452 51808
rect 173572 51756 173578 51808
rect 173630 51756 173636 51808
rect 173406 51672 173434 51756
rect 172946 51632 172980 51672
rect 172204 51620 172210 51632
rect 172974 51620 172980 51632
rect 173032 51620 173038 51672
rect 173066 51620 173072 51672
rect 173124 51620 173130 51672
rect 173158 51620 173164 51672
rect 173216 51620 173222 51672
rect 173342 51620 173348 51672
rect 173400 51632 173434 51672
rect 173590 51672 173618 51756
rect 173590 51632 173624 51672
rect 173400 51620 173406 51632
rect 173618 51620 173624 51632
rect 173676 51620 173682 51672
rect 174694 51660 174722 51892
rect 175016 51864 175044 51972
rect 175706 51944 175734 52040
rect 175982 51972 178034 52000
rect 175688 51892 175694 51944
rect 175746 51892 175752 51944
rect 175982 51864 176010 51972
rect 176516 51892 176522 51944
rect 176574 51932 176580 51944
rect 176574 51904 176746 51932
rect 176574 51892 176580 51904
rect 175016 51836 176010 51864
rect 176056 51824 176062 51876
rect 176114 51824 176120 51876
rect 175734 51688 175740 51740
rect 175792 51728 175798 51740
rect 176074 51728 176102 51824
rect 176608 51796 176614 51808
rect 175792 51700 176102 51728
rect 176258 51768 176614 51796
rect 175792 51688 175798 51700
rect 174694 51632 175964 51660
rect 175642 51592 175648 51604
rect 170784 51564 175648 51592
rect 170674 51524 170680 51536
rect 170600 51496 170680 51524
rect 170674 51484 170680 51496
rect 170732 51484 170738 51536
rect 166500 51428 166626 51456
rect 166500 51416 166506 51428
rect 169754 51388 169760 51400
rect 160664 51360 169760 51388
rect 169754 51348 169760 51360
rect 169812 51348 169818 51400
rect 160526 51292 169754 51320
rect 157306 51224 158714 51252
rect 135346 50940 135352 50992
rect 135404 50980 135410 50992
rect 137370 50980 137376 50992
rect 135404 50952 137376 50980
rect 135404 50940 135410 50952
rect 137370 50940 137376 50952
rect 137428 50940 137434 50992
rect 158686 50980 158714 51224
rect 159818 51212 159824 51264
rect 159876 51252 159882 51264
rect 166902 51252 166908 51264
rect 159876 51224 166908 51252
rect 159876 51212 159882 51224
rect 166902 51212 166908 51224
rect 166960 51212 166966 51264
rect 169726 51252 169754 51292
rect 170784 51252 170812 51564
rect 175642 51552 175648 51564
rect 175700 51552 175706 51604
rect 175734 51552 175740 51604
rect 175792 51552 175798 51604
rect 170950 51484 170956 51536
rect 171008 51524 171014 51536
rect 175752 51524 175780 51552
rect 171008 51496 175780 51524
rect 171008 51484 171014 51496
rect 171870 51416 171876 51468
rect 171928 51456 171934 51468
rect 175642 51456 175648 51468
rect 171928 51428 175648 51456
rect 171928 51416 171934 51428
rect 175642 51416 175648 51428
rect 175700 51416 175706 51468
rect 175936 51456 175964 51632
rect 176010 51552 176016 51604
rect 176068 51592 176074 51604
rect 176258 51592 176286 51768
rect 176608 51756 176614 51768
rect 176666 51756 176672 51808
rect 176562 51620 176568 51672
rect 176620 51660 176626 51672
rect 176718 51660 176746 51904
rect 176792 51892 176798 51944
rect 176850 51892 176856 51944
rect 176620 51632 176746 51660
rect 176620 51620 176626 51632
rect 176068 51564 176286 51592
rect 176068 51552 176074 51564
rect 176378 51552 176384 51604
rect 176436 51592 176442 51604
rect 176810 51592 176838 51892
rect 178006 51864 178034 51972
rect 178374 51944 178402 52244
rect 178356 51892 178362 51944
rect 178414 51892 178420 51944
rect 178466 51864 178494 52584
rect 183526 52476 183554 52584
rect 183526 52448 184934 52476
rect 184906 52272 184934 52448
rect 190426 52340 190454 52788
rect 212506 52748 212534 52788
rect 216674 52776 216680 52828
rect 216732 52816 216738 52828
rect 216732 52788 220814 52816
rect 216732 52776 216738 52788
rect 216030 52748 216036 52760
rect 202846 52720 209774 52748
rect 212506 52720 216036 52748
rect 195992 52652 198734 52680
rect 195992 52454 196020 52652
rect 195716 52426 196020 52454
rect 198706 52476 198734 52652
rect 202846 52476 202874 52720
rect 209746 52544 209774 52720
rect 216030 52708 216036 52720
rect 216088 52708 216094 52760
rect 211126 52652 212534 52680
rect 211126 52544 211154 52652
rect 212506 52612 212534 52652
rect 212506 52584 219434 52612
rect 209746 52516 211154 52544
rect 198706 52448 202874 52476
rect 219406 52476 219434 52584
rect 220786 52544 220814 52788
rect 255866 52544 255872 52556
rect 220786 52516 255872 52544
rect 255866 52504 255872 52516
rect 255924 52504 255930 52556
rect 253382 52476 253388 52488
rect 219406 52448 253388 52476
rect 253382 52436 253388 52448
rect 253440 52436 253446 52488
rect 195716 52408 195744 52426
rect 194428 52380 195744 52408
rect 194428 52340 194456 52380
rect 200252 52368 200258 52420
rect 200310 52408 200316 52420
rect 200310 52380 209682 52408
rect 200310 52368 200316 52380
rect 186286 52312 190454 52340
rect 193554 52312 194456 52340
rect 186286 52272 186314 52312
rect 184906 52244 186314 52272
rect 189230 52244 193398 52272
rect 182772 52028 182778 52080
rect 182830 52028 182836 52080
rect 184336 52028 184342 52080
rect 184394 52028 184400 52080
rect 188108 52028 188114 52080
rect 188166 52028 188172 52080
rect 182790 52000 182818 52028
rect 181226 51972 181990 52000
rect 182790 51972 183048 52000
rect 181226 51944 181254 51972
rect 179000 51892 179006 51944
rect 179058 51892 179064 51944
rect 179092 51892 179098 51944
rect 179150 51892 179156 51944
rect 179368 51892 179374 51944
rect 179426 51932 179432 51944
rect 179426 51904 179736 51932
rect 179426 51892 179432 51904
rect 178006 51836 178494 51864
rect 178816 51824 178822 51876
rect 178874 51824 178880 51876
rect 179018 51864 179046 51892
rect 178926 51836 179046 51864
rect 177068 51756 177074 51808
rect 177126 51756 177132 51808
rect 178834 51796 178862 51824
rect 177638 51768 178862 51796
rect 176436 51564 176838 51592
rect 177086 51604 177114 51756
rect 177086 51564 177120 51604
rect 176436 51552 176442 51564
rect 177114 51552 177120 51564
rect 177172 51552 177178 51604
rect 176102 51484 176108 51536
rect 176160 51524 176166 51536
rect 177638 51524 177666 51768
rect 178494 51552 178500 51604
rect 178552 51592 178558 51604
rect 178926 51592 178954 51836
rect 179110 51740 179138 51892
rect 179276 51824 179282 51876
rect 179334 51824 179340 51876
rect 179460 51824 179466 51876
rect 179518 51824 179524 51876
rect 179552 51824 179558 51876
rect 179610 51864 179616 51876
rect 179610 51824 179644 51864
rect 179046 51688 179052 51740
rect 179104 51700 179138 51740
rect 179104 51688 179110 51700
rect 178552 51564 178954 51592
rect 178552 51552 178558 51564
rect 176160 51496 177666 51524
rect 176160 51484 176166 51496
rect 178954 51456 178960 51468
rect 175936 51428 178960 51456
rect 178954 51416 178960 51428
rect 179012 51416 179018 51468
rect 173434 51348 173440 51400
rect 173492 51388 173498 51400
rect 175734 51388 175740 51400
rect 173492 51360 175740 51388
rect 173492 51348 173498 51360
rect 175734 51348 175740 51360
rect 175792 51348 175798 51400
rect 179294 51388 179322 51824
rect 179478 51672 179506 51824
rect 179616 51740 179644 51824
rect 179598 51688 179604 51740
rect 179656 51688 179662 51740
rect 179414 51620 179420 51672
rect 179472 51632 179506 51672
rect 179472 51620 179478 51632
rect 179506 51552 179512 51604
rect 179564 51592 179570 51604
rect 179708 51592 179736 51904
rect 180104 51892 180110 51944
rect 180162 51892 180168 51944
rect 180196 51892 180202 51944
rect 180254 51892 180260 51944
rect 180472 51892 180478 51944
rect 180530 51892 180536 51944
rect 181116 51892 181122 51944
rect 181174 51892 181180 51944
rect 181208 51892 181214 51944
rect 181266 51892 181272 51944
rect 180012 51824 180018 51876
rect 180070 51824 180076 51876
rect 179564 51564 179736 51592
rect 179564 51552 179570 51564
rect 177270 51360 179322 51388
rect 180030 51400 180058 51824
rect 180122 51456 180150 51892
rect 180214 51524 180242 51892
rect 180490 51808 180518 51892
rect 180564 51824 180570 51876
rect 180622 51824 180628 51876
rect 180426 51756 180432 51808
rect 180484 51768 180518 51808
rect 180484 51756 180490 51768
rect 180582 51740 180610 51824
rect 180656 51756 180662 51808
rect 180714 51756 180720 51808
rect 180840 51756 180846 51808
rect 180898 51756 180904 51808
rect 180518 51688 180524 51740
rect 180576 51700 180610 51740
rect 180576 51688 180582 51700
rect 180674 51672 180702 51756
rect 180610 51620 180616 51672
rect 180668 51632 180702 51672
rect 180668 51620 180674 51632
rect 180334 51524 180340 51536
rect 180214 51496 180340 51524
rect 180334 51484 180340 51496
rect 180392 51484 180398 51536
rect 180858 51524 180886 51756
rect 181134 51672 181162 51892
rect 181576 51864 181582 51876
rect 181272 51836 181582 51864
rect 181272 51808 181300 51836
rect 181576 51824 181582 51836
rect 181634 51824 181640 51876
rect 181254 51756 181260 51808
rect 181312 51756 181318 51808
rect 181852 51796 181858 51808
rect 181456 51768 181858 51796
rect 181134 51632 181168 51672
rect 181162 51620 181168 51632
rect 181220 51620 181226 51672
rect 181456 51536 181484 51768
rect 181852 51756 181858 51768
rect 181910 51756 181916 51808
rect 181622 51688 181628 51740
rect 181680 51688 181686 51740
rect 181162 51524 181168 51536
rect 180858 51496 181168 51524
rect 181162 51484 181168 51496
rect 181220 51484 181226 51536
rect 181438 51484 181444 51536
rect 181496 51484 181502 51536
rect 181640 51524 181668 51688
rect 181714 51524 181720 51536
rect 181640 51496 181720 51524
rect 181714 51484 181720 51496
rect 181772 51484 181778 51536
rect 180794 51456 180800 51468
rect 180122 51428 180800 51456
rect 180794 51416 180800 51428
rect 180852 51416 180858 51468
rect 180030 51360 180064 51400
rect 173710 51280 173716 51332
rect 173768 51320 173774 51332
rect 177270 51320 177298 51360
rect 180058 51348 180064 51360
rect 180116 51348 180122 51400
rect 181070 51348 181076 51400
rect 181128 51388 181134 51400
rect 181962 51388 181990 51972
rect 182220 51892 182226 51944
rect 182278 51892 182284 51944
rect 182312 51892 182318 51944
rect 182370 51892 182376 51944
rect 182496 51892 182502 51944
rect 182554 51892 182560 51944
rect 182588 51892 182594 51944
rect 182646 51892 182652 51944
rect 182680 51892 182686 51944
rect 182738 51932 182744 51944
rect 182738 51892 182772 51932
rect 182864 51892 182870 51944
rect 182922 51932 182928 51944
rect 182922 51892 182956 51932
rect 182128 51824 182134 51876
rect 182186 51824 182192 51876
rect 182146 51536 182174 51824
rect 182238 51672 182266 51892
rect 182330 51808 182358 51892
rect 182330 51768 182364 51808
rect 182358 51756 182364 51768
rect 182416 51756 182422 51808
rect 182514 51740 182542 51892
rect 182606 51864 182634 51892
rect 182606 51836 182680 51864
rect 182514 51700 182548 51740
rect 182542 51688 182548 51700
rect 182600 51688 182606 51740
rect 182238 51632 182272 51672
rect 182266 51620 182272 51632
rect 182324 51620 182330 51672
rect 182652 51604 182680 51836
rect 182744 51672 182772 51892
rect 182726 51620 182732 51672
rect 182784 51620 182790 51672
rect 182928 51604 182956 51892
rect 182634 51552 182640 51604
rect 182692 51552 182698 51604
rect 182910 51552 182916 51604
rect 182968 51552 182974 51604
rect 183020 51536 183048 51972
rect 183140 51892 183146 51944
rect 183198 51892 183204 51944
rect 183232 51892 183238 51944
rect 183290 51892 183296 51944
rect 183324 51892 183330 51944
rect 183382 51932 183388 51944
rect 183382 51892 183416 51932
rect 183692 51892 183698 51944
rect 183750 51892 183756 51944
rect 183876 51892 183882 51944
rect 183934 51892 183940 51944
rect 183968 51892 183974 51944
rect 184026 51892 184032 51944
rect 184060 51892 184066 51944
rect 184118 51892 184124 51944
rect 184244 51892 184250 51944
rect 184302 51892 184308 51944
rect 184354 51932 184382 52028
rect 185182 51972 185716 52000
rect 185182 51944 185210 51972
rect 184354 51904 184520 51932
rect 183158 51740 183186 51892
rect 183250 51864 183278 51892
rect 183250 51836 183324 51864
rect 183296 51808 183324 51836
rect 183278 51756 183284 51808
rect 183336 51756 183342 51808
rect 183158 51700 183192 51740
rect 183186 51688 183192 51700
rect 183244 51688 183250 51740
rect 182082 51484 182088 51536
rect 182140 51496 182174 51536
rect 182140 51484 182146 51496
rect 183002 51484 183008 51536
rect 183060 51484 183066 51536
rect 181128 51360 181990 51388
rect 181128 51348 181134 51360
rect 182726 51348 182732 51400
rect 182784 51388 182790 51400
rect 183388 51388 183416 51892
rect 183710 51808 183738 51892
rect 183646 51756 183652 51808
rect 183704 51768 183738 51808
rect 183704 51756 183710 51768
rect 183894 51672 183922 51892
rect 183986 51740 184014 51892
rect 184078 51796 184106 51892
rect 184262 51808 184290 51892
rect 184382 51824 184388 51876
rect 184440 51824 184446 51876
rect 184078 51768 184152 51796
rect 184124 51740 184152 51768
rect 184198 51756 184204 51808
rect 184256 51768 184290 51808
rect 184256 51756 184262 51768
rect 184400 51740 184428 51824
rect 183986 51700 184020 51740
rect 184014 51688 184020 51700
rect 184072 51688 184078 51740
rect 184106 51688 184112 51740
rect 184164 51688 184170 51740
rect 184382 51688 184388 51740
rect 184440 51688 184446 51740
rect 183894 51632 183928 51672
rect 183922 51620 183928 51632
rect 183980 51620 183986 51672
rect 184290 51620 184296 51672
rect 184348 51660 184354 51672
rect 184492 51660 184520 51904
rect 184888 51892 184894 51944
rect 184946 51892 184952 51944
rect 185164 51892 185170 51944
rect 185222 51892 185228 51944
rect 185256 51892 185262 51944
rect 185314 51892 185320 51944
rect 185348 51892 185354 51944
rect 185406 51892 185412 51944
rect 185440 51892 185446 51944
rect 185498 51892 185504 51944
rect 184348 51632 184520 51660
rect 184348 51620 184354 51632
rect 184906 51536 184934 51892
rect 185274 51864 185302 51892
rect 185228 51836 185302 51864
rect 185072 51796 185078 51808
rect 185044 51756 185078 51796
rect 185130 51756 185136 51808
rect 185044 51672 185072 51756
rect 185228 51740 185256 51836
rect 185366 51796 185394 51892
rect 185320 51768 185394 51796
rect 185320 51740 185348 51768
rect 185458 51740 185486 51892
rect 185210 51688 185216 51740
rect 185268 51688 185274 51740
rect 185302 51688 185308 51740
rect 185360 51688 185366 51740
rect 185394 51688 185400 51740
rect 185452 51700 185486 51740
rect 185452 51688 185458 51700
rect 185026 51620 185032 51672
rect 185084 51620 185090 51672
rect 185118 51620 185124 51672
rect 185176 51660 185182 51672
rect 185578 51660 185584 51672
rect 185176 51632 185584 51660
rect 185176 51620 185182 51632
rect 185578 51620 185584 51632
rect 185636 51620 185642 51672
rect 184842 51484 184848 51536
rect 184900 51496 184934 51536
rect 184900 51484 184906 51496
rect 185578 51484 185584 51536
rect 185636 51524 185642 51536
rect 185688 51524 185716 51972
rect 185900 51892 185906 51944
rect 185958 51892 185964 51944
rect 186268 51932 186274 51944
rect 186010 51904 186274 51932
rect 185808 51824 185814 51876
rect 185866 51824 185872 51876
rect 185636 51496 185716 51524
rect 185636 51484 185642 51496
rect 185826 51468 185854 51824
rect 185762 51416 185768 51468
rect 185820 51428 185854 51468
rect 185820 51416 185826 51428
rect 185918 51400 185946 51892
rect 186010 51536 186038 51904
rect 186268 51892 186274 51904
rect 186326 51892 186332 51944
rect 186544 51892 186550 51944
rect 186602 51932 186608 51944
rect 186602 51904 187142 51932
rect 186602 51892 186608 51904
rect 186084 51824 186090 51876
rect 186142 51824 186148 51876
rect 186360 51824 186366 51876
rect 186418 51824 186424 51876
rect 186820 51824 186826 51876
rect 186878 51824 186884 51876
rect 187114 51864 187142 51904
rect 187464 51892 187470 51944
rect 187522 51892 187528 51944
rect 187832 51892 187838 51944
rect 187890 51892 187896 51944
rect 188126 51932 188154 52028
rect 189230 51944 189258 52244
rect 189488 52164 189494 52216
rect 189546 52204 189552 52216
rect 189546 52176 191834 52204
rect 189546 52164 189552 52176
rect 191806 52136 191834 52176
rect 191806 52108 193306 52136
rect 190408 52028 190414 52080
rect 190466 52028 190472 52080
rect 192248 52028 192254 52080
rect 192306 52028 192312 52080
rect 188126 51904 188890 51932
rect 187114 51836 187188 51864
rect 186102 51660 186130 51824
rect 186222 51660 186228 51672
rect 186102 51632 186228 51660
rect 186222 51620 186228 51632
rect 186280 51620 186286 51672
rect 186378 51660 186406 51824
rect 186498 51660 186504 51672
rect 186378 51632 186504 51660
rect 186498 51620 186504 51632
rect 186556 51620 186562 51672
rect 186838 51660 186866 51824
rect 187160 51672 187188 51836
rect 187280 51824 187286 51876
rect 187338 51824 187344 51876
rect 187372 51824 187378 51876
rect 187430 51824 187436 51876
rect 186958 51660 186964 51672
rect 186838 51632 186964 51660
rect 186958 51620 186964 51632
rect 187016 51620 187022 51672
rect 187142 51620 187148 51672
rect 187200 51620 187206 51672
rect 186314 51552 186320 51604
rect 186372 51592 186378 51604
rect 187298 51592 187326 51824
rect 187390 51672 187418 51824
rect 187482 51728 187510 51892
rect 187482 51700 187556 51728
rect 187528 51672 187556 51700
rect 187390 51632 187424 51672
rect 187418 51620 187424 51632
rect 187476 51620 187482 51672
rect 187510 51620 187516 51672
rect 187568 51620 187574 51672
rect 186372 51564 187326 51592
rect 186372 51552 186378 51564
rect 186010 51496 186044 51536
rect 186038 51484 186044 51496
rect 186096 51484 186102 51536
rect 186590 51484 186596 51536
rect 186648 51524 186654 51536
rect 186774 51524 186780 51536
rect 186648 51496 186780 51524
rect 186648 51484 186654 51496
rect 186774 51484 186780 51496
rect 186832 51484 186838 51536
rect 187694 51484 187700 51536
rect 187752 51524 187758 51536
rect 187850 51524 187878 51892
rect 188200 51824 188206 51876
rect 188258 51824 188264 51876
rect 188292 51824 188298 51876
rect 188350 51824 188356 51876
rect 188476 51824 188482 51876
rect 188534 51824 188540 51876
rect 187752 51496 187878 51524
rect 187752 51484 187758 51496
rect 187970 51484 187976 51536
rect 188028 51524 188034 51536
rect 188218 51524 188246 51824
rect 188310 51672 188338 51824
rect 188310 51632 188344 51672
rect 188338 51620 188344 51632
rect 188396 51620 188402 51672
rect 188028 51496 188246 51524
rect 188028 51484 188034 51496
rect 182784 51360 183416 51388
rect 184676 51360 184888 51388
rect 182784 51348 182790 51360
rect 173768 51292 177298 51320
rect 173768 51280 173774 51292
rect 178954 51280 178960 51332
rect 179012 51320 179018 51332
rect 180886 51320 180892 51332
rect 179012 51292 180892 51320
rect 179012 51280 179018 51292
rect 180886 51280 180892 51292
rect 180944 51280 180950 51332
rect 184676 51320 184704 51360
rect 180996 51292 184704 51320
rect 184860 51320 184888 51360
rect 185854 51348 185860 51400
rect 185912 51360 185946 51400
rect 185912 51348 185918 51360
rect 187970 51348 187976 51400
rect 188028 51388 188034 51400
rect 188494 51388 188522 51824
rect 188660 51756 188666 51808
rect 188718 51756 188724 51808
rect 188028 51360 188522 51388
rect 188028 51348 188034 51360
rect 184860 51292 188384 51320
rect 169726 51224 170812 51252
rect 175090 51212 175096 51264
rect 175148 51252 175154 51264
rect 180996 51252 181024 51292
rect 188356 51252 188384 51292
rect 188430 51280 188436 51332
rect 188488 51320 188494 51332
rect 188678 51320 188706 51756
rect 188862 51468 188890 51904
rect 189212 51892 189218 51944
rect 189270 51892 189276 51944
rect 190132 51932 190138 51944
rect 189368 51904 190138 51932
rect 188936 51824 188942 51876
rect 188994 51824 189000 51876
rect 188954 51524 188982 51824
rect 189166 51524 189172 51536
rect 188954 51496 189172 51524
rect 189166 51484 189172 51496
rect 189224 51484 189230 51536
rect 189258 51484 189264 51536
rect 189316 51524 189322 51536
rect 189368 51524 189396 51904
rect 190132 51892 190138 51904
rect 190190 51892 190196 51944
rect 190224 51892 190230 51944
rect 190282 51892 190288 51944
rect 189580 51864 189586 51876
rect 189460 51836 189586 51864
rect 189460 51672 189488 51836
rect 189580 51824 189586 51836
rect 189638 51824 189644 51876
rect 189764 51824 189770 51876
rect 189822 51824 189828 51876
rect 189782 51728 189810 51824
rect 190242 51808 190270 51892
rect 190178 51756 190184 51808
rect 190236 51768 190270 51808
rect 190236 51756 190242 51768
rect 189644 51700 189810 51728
rect 189442 51620 189448 51672
rect 189500 51620 189506 51672
rect 189316 51496 189396 51524
rect 189644 51524 189672 51700
rect 189718 51620 189724 51672
rect 189776 51660 189782 51672
rect 190426 51660 190454 52028
rect 191328 51932 191334 51944
rect 189776 51632 190454 51660
rect 190564 51904 191334 51932
rect 189776 51620 189782 51632
rect 190564 51536 190592 51904
rect 191328 51892 191334 51904
rect 191386 51892 191392 51944
rect 191604 51932 191610 51944
rect 191438 51904 191610 51932
rect 190776 51824 190782 51876
rect 190834 51824 190840 51876
rect 190868 51824 190874 51876
rect 190926 51824 190932 51876
rect 191236 51824 191242 51876
rect 191294 51824 191300 51876
rect 190362 51524 190368 51536
rect 189644 51496 190368 51524
rect 189316 51484 189322 51496
rect 190362 51484 190368 51496
rect 190420 51484 190426 51536
rect 190546 51484 190552 51536
rect 190604 51484 190610 51536
rect 190794 51524 190822 51824
rect 190748 51496 190822 51524
rect 190886 51524 190914 51824
rect 191098 51524 191104 51536
rect 190886 51496 191104 51524
rect 188862 51428 188896 51468
rect 188890 51416 188896 51428
rect 188948 51416 188954 51468
rect 190748 51388 190776 51496
rect 191098 51484 191104 51496
rect 191156 51484 191162 51536
rect 190822 51416 190828 51468
rect 190880 51456 190886 51468
rect 191254 51456 191282 51824
rect 191438 51468 191466 51904
rect 191604 51892 191610 51904
rect 191662 51892 191668 51944
rect 192064 51892 192070 51944
rect 192122 51892 192128 51944
rect 191696 51864 191702 51876
rect 191668 51824 191702 51864
rect 191754 51824 191760 51876
rect 191668 51536 191696 51824
rect 191788 51796 191794 51808
rect 191760 51756 191794 51796
rect 191846 51756 191852 51808
rect 191880 51756 191886 51808
rect 191938 51756 191944 51808
rect 191972 51756 191978 51808
rect 192030 51756 192036 51808
rect 191760 51604 191788 51756
rect 191898 51604 191926 51756
rect 191742 51552 191748 51604
rect 191800 51552 191806 51604
rect 191834 51552 191840 51604
rect 191892 51564 191926 51604
rect 191990 51604 192018 51756
rect 192082 51740 192110 51892
rect 192082 51700 192116 51740
rect 192110 51688 192116 51700
rect 192168 51688 192174 51740
rect 191990 51564 192024 51604
rect 191892 51552 191898 51564
rect 192018 51552 192024 51564
rect 192076 51552 192082 51604
rect 191650 51484 191656 51536
rect 191708 51484 191714 51536
rect 190880 51428 191282 51456
rect 190880 51416 190886 51428
rect 191374 51416 191380 51468
rect 191432 51428 191466 51468
rect 191432 51416 191438 51428
rect 191926 51416 191932 51468
rect 191984 51456 191990 51468
rect 192266 51456 192294 52028
rect 192616 51892 192622 51944
rect 192674 51892 192680 51944
rect 192634 51808 192662 51892
rect 193168 51824 193174 51876
rect 193226 51824 193232 51876
rect 192570 51756 192576 51808
rect 192628 51768 192662 51808
rect 192628 51756 192634 51768
rect 192938 51484 192944 51536
rect 192996 51524 193002 51536
rect 193186 51524 193214 51824
rect 192996 51496 193214 51524
rect 193278 51524 193306 52108
rect 193370 51728 193398 52244
rect 193444 51824 193450 51876
rect 193502 51864 193508 51876
rect 193554 51864 193582 52312
rect 209654 52272 209682 52380
rect 216030 52368 216036 52420
rect 216088 52408 216094 52420
rect 216088 52380 220814 52408
rect 216088 52368 216094 52380
rect 216214 52340 216220 52352
rect 209746 52312 216220 52340
rect 209746 52272 209774 52312
rect 216214 52300 216220 52312
rect 216272 52300 216278 52352
rect 220786 52272 220814 52380
rect 197648 52244 198274 52272
rect 197648 52204 197676 52244
rect 197326 52176 197676 52204
rect 198246 52204 198274 52244
rect 200086 52244 202874 52272
rect 209654 52244 209774 52272
rect 212506 52244 219434 52272
rect 220786 52244 224954 52272
rect 200086 52204 200114 52244
rect 198246 52176 198642 52204
rect 197326 52136 197354 52176
rect 193502 51836 193582 51864
rect 193784 52108 197354 52136
rect 198614 52136 198642 52176
rect 198706 52176 200114 52204
rect 202846 52204 202874 52244
rect 212506 52204 212534 52244
rect 202846 52176 212534 52204
rect 198706 52136 198734 52176
rect 214420 52164 214426 52216
rect 214478 52204 214484 52216
rect 216306 52204 216312 52216
rect 214478 52176 216312 52204
rect 214478 52164 214484 52176
rect 216306 52164 216312 52176
rect 216364 52164 216370 52216
rect 219406 52204 219434 52244
rect 219406 52176 222194 52204
rect 216122 52136 216128 52148
rect 198614 52108 198734 52136
rect 210850 52108 216128 52136
rect 193502 51824 193508 51836
rect 193784 51728 193812 52108
rect 194060 52040 201218 52068
rect 194060 52000 194088 52040
rect 193370 51700 193812 51728
rect 193876 51972 194088 52000
rect 195072 51972 195606 52000
rect 193876 51524 193904 51972
rect 193996 51932 194002 51944
rect 193278 51496 193904 51524
rect 193968 51892 194002 51932
rect 194054 51892 194060 51944
rect 194088 51892 194094 51944
rect 194146 51892 194152 51944
rect 194180 51892 194186 51944
rect 194238 51892 194244 51944
rect 194272 51892 194278 51944
rect 194330 51932 194336 51944
rect 194330 51904 194594 51932
rect 194330 51892 194336 51904
rect 192996 51484 193002 51496
rect 191984 51428 192294 51456
rect 191984 51416 191990 51428
rect 191558 51388 191564 51400
rect 190748 51360 191564 51388
rect 191558 51348 191564 51360
rect 191616 51348 191622 51400
rect 193968 51388 193996 51892
rect 194106 51864 194134 51892
rect 194060 51836 194134 51864
rect 194060 51740 194088 51836
rect 194198 51740 194226 51892
rect 194364 51824 194370 51876
rect 194422 51824 194428 51876
rect 194456 51824 194462 51876
rect 194514 51824 194520 51876
rect 194042 51688 194048 51740
rect 194100 51688 194106 51740
rect 194134 51688 194140 51740
rect 194192 51700 194226 51740
rect 194382 51728 194410 51824
rect 194336 51700 194410 51728
rect 194192 51688 194198 51700
rect 194336 51604 194364 51700
rect 194474 51604 194502 51824
rect 194318 51552 194324 51604
rect 194376 51552 194382 51604
rect 194410 51552 194416 51604
rect 194468 51564 194502 51604
rect 194468 51552 194474 51564
rect 194566 51536 194594 51904
rect 194732 51892 194738 51944
rect 194790 51892 194796 51944
rect 194916 51892 194922 51944
rect 194974 51892 194980 51944
rect 194750 51808 194778 51892
rect 194750 51768 194784 51808
rect 194778 51756 194784 51768
rect 194836 51756 194842 51808
rect 194934 51592 194962 51892
rect 195072 51672 195100 51972
rect 195578 51944 195606 51972
rect 197326 51972 198274 52000
rect 197326 51944 197354 51972
rect 195192 51892 195198 51944
rect 195250 51892 195256 51944
rect 195284 51892 195290 51944
rect 195342 51892 195348 51944
rect 195376 51892 195382 51944
rect 195434 51892 195440 51944
rect 195560 51892 195566 51944
rect 195618 51892 195624 51944
rect 196020 51892 196026 51944
rect 196078 51892 196084 51944
rect 196204 51892 196210 51944
rect 196262 51892 196268 51944
rect 196480 51892 196486 51944
rect 196538 51892 196544 51944
rect 196848 51892 196854 51944
rect 196906 51892 196912 51944
rect 197216 51892 197222 51944
rect 197274 51892 197280 51944
rect 197308 51892 197314 51944
rect 197366 51892 197372 51944
rect 197676 51932 197682 51944
rect 197648 51892 197682 51932
rect 197734 51892 197740 51944
rect 198044 51892 198050 51944
rect 198102 51892 198108 51944
rect 195054 51620 195060 51672
rect 195112 51620 195118 51672
rect 195210 51660 195238 51892
rect 195302 51740 195330 51892
rect 195394 51796 195422 51892
rect 195652 51864 195658 51876
rect 195624 51824 195658 51864
rect 195710 51824 195716 51876
rect 195394 51768 195560 51796
rect 195302 51700 195336 51740
rect 195330 51688 195336 51700
rect 195388 51688 195394 51740
rect 195422 51660 195428 51672
rect 195210 51632 195428 51660
rect 195422 51620 195428 51632
rect 195480 51620 195486 51672
rect 195532 51604 195560 51768
rect 195624 51672 195652 51824
rect 195606 51620 195612 51672
rect 195664 51620 195670 51672
rect 195238 51592 195244 51604
rect 194934 51564 195244 51592
rect 195238 51552 195244 51564
rect 195296 51552 195302 51604
rect 195514 51552 195520 51604
rect 195572 51552 195578 51604
rect 196038 51536 196066 51892
rect 194566 51496 194600 51536
rect 194594 51484 194600 51496
rect 194652 51484 194658 51536
rect 195974 51484 195980 51536
rect 196032 51496 196066 51536
rect 196032 51484 196038 51496
rect 196222 51456 196250 51892
rect 196498 51672 196526 51892
rect 196498 51632 196532 51672
rect 196526 51620 196532 51632
rect 196584 51620 196590 51672
rect 196866 51660 196894 51892
rect 197234 51740 197262 51892
rect 197400 51824 197406 51876
rect 197458 51824 197464 51876
rect 197492 51824 197498 51876
rect 197550 51824 197556 51876
rect 197418 51740 197446 51824
rect 197234 51700 197268 51740
rect 197262 51688 197268 51700
rect 197320 51688 197326 51740
rect 197354 51688 197360 51740
rect 197412 51700 197446 51740
rect 197412 51688 197418 51700
rect 196636 51632 196894 51660
rect 196636 51524 196664 51632
rect 197510 51604 197538 51824
rect 196710 51552 196716 51604
rect 196768 51592 196774 51604
rect 197170 51592 197176 51604
rect 196768 51564 197176 51592
rect 196768 51552 196774 51564
rect 197170 51552 197176 51564
rect 197228 51552 197234 51604
rect 197510 51564 197544 51604
rect 197538 51552 197544 51564
rect 197596 51552 197602 51604
rect 196802 51524 196808 51536
rect 196636 51496 196808 51524
rect 196802 51484 196808 51496
rect 196860 51484 196866 51536
rect 196894 51484 196900 51536
rect 196952 51524 196958 51536
rect 197648 51524 197676 51892
rect 197860 51824 197866 51876
rect 197918 51824 197924 51876
rect 197722 51552 197728 51604
rect 197780 51592 197786 51604
rect 197878 51592 197906 51824
rect 197952 51756 197958 51808
rect 198010 51756 198016 51808
rect 197970 51672 197998 51756
rect 198062 51728 198090 51892
rect 198062 51700 198136 51728
rect 197970 51632 198004 51672
rect 197998 51620 198004 51632
rect 198056 51620 198062 51672
rect 197780 51564 197906 51592
rect 197780 51552 197786 51564
rect 196952 51496 197676 51524
rect 196952 51484 196958 51496
rect 197814 51484 197820 51536
rect 197872 51524 197878 51536
rect 198108 51524 198136 51700
rect 198246 51604 198274 51972
rect 199056 51892 199062 51944
rect 199114 51892 199120 51944
rect 200224 51904 200850 51932
rect 198780 51824 198786 51876
rect 198838 51824 198844 51876
rect 198504 51756 198510 51808
rect 198562 51756 198568 51808
rect 198522 51672 198550 51756
rect 198798 51672 198826 51824
rect 198458 51620 198464 51672
rect 198516 51632 198550 51672
rect 198516 51620 198522 51632
rect 198734 51620 198740 51672
rect 198792 51632 198826 51672
rect 198792 51620 198798 51632
rect 198246 51564 198280 51604
rect 198274 51552 198280 51564
rect 198332 51552 198338 51604
rect 198642 51552 198648 51604
rect 198700 51552 198706 51604
rect 199074 51592 199102 51892
rect 199332 51824 199338 51876
rect 199390 51824 199396 51876
rect 199516 51824 199522 51876
rect 199574 51824 199580 51876
rect 199792 51824 199798 51876
rect 199850 51824 199856 51876
rect 199976 51824 199982 51876
rect 200034 51824 200040 51876
rect 200068 51824 200074 51876
rect 200126 51824 200132 51876
rect 199194 51620 199200 51672
rect 199252 51660 199258 51672
rect 199350 51660 199378 51824
rect 199252 51632 199378 51660
rect 199534 51660 199562 51824
rect 199810 51672 199838 51824
rect 199994 51672 200022 51824
rect 199654 51660 199660 51672
rect 199534 51632 199660 51660
rect 199252 51620 199258 51632
rect 199654 51620 199660 51632
rect 199712 51620 199718 51672
rect 199810 51632 199844 51672
rect 199838 51620 199844 51632
rect 199896 51620 199902 51672
rect 199930 51620 199936 51672
rect 199988 51632 200022 51672
rect 199988 51620 199994 51632
rect 199378 51592 199384 51604
rect 199074 51564 199384 51592
rect 199378 51552 199384 51564
rect 199436 51552 199442 51604
rect 198660 51524 198688 51552
rect 197872 51496 198136 51524
rect 198568 51496 198688 51524
rect 197872 51484 197878 51496
rect 198568 51468 198596 51496
rect 199010 51484 199016 51536
rect 199068 51524 199074 51536
rect 200086 51524 200114 51824
rect 200224 51672 200252 51904
rect 200712 51824 200718 51876
rect 200770 51824 200776 51876
rect 200822 51864 200850 51904
rect 201080 51864 201086 51876
rect 200822 51836 201086 51864
rect 201080 51824 201086 51836
rect 201138 51824 201144 51876
rect 200206 51620 200212 51672
rect 200264 51620 200270 51672
rect 199068 51496 200114 51524
rect 200730 51524 200758 51824
rect 201190 51796 201218 52040
rect 205790 52040 206830 52068
rect 205790 51944 205818 52040
rect 201724 51892 201730 51944
rect 201782 51892 201788 51944
rect 202184 51892 202190 51944
rect 202242 51892 202248 51944
rect 203012 51892 203018 51944
rect 203070 51932 203076 51944
rect 203070 51904 204300 51932
rect 203070 51892 203076 51904
rect 201742 51808 201770 51892
rect 202000 51824 202006 51876
rect 202058 51824 202064 51876
rect 201052 51768 201218 51796
rect 201052 51604 201080 51768
rect 201632 51756 201638 51808
rect 201690 51756 201696 51808
rect 201742 51768 201776 51808
rect 201770 51756 201776 51768
rect 201828 51756 201834 51808
rect 201650 51672 201678 51756
rect 201650 51632 201684 51672
rect 201678 51620 201684 51632
rect 201736 51620 201742 51672
rect 201862 51620 201868 51672
rect 201920 51660 201926 51672
rect 202018 51660 202046 51824
rect 201920 51632 202046 51660
rect 202202 51672 202230 51892
rect 202644 51824 202650 51876
rect 202702 51824 202708 51876
rect 202920 51824 202926 51876
rect 202978 51824 202984 51876
rect 203380 51824 203386 51876
rect 203438 51824 203444 51876
rect 203564 51824 203570 51876
rect 203622 51824 203628 51876
rect 203656 51824 203662 51876
rect 203714 51824 203720 51876
rect 203748 51824 203754 51876
rect 203806 51824 203812 51876
rect 204024 51824 204030 51876
rect 204082 51824 204088 51876
rect 202202 51632 202236 51672
rect 201920 51620 201926 51632
rect 202230 51620 202236 51632
rect 202288 51620 202294 51672
rect 201034 51552 201040 51604
rect 201092 51552 201098 51604
rect 201604 51564 202230 51592
rect 200942 51524 200948 51536
rect 200730 51496 200948 51524
rect 199068 51484 199074 51496
rect 200942 51484 200948 51496
rect 201000 51484 201006 51536
rect 196710 51456 196716 51468
rect 196222 51428 196716 51456
rect 196710 51416 196716 51428
rect 196768 51416 196774 51468
rect 198550 51416 198556 51468
rect 198608 51416 198614 51468
rect 201604 51400 201632 51564
rect 202202 51456 202230 51564
rect 202662 51536 202690 51824
rect 202938 51660 202966 51824
rect 203398 51672 203426 51824
rect 203582 51672 203610 51824
rect 203058 51660 203064 51672
rect 202938 51632 203064 51660
rect 203058 51620 203064 51632
rect 203116 51620 203122 51672
rect 203398 51632 203432 51672
rect 203426 51620 203432 51632
rect 203484 51620 203490 51672
rect 203518 51620 203524 51672
rect 203576 51632 203610 51672
rect 203576 51620 203582 51632
rect 203674 51604 203702 51824
rect 203610 51552 203616 51604
rect 203668 51564 203702 51604
rect 203668 51552 203674 51564
rect 202598 51484 202604 51536
rect 202656 51496 202690 51536
rect 202656 51484 202662 51496
rect 203242 51484 203248 51536
rect 203300 51524 203306 51536
rect 203766 51524 203794 51824
rect 203886 51620 203892 51672
rect 203944 51660 203950 51672
rect 204042 51660 204070 51824
rect 204272 51672 204300 51904
rect 204392 51892 204398 51944
rect 204450 51892 204456 51944
rect 204576 51932 204582 51944
rect 204502 51904 204582 51932
rect 203944 51632 204070 51660
rect 203944 51620 203950 51632
rect 204254 51620 204260 51672
rect 204312 51620 204318 51672
rect 204070 51552 204076 51604
rect 204128 51592 204134 51604
rect 204410 51592 204438 51892
rect 204128 51564 204438 51592
rect 204128 51552 204134 51564
rect 204502 51536 204530 51904
rect 204576 51892 204582 51904
rect 204634 51892 204640 51944
rect 204668 51892 204674 51944
rect 204726 51892 204732 51944
rect 204760 51892 204766 51944
rect 204818 51892 204824 51944
rect 204852 51892 204858 51944
rect 204910 51892 204916 51944
rect 204944 51892 204950 51944
rect 205002 51892 205008 51944
rect 205036 51892 205042 51944
rect 205094 51892 205100 51944
rect 205312 51892 205318 51944
rect 205370 51892 205376 51944
rect 205496 51892 205502 51944
rect 205554 51892 205560 51944
rect 205588 51892 205594 51944
rect 205646 51892 205652 51944
rect 205680 51892 205686 51944
rect 205738 51892 205744 51944
rect 205772 51892 205778 51944
rect 205830 51892 205836 51944
rect 206232 51892 206238 51944
rect 206290 51892 206296 51944
rect 206600 51892 206606 51944
rect 206658 51892 206664 51944
rect 206692 51892 206698 51944
rect 206750 51892 206756 51944
rect 206802 51932 206830 52040
rect 208624 52028 208630 52080
rect 208682 52028 208688 52080
rect 208642 52000 208670 52028
rect 210850 52000 210878 52108
rect 216122 52096 216128 52108
rect 216180 52096 216186 52148
rect 222166 52068 222194 52176
rect 224926 52136 224954 52244
rect 258718 52136 258724 52148
rect 224926 52108 258724 52136
rect 258718 52096 258724 52108
rect 258776 52096 258782 52148
rect 212506 52040 219434 52068
rect 222166 52040 224954 52068
rect 212506 52000 212534 52040
rect 219406 52000 219434 52040
rect 208642 51972 209590 52000
rect 206802 51904 206922 51932
rect 204686 51864 204714 51892
rect 204640 51836 204714 51864
rect 204640 51740 204668 51836
rect 204778 51740 204806 51892
rect 204622 51688 204628 51740
rect 204680 51688 204686 51740
rect 204714 51688 204720 51740
rect 204772 51700 204806 51740
rect 204772 51688 204778 51700
rect 203300 51496 203794 51524
rect 203300 51484 203306 51496
rect 204438 51484 204444 51536
rect 204496 51496 204530 51536
rect 204870 51524 204898 51892
rect 204962 51808 204990 51892
rect 204944 51756 204950 51808
rect 205002 51756 205008 51808
rect 205054 51592 205082 51892
rect 205330 51808 205358 51892
rect 205514 51808 205542 51892
rect 205266 51756 205272 51808
rect 205324 51768 205358 51808
rect 205324 51756 205330 51768
rect 205450 51756 205456 51808
rect 205508 51768 205542 51808
rect 205508 51756 205514 51768
rect 205606 51740 205634 51892
rect 205698 51808 205726 51892
rect 205864 51824 205870 51876
rect 205922 51824 205928 51876
rect 205698 51768 205732 51808
rect 205726 51756 205732 51768
rect 205784 51756 205790 51808
rect 205606 51700 205640 51740
rect 205634 51688 205640 51700
rect 205692 51688 205698 51740
rect 205358 51620 205364 51672
rect 205416 51660 205422 51672
rect 205882 51660 205910 51824
rect 205956 51756 205962 51808
rect 206014 51756 206020 51808
rect 205416 51632 205910 51660
rect 205416 51620 205422 51632
rect 205974 51604 206002 51756
rect 206250 51604 206278 51892
rect 206416 51824 206422 51876
rect 206474 51824 206480 51876
rect 206434 51604 206462 51824
rect 206618 51808 206646 51892
rect 206600 51756 206606 51808
rect 206658 51756 206664 51808
rect 206710 51740 206738 51892
rect 206784 51824 206790 51876
rect 206842 51824 206848 51876
rect 206894 51864 206922 51904
rect 206968 51892 206974 51944
rect 207026 51932 207032 51944
rect 207152 51932 207158 51944
rect 207026 51892 207060 51932
rect 206894 51836 206968 51864
rect 206802 51796 206830 51824
rect 206940 51808 206968 51836
rect 206802 51768 206876 51796
rect 206710 51700 206744 51740
rect 206738 51688 206744 51700
rect 206796 51688 206802 51740
rect 205634 51592 205640 51604
rect 205054 51564 205640 51592
rect 205634 51552 205640 51564
rect 205692 51552 205698 51604
rect 205910 51552 205916 51604
rect 205968 51564 206002 51604
rect 205968 51552 205974 51564
rect 206186 51552 206192 51604
rect 206244 51564 206278 51604
rect 206244 51552 206250 51564
rect 206370 51552 206376 51604
rect 206428 51564 206462 51604
rect 206428 51552 206434 51564
rect 206278 51524 206284 51536
rect 204870 51496 206284 51524
rect 204496 51484 204502 51496
rect 206278 51484 206284 51496
rect 206336 51484 206342 51536
rect 206848 51524 206876 51768
rect 206922 51756 206928 51808
rect 206980 51756 206986 51808
rect 206922 51620 206928 51672
rect 206980 51660 206986 51672
rect 207032 51660 207060 51892
rect 206980 51632 207060 51660
rect 207124 51892 207158 51932
rect 207210 51892 207216 51944
rect 207888 51932 207894 51944
rect 207860 51892 207894 51932
rect 207946 51892 207952 51944
rect 208256 51892 208262 51944
rect 208314 51892 208320 51944
rect 208348 51892 208354 51944
rect 208406 51892 208412 51944
rect 208440 51892 208446 51944
rect 208498 51892 208504 51944
rect 209084 51892 209090 51944
rect 209142 51892 209148 51944
rect 209452 51932 209458 51944
rect 209424 51892 209458 51932
rect 209510 51892 209516 51944
rect 206980 51620 206986 51632
rect 207014 51552 207020 51604
rect 207072 51592 207078 51604
rect 207124 51592 207152 51892
rect 207428 51824 207434 51876
rect 207486 51864 207492 51876
rect 207486 51824 207520 51864
rect 207704 51824 207710 51876
rect 207762 51864 207768 51876
rect 207762 51824 207796 51864
rect 207244 51756 207250 51808
rect 207302 51756 207308 51808
rect 207262 51604 207290 51756
rect 207072 51564 207152 51592
rect 207072 51552 207078 51564
rect 207198 51552 207204 51604
rect 207256 51564 207290 51604
rect 207256 51552 207262 51564
rect 207492 51536 207520 51824
rect 207768 51672 207796 51824
rect 207750 51620 207756 51672
rect 207808 51620 207814 51672
rect 207658 51552 207664 51604
rect 207716 51592 207722 51604
rect 207860 51592 207888 51892
rect 208274 51796 208302 51892
rect 208228 51768 208302 51796
rect 208228 51740 208256 51768
rect 208366 51740 208394 51892
rect 208210 51688 208216 51740
rect 208268 51688 208274 51740
rect 208302 51688 208308 51740
rect 208360 51700 208394 51740
rect 208360 51688 208366 51700
rect 208458 51672 208486 51892
rect 208532 51824 208538 51876
rect 208590 51824 208596 51876
rect 208900 51824 208906 51876
rect 208958 51824 208964 51876
rect 208394 51620 208400 51672
rect 208452 51632 208486 51672
rect 208452 51620 208458 51632
rect 207716 51564 207888 51592
rect 207716 51552 207722 51564
rect 207382 51524 207388 51536
rect 206848 51496 207388 51524
rect 207382 51484 207388 51496
rect 207440 51484 207446 51536
rect 207474 51484 207480 51536
rect 207532 51484 207538 51536
rect 208550 51524 208578 51824
rect 208670 51688 208676 51740
rect 208728 51688 208734 51740
rect 208688 51604 208716 51688
rect 208918 51672 208946 51824
rect 209102 51672 209130 51892
rect 208918 51632 208952 51672
rect 208946 51620 208952 51632
rect 209004 51620 209010 51672
rect 209038 51620 209044 51672
rect 209096 51632 209130 51672
rect 209096 51620 209102 51632
rect 208670 51552 208676 51604
rect 208728 51552 208734 51604
rect 209424 51592 209452 51892
rect 209562 51672 209590 51972
rect 210574 51972 210878 52000
rect 211264 51972 212534 52000
rect 215450 51972 215984 52000
rect 219406 51972 222194 52000
rect 210004 51892 210010 51944
rect 210062 51892 210068 51944
rect 209912 51824 209918 51876
rect 209970 51824 209976 51876
rect 209498 51620 209504 51672
rect 209556 51632 209590 51672
rect 209556 51620 209562 51632
rect 209590 51592 209596 51604
rect 209424 51564 209596 51592
rect 209590 51552 209596 51564
rect 209648 51552 209654 51604
rect 209682 51524 209688 51536
rect 208550 51496 209688 51524
rect 209682 51484 209688 51496
rect 209740 51484 209746 51536
rect 209930 51524 209958 51824
rect 210022 51728 210050 51892
rect 210574 51808 210602 51972
rect 210648 51892 210654 51944
rect 210706 51932 210712 51944
rect 210706 51904 211016 51932
rect 210706 51892 210712 51904
rect 210832 51824 210838 51876
rect 210890 51824 210896 51876
rect 210574 51768 210608 51808
rect 210602 51756 210608 51768
rect 210660 51756 210666 51808
rect 210022 51700 210096 51728
rect 210068 51604 210096 51700
rect 210850 51672 210878 51824
rect 210786 51620 210792 51672
rect 210844 51632 210878 51672
rect 210844 51620 210850 51632
rect 210050 51552 210056 51604
rect 210108 51552 210114 51604
rect 210988 51536 211016 51904
rect 211264 51604 211292 51972
rect 215450 51944 215478 51972
rect 215956 51944 215984 51972
rect 211384 51892 211390 51944
rect 211442 51932 211448 51944
rect 211442 51904 211614 51932
rect 211442 51892 211448 51904
rect 211476 51756 211482 51808
rect 211534 51756 211540 51808
rect 211494 51728 211522 51756
rect 211448 51700 211522 51728
rect 211448 51604 211476 51700
rect 211246 51552 211252 51604
rect 211304 51552 211310 51604
rect 211430 51552 211436 51604
rect 211488 51552 211494 51604
rect 211586 51536 211614 51904
rect 212764 51892 212770 51944
rect 212822 51892 212828 51944
rect 212856 51892 212862 51944
rect 212914 51892 212920 51944
rect 212948 51892 212954 51944
rect 213006 51892 213012 51944
rect 213224 51892 213230 51944
rect 213282 51892 213288 51944
rect 213408 51892 213414 51944
rect 213466 51892 213472 51944
rect 213684 51892 213690 51944
rect 213742 51892 213748 51944
rect 213776 51892 213782 51944
rect 213834 51892 213840 51944
rect 213960 51932 213966 51944
rect 213932 51892 213966 51932
rect 214018 51892 214024 51944
rect 214880 51892 214886 51944
rect 214938 51892 214944 51944
rect 215064 51892 215070 51944
rect 215122 51892 215128 51944
rect 215156 51892 215162 51944
rect 215214 51892 215220 51944
rect 215248 51892 215254 51944
rect 215306 51932 215312 51944
rect 215306 51892 215340 51932
rect 215432 51892 215438 51944
rect 215490 51892 215496 51944
rect 215708 51892 215714 51944
rect 215766 51892 215772 51944
rect 215800 51892 215806 51944
rect 215858 51892 215864 51944
rect 215938 51892 215944 51944
rect 215996 51892 216002 51944
rect 211752 51824 211758 51876
rect 211810 51824 211816 51876
rect 212028 51824 212034 51876
rect 212086 51824 212092 51876
rect 212580 51824 212586 51876
rect 212638 51824 212644 51876
rect 212782 51864 212810 51892
rect 212736 51836 212810 51864
rect 211770 51672 211798 51824
rect 211706 51620 211712 51672
rect 211764 51632 211798 51672
rect 211764 51620 211770 51632
rect 212046 51592 212074 51824
rect 212598 51740 212626 51824
rect 212534 51688 212540 51740
rect 212592 51700 212626 51740
rect 212592 51688 212598 51700
rect 212736 51604 212764 51836
rect 212874 51808 212902 51892
rect 212810 51756 212816 51808
rect 212868 51768 212902 51808
rect 212868 51756 212874 51768
rect 212966 51740 212994 51892
rect 213040 51824 213046 51876
rect 213098 51824 213104 51876
rect 212902 51688 212908 51740
rect 212960 51700 212994 51740
rect 212960 51688 212966 51700
rect 213058 51604 213086 51824
rect 213242 51740 213270 51892
rect 213242 51700 213276 51740
rect 213270 51688 213276 51700
rect 213328 51688 213334 51740
rect 213426 51660 213454 51892
rect 213500 51824 213506 51876
rect 213558 51824 213564 51876
rect 212166 51592 212172 51604
rect 212046 51564 212172 51592
rect 212166 51552 212172 51564
rect 212224 51552 212230 51604
rect 212718 51552 212724 51604
rect 212776 51552 212782 51604
rect 212994 51552 213000 51604
rect 213052 51564 213086 51604
rect 213150 51632 213454 51660
rect 213052 51552 213058 51564
rect 210326 51524 210332 51536
rect 209930 51496 210332 51524
rect 210326 51484 210332 51496
rect 210384 51484 210390 51536
rect 210970 51484 210976 51536
rect 211028 51484 211034 51536
rect 211586 51496 211620 51536
rect 211614 51484 211620 51496
rect 211672 51484 211678 51536
rect 212442 51484 212448 51536
rect 212500 51524 212506 51536
rect 213150 51524 213178 51632
rect 213518 51604 213546 51824
rect 213702 51808 213730 51892
rect 213684 51756 213690 51808
rect 213742 51756 213748 51808
rect 213518 51564 213552 51604
rect 213546 51552 213552 51564
rect 213604 51552 213610 51604
rect 213638 51552 213644 51604
rect 213696 51592 213702 51604
rect 213794 51592 213822 51892
rect 213932 51740 213960 51892
rect 214052 51864 214058 51876
rect 214024 51824 214058 51864
rect 214110 51824 214116 51876
rect 214144 51824 214150 51876
rect 214202 51824 214208 51876
rect 214024 51740 214052 51824
rect 213914 51688 213920 51740
rect 213972 51688 213978 51740
rect 214006 51688 214012 51740
rect 214064 51688 214070 51740
rect 214162 51672 214190 51824
rect 214898 51740 214926 51892
rect 215082 51808 215110 51892
rect 215174 51864 215202 51892
rect 215174 51836 215248 51864
rect 215220 51808 215248 51836
rect 215082 51768 215116 51808
rect 215110 51756 215116 51768
rect 215168 51756 215174 51808
rect 215202 51756 215208 51808
rect 215260 51756 215266 51808
rect 214834 51688 214840 51740
rect 214892 51700 214926 51740
rect 214892 51688 214898 51700
rect 214098 51620 214104 51672
rect 214156 51632 214190 51672
rect 214156 51620 214162 51632
rect 213696 51564 213822 51592
rect 214484 51564 214880 51592
rect 213696 51552 213702 51564
rect 214484 51524 214512 51564
rect 212500 51496 213178 51524
rect 213242 51496 214512 51524
rect 214852 51524 214880 51564
rect 214926 51552 214932 51604
rect 214984 51592 214990 51604
rect 215312 51592 215340 51892
rect 215726 51808 215754 51892
rect 215818 51864 215846 51892
rect 215818 51836 215892 51864
rect 215864 51808 215892 51836
rect 215726 51768 215760 51808
rect 215754 51756 215760 51768
rect 215812 51756 215818 51808
rect 215846 51756 215852 51808
rect 215904 51756 215910 51808
rect 222166 51796 222194 51972
rect 224926 51864 224954 52040
rect 234706 51864 234712 51876
rect 224926 51836 234712 51864
rect 234706 51824 234712 51836
rect 234764 51824 234770 51876
rect 253566 51796 253572 51808
rect 222166 51768 253572 51796
rect 253566 51756 253572 51768
rect 253624 51756 253630 51808
rect 216582 51688 216588 51740
rect 216640 51728 216646 51740
rect 238754 51728 238760 51740
rect 216640 51700 238760 51728
rect 216640 51688 216646 51700
rect 238754 51688 238760 51700
rect 238812 51688 238818 51740
rect 216122 51620 216128 51672
rect 216180 51660 216186 51672
rect 253474 51660 253480 51672
rect 216180 51632 253480 51660
rect 216180 51620 216186 51632
rect 253474 51620 253480 51632
rect 253532 51620 253538 51672
rect 214984 51564 215340 51592
rect 214984 51552 214990 51564
rect 216398 51552 216404 51604
rect 216456 51592 216462 51604
rect 258810 51592 258816 51604
rect 216456 51564 258816 51592
rect 216456 51552 216462 51564
rect 258810 51552 258816 51564
rect 258868 51552 258874 51604
rect 242894 51524 242900 51536
rect 214852 51496 242900 51524
rect 212500 51484 212506 51496
rect 213242 51456 213270 51496
rect 242894 51484 242900 51496
rect 242952 51484 242958 51536
rect 202202 51428 213270 51456
rect 216214 51416 216220 51468
rect 216272 51456 216278 51468
rect 256326 51456 256332 51468
rect 216272 51428 256332 51456
rect 216272 51416 216278 51428
rect 256326 51416 256332 51428
rect 256384 51416 256390 51468
rect 194502 51388 194508 51400
rect 193968 51360 194508 51388
rect 194502 51348 194508 51360
rect 194560 51348 194566 51400
rect 194778 51348 194784 51400
rect 194836 51388 194842 51400
rect 194836 51360 200114 51388
rect 194836 51348 194842 51360
rect 188488 51292 188706 51320
rect 200086 51320 200114 51360
rect 201586 51348 201592 51400
rect 201644 51348 201650 51400
rect 202046 51348 202052 51400
rect 202104 51388 202110 51400
rect 256234 51388 256240 51400
rect 202104 51360 256240 51388
rect 202104 51348 202110 51360
rect 256234 51348 256240 51360
rect 256292 51348 256298 51400
rect 256142 51320 256148 51332
rect 200086 51292 256148 51320
rect 188488 51280 188494 51292
rect 256142 51280 256148 51292
rect 256200 51280 256206 51332
rect 238018 51252 238024 51264
rect 175148 51224 181024 51252
rect 183526 51224 183738 51252
rect 188356 51224 238024 51252
rect 175148 51212 175154 51224
rect 159450 51144 159456 51196
rect 159508 51184 159514 51196
rect 176378 51184 176384 51196
rect 159508 51156 176384 51184
rect 159508 51144 159514 51156
rect 176378 51144 176384 51156
rect 176436 51144 176442 51196
rect 178770 51144 178776 51196
rect 178828 51184 178834 51196
rect 179138 51184 179144 51196
rect 178828 51156 179144 51184
rect 178828 51144 178834 51156
rect 179138 51144 179144 51156
rect 179196 51144 179202 51196
rect 183526 51184 183554 51224
rect 179294 51156 183554 51184
rect 183710 51184 183738 51224
rect 238018 51212 238024 51224
rect 238076 51212 238082 51264
rect 253198 51184 253204 51196
rect 183710 51156 253204 51184
rect 171870 51116 171876 51128
rect 160250 51088 171876 51116
rect 160250 51060 160278 51088
rect 171870 51076 171876 51088
rect 171928 51076 171934 51128
rect 174998 51076 175004 51128
rect 175056 51116 175062 51128
rect 179294 51116 179322 51156
rect 253198 51144 253204 51156
rect 253256 51144 253262 51196
rect 175056 51088 179322 51116
rect 175056 51076 175062 51088
rect 180242 51076 180248 51128
rect 180300 51116 180306 51128
rect 180794 51116 180800 51128
rect 180300 51088 180800 51116
rect 180300 51076 180306 51088
rect 180794 51076 180800 51088
rect 180852 51076 180858 51128
rect 188890 51076 188896 51128
rect 188948 51116 188954 51128
rect 220814 51116 220820 51128
rect 188948 51088 220820 51116
rect 188948 51076 188954 51088
rect 220814 51076 220820 51088
rect 220872 51076 220878 51128
rect 160186 51008 160192 51060
rect 160244 51020 160278 51060
rect 160244 51008 160250 51020
rect 162854 51008 162860 51060
rect 162912 51048 162918 51060
rect 173434 51048 173440 51060
rect 162912 51020 173440 51048
rect 162912 51008 162918 51020
rect 173434 51008 173440 51020
rect 173492 51008 173498 51060
rect 174906 51008 174912 51060
rect 174964 51048 174970 51060
rect 246482 51048 246488 51060
rect 174964 51020 246488 51048
rect 174964 51008 174970 51020
rect 246482 51008 246488 51020
rect 246540 51008 246546 51060
rect 255958 51008 255964 51060
rect 256016 51048 256022 51060
rect 256694 51048 256700 51060
rect 256016 51020 256700 51048
rect 256016 51008 256022 51020
rect 256694 51008 256700 51020
rect 256752 51008 256758 51060
rect 173710 50980 173716 50992
rect 158686 50952 173716 50980
rect 173710 50940 173716 50952
rect 173768 50940 173774 50992
rect 175274 50940 175280 50992
rect 175332 50980 175338 50992
rect 246390 50980 246396 50992
rect 175332 50952 246396 50980
rect 175332 50940 175338 50952
rect 246390 50940 246396 50952
rect 246448 50940 246454 50992
rect 170950 50912 170956 50924
rect 168346 50884 170956 50912
rect 156690 50804 156696 50856
rect 156748 50844 156754 50856
rect 159818 50844 159824 50856
rect 156748 50816 159824 50844
rect 156748 50804 156754 50816
rect 159818 50804 159824 50816
rect 159876 50804 159882 50856
rect 159266 50736 159272 50788
rect 159324 50776 159330 50788
rect 168346 50776 168374 50884
rect 170950 50872 170956 50884
rect 171008 50872 171014 50924
rect 172238 50872 172244 50924
rect 172296 50912 172302 50924
rect 231118 50912 231124 50924
rect 172296 50884 231124 50912
rect 172296 50872 172302 50884
rect 231118 50872 231124 50884
rect 231176 50872 231182 50924
rect 171778 50804 171784 50856
rect 171836 50844 171842 50856
rect 220170 50844 220176 50856
rect 171836 50816 220176 50844
rect 171836 50804 171842 50816
rect 220170 50804 220176 50816
rect 220228 50804 220234 50856
rect 159324 50748 168374 50776
rect 159324 50736 159330 50748
rect 175550 50736 175556 50788
rect 175608 50776 175614 50788
rect 175608 50748 176654 50776
rect 175608 50736 175614 50748
rect 148318 50668 148324 50720
rect 148376 50708 148382 50720
rect 175918 50708 175924 50720
rect 148376 50680 175924 50708
rect 148376 50668 148382 50680
rect 175918 50668 175924 50680
rect 175976 50668 175982 50720
rect 176626 50708 176654 50748
rect 179230 50736 179236 50788
rect 179288 50776 179294 50788
rect 220078 50776 220084 50788
rect 179288 50748 220084 50776
rect 179288 50736 179294 50748
rect 220078 50736 220084 50748
rect 220136 50736 220142 50788
rect 218054 50708 218060 50720
rect 176626 50680 218060 50708
rect 218054 50668 218060 50680
rect 218112 50668 218118 50720
rect 151354 50600 151360 50652
rect 151412 50640 151418 50652
rect 179046 50640 179052 50652
rect 151412 50612 179052 50640
rect 151412 50600 151418 50612
rect 179046 50600 179052 50612
rect 179104 50600 179110 50652
rect 179782 50600 179788 50652
rect 179840 50640 179846 50652
rect 180518 50640 180524 50652
rect 179840 50612 180524 50640
rect 179840 50600 179846 50612
rect 180518 50600 180524 50612
rect 180576 50600 180582 50652
rect 188706 50600 188712 50652
rect 188764 50600 188770 50652
rect 188890 50600 188896 50652
rect 188948 50640 188954 50652
rect 189166 50640 189172 50652
rect 188948 50612 189172 50640
rect 188948 50600 188954 50612
rect 189166 50600 189172 50612
rect 189224 50600 189230 50652
rect 190362 50600 190368 50652
rect 190420 50640 190426 50652
rect 201586 50640 201592 50652
rect 190420 50612 201592 50640
rect 190420 50600 190426 50612
rect 201586 50600 201592 50612
rect 201644 50600 201650 50652
rect 204622 50600 204628 50652
rect 204680 50640 204686 50652
rect 253198 50640 253204 50652
rect 204680 50612 253204 50640
rect 204680 50600 204686 50612
rect 253198 50600 253204 50612
rect 253256 50600 253262 50652
rect 159818 50532 159824 50584
rect 159876 50572 159882 50584
rect 178034 50572 178040 50584
rect 159876 50544 178040 50572
rect 159876 50532 159882 50544
rect 178034 50532 178040 50544
rect 178092 50532 178098 50584
rect 178402 50532 178408 50584
rect 178460 50572 178466 50584
rect 179506 50572 179512 50584
rect 178460 50544 179512 50572
rect 178460 50532 178466 50544
rect 179506 50532 179512 50544
rect 179564 50532 179570 50584
rect 134518 50464 134524 50516
rect 134576 50504 134582 50516
rect 177942 50504 177948 50516
rect 134576 50476 177948 50504
rect 134576 50464 134582 50476
rect 177942 50464 177948 50476
rect 178000 50464 178006 50516
rect 188724 50448 188752 50600
rect 196434 50532 196440 50584
rect 196492 50572 196498 50584
rect 202046 50572 202052 50584
rect 196492 50544 202052 50572
rect 196492 50532 196498 50544
rect 202046 50532 202052 50544
rect 202104 50532 202110 50584
rect 205634 50532 205640 50584
rect 205692 50572 205698 50584
rect 206094 50572 206100 50584
rect 205692 50544 206100 50572
rect 205692 50532 205698 50544
rect 206094 50532 206100 50544
rect 206152 50532 206158 50584
rect 206278 50532 206284 50584
rect 206336 50572 206342 50584
rect 208026 50572 208032 50584
rect 206336 50544 208032 50572
rect 206336 50532 206342 50544
rect 208026 50532 208032 50544
rect 208084 50532 208090 50584
rect 212506 50544 214834 50572
rect 200482 50464 200488 50516
rect 200540 50504 200546 50516
rect 212506 50504 212534 50544
rect 200540 50476 212534 50504
rect 214806 50504 214834 50544
rect 214926 50532 214932 50584
rect 214984 50572 214990 50584
rect 258718 50572 258724 50584
rect 214984 50544 258724 50572
rect 214984 50532 214990 50544
rect 258718 50532 258724 50544
rect 258776 50532 258782 50584
rect 253290 50504 253296 50516
rect 214806 50476 253296 50504
rect 200540 50464 200546 50476
rect 253290 50464 253296 50476
rect 253348 50464 253354 50516
rect 154022 50396 154028 50448
rect 154080 50436 154086 50448
rect 177758 50436 177764 50448
rect 154080 50408 177764 50436
rect 154080 50396 154086 50408
rect 177758 50396 177764 50408
rect 177816 50396 177822 50448
rect 179506 50396 179512 50448
rect 179564 50436 179570 50448
rect 179874 50436 179880 50448
rect 179564 50408 179880 50436
rect 179564 50396 179570 50408
rect 179874 50396 179880 50408
rect 179932 50396 179938 50448
rect 183830 50396 183836 50448
rect 183888 50436 183894 50448
rect 184934 50436 184940 50448
rect 183888 50408 184940 50436
rect 183888 50396 183894 50408
rect 184934 50396 184940 50408
rect 184992 50396 184998 50448
rect 188706 50396 188712 50448
rect 188764 50396 188770 50448
rect 197538 50396 197544 50448
rect 197596 50436 197602 50448
rect 197596 50408 212534 50436
rect 197596 50396 197602 50408
rect 160370 50328 160376 50380
rect 160428 50368 160434 50380
rect 160554 50368 160560 50380
rect 160428 50340 160560 50368
rect 160428 50328 160434 50340
rect 160554 50328 160560 50340
rect 160612 50328 160618 50380
rect 172330 50328 172336 50380
rect 172388 50368 172394 50380
rect 179230 50368 179236 50380
rect 172388 50340 179236 50368
rect 172388 50328 172394 50340
rect 179230 50328 179236 50340
rect 179288 50328 179294 50380
rect 190638 50328 190644 50380
rect 190696 50368 190702 50380
rect 207106 50368 207112 50380
rect 190696 50340 207112 50368
rect 190696 50328 190702 50340
rect 207106 50328 207112 50340
rect 207164 50328 207170 50380
rect 207290 50328 207296 50380
rect 207348 50368 207354 50380
rect 207474 50368 207480 50380
rect 207348 50340 207480 50368
rect 207348 50328 207354 50340
rect 207474 50328 207480 50340
rect 207532 50328 207538 50380
rect 210602 50368 210608 50380
rect 210252 50340 210608 50368
rect 144178 50260 144184 50312
rect 144236 50300 144242 50312
rect 176562 50300 176568 50312
rect 144236 50272 176568 50300
rect 144236 50260 144242 50272
rect 176562 50260 176568 50272
rect 176620 50260 176626 50312
rect 188338 50260 188344 50312
rect 188396 50300 188402 50312
rect 188396 50272 195974 50300
rect 188396 50260 188402 50272
rect 141418 50192 141424 50244
rect 141476 50232 141482 50244
rect 176010 50232 176016 50244
rect 141476 50204 176016 50232
rect 141476 50192 141482 50204
rect 176010 50192 176016 50204
rect 176068 50192 176074 50244
rect 188062 50192 188068 50244
rect 188120 50232 188126 50244
rect 188798 50232 188804 50244
rect 188120 50204 188804 50232
rect 188120 50192 188126 50204
rect 188798 50192 188804 50204
rect 188856 50192 188862 50244
rect 159450 50124 159456 50176
rect 159508 50164 159514 50176
rect 161842 50164 161848 50176
rect 159508 50136 161848 50164
rect 159508 50124 159514 50136
rect 161842 50124 161848 50136
rect 161900 50124 161906 50176
rect 171226 50124 171232 50176
rect 171284 50164 171290 50176
rect 171870 50164 171876 50176
rect 171284 50136 171876 50164
rect 171284 50124 171290 50136
rect 171870 50124 171876 50136
rect 171928 50124 171934 50176
rect 174262 50124 174268 50176
rect 174320 50164 174326 50176
rect 178862 50164 178868 50176
rect 174320 50136 178868 50164
rect 174320 50124 174326 50136
rect 178862 50124 178868 50136
rect 178920 50124 178926 50176
rect 184934 50124 184940 50176
rect 184992 50164 184998 50176
rect 185578 50164 185584 50176
rect 184992 50136 185584 50164
rect 184992 50124 184998 50136
rect 185578 50124 185584 50136
rect 185636 50124 185642 50176
rect 190178 50124 190184 50176
rect 190236 50164 190242 50176
rect 190362 50164 190368 50176
rect 190236 50136 190368 50164
rect 190236 50124 190242 50136
rect 190362 50124 190368 50136
rect 190420 50124 190426 50176
rect 193398 50124 193404 50176
rect 193456 50164 193462 50176
rect 193950 50164 193956 50176
rect 193456 50136 193956 50164
rect 193456 50124 193462 50136
rect 193950 50124 193956 50136
rect 194008 50124 194014 50176
rect 138658 50056 138664 50108
rect 138716 50096 138722 50108
rect 176286 50096 176292 50108
rect 138716 50068 176292 50096
rect 138716 50056 138722 50068
rect 176286 50056 176292 50068
rect 176344 50056 176350 50108
rect 195946 50096 195974 50272
rect 204254 50260 204260 50312
rect 204312 50300 204318 50312
rect 210252 50300 210280 50340
rect 210602 50328 210608 50340
rect 210660 50328 210666 50380
rect 210694 50328 210700 50380
rect 210752 50368 210758 50380
rect 210878 50368 210884 50380
rect 210752 50340 210884 50368
rect 210752 50328 210758 50340
rect 210878 50328 210884 50340
rect 210936 50328 210942 50380
rect 211798 50328 211804 50380
rect 211856 50368 211862 50380
rect 211982 50368 211988 50380
rect 211856 50340 211988 50368
rect 211856 50328 211862 50340
rect 211982 50328 211988 50340
rect 212040 50328 212046 50380
rect 212506 50368 212534 50408
rect 213454 50396 213460 50448
rect 213512 50436 213518 50448
rect 214190 50436 214196 50448
rect 213512 50408 214196 50436
rect 213512 50396 213518 50408
rect 214190 50396 214196 50408
rect 214248 50396 214254 50448
rect 256602 50436 256608 50448
rect 214806 50408 256608 50436
rect 214806 50368 214834 50408
rect 256602 50396 256608 50408
rect 256660 50396 256666 50448
rect 252554 50368 252560 50380
rect 212506 50340 214834 50368
rect 215266 50340 252560 50368
rect 204312 50272 210280 50300
rect 204312 50260 204318 50272
rect 210326 50260 210332 50312
rect 210384 50300 210390 50312
rect 214926 50300 214932 50312
rect 210384 50272 214932 50300
rect 210384 50260 210390 50272
rect 214926 50260 214932 50272
rect 214984 50260 214990 50312
rect 204990 50192 204996 50244
rect 205048 50232 205054 50244
rect 206186 50232 206192 50244
rect 205048 50204 206192 50232
rect 205048 50192 205054 50204
rect 206186 50192 206192 50204
rect 206244 50192 206250 50244
rect 207474 50192 207480 50244
rect 207532 50232 207538 50244
rect 207842 50232 207848 50244
rect 207532 50204 207848 50232
rect 207532 50192 207538 50204
rect 207842 50192 207848 50204
rect 207900 50192 207906 50244
rect 208026 50192 208032 50244
rect 208084 50232 208090 50244
rect 208302 50232 208308 50244
rect 208084 50204 208308 50232
rect 208084 50192 208090 50204
rect 208302 50192 208308 50204
rect 208360 50192 208366 50244
rect 208486 50192 208492 50244
rect 208544 50232 208550 50244
rect 209406 50232 209412 50244
rect 208544 50204 209412 50232
rect 208544 50192 208550 50204
rect 209406 50192 209412 50204
rect 209464 50192 209470 50244
rect 211982 50192 211988 50244
rect 212040 50232 212046 50244
rect 215266 50232 215294 50340
rect 252554 50328 252560 50340
rect 252612 50328 252618 50380
rect 580074 50328 580080 50380
rect 580132 50368 580138 50380
rect 580810 50368 580816 50380
rect 580132 50340 580816 50368
rect 580132 50328 580138 50340
rect 580810 50328 580816 50340
rect 580868 50328 580874 50380
rect 212040 50204 215294 50232
rect 212040 50192 212046 50204
rect 204806 50124 204812 50176
rect 204864 50164 204870 50176
rect 205082 50164 205088 50176
rect 204864 50136 205088 50164
rect 204864 50124 204870 50136
rect 205082 50124 205088 50136
rect 205140 50124 205146 50176
rect 205174 50124 205180 50176
rect 205232 50164 205238 50176
rect 205634 50164 205640 50176
rect 205232 50136 205640 50164
rect 205232 50124 205238 50136
rect 205634 50124 205640 50136
rect 205692 50124 205698 50176
rect 206094 50124 206100 50176
rect 206152 50164 206158 50176
rect 206370 50164 206376 50176
rect 206152 50136 206376 50164
rect 206152 50124 206158 50136
rect 206370 50124 206376 50136
rect 206428 50124 206434 50176
rect 208394 50124 208400 50176
rect 208452 50164 208458 50176
rect 208578 50164 208584 50176
rect 208452 50136 208584 50164
rect 208452 50124 208458 50136
rect 208578 50124 208584 50136
rect 208636 50124 208642 50176
rect 211126 50136 213546 50164
rect 211126 50096 211154 50136
rect 195946 50068 211154 50096
rect 213518 50096 213546 50136
rect 223574 50096 223580 50108
rect 213518 50068 223580 50096
rect 223574 50056 223580 50068
rect 223632 50056 223638 50108
rect 158070 49988 158076 50040
rect 158128 50028 158134 50040
rect 161474 50028 161480 50040
rect 158128 50000 161480 50028
rect 158128 49988 158134 50000
rect 161474 49988 161480 50000
rect 161532 49988 161538 50040
rect 175642 49988 175648 50040
rect 175700 50028 175706 50040
rect 178126 50028 178132 50040
rect 175700 50000 178132 50028
rect 175700 49988 175706 50000
rect 178126 49988 178132 50000
rect 178184 49988 178190 50040
rect 205358 49988 205364 50040
rect 205416 50028 205422 50040
rect 205910 50028 205916 50040
rect 205416 50000 205916 50028
rect 205416 49988 205422 50000
rect 205910 49988 205916 50000
rect 205968 49988 205974 50040
rect 207198 49988 207204 50040
rect 207256 50028 207262 50040
rect 207382 50028 207388 50040
rect 207256 50000 207388 50028
rect 207256 49988 207262 50000
rect 207382 49988 207388 50000
rect 207440 49988 207446 50040
rect 208394 49988 208400 50040
rect 208452 50028 208458 50040
rect 209130 50028 209136 50040
rect 208452 50000 209136 50028
rect 208452 49988 208458 50000
rect 209130 49988 209136 50000
rect 209188 49988 209194 50040
rect 212718 49988 212724 50040
rect 212776 50028 212782 50040
rect 213086 50028 213092 50040
rect 212776 50000 213092 50028
rect 212776 49988 212782 50000
rect 213086 49988 213092 50000
rect 213144 49988 213150 50040
rect 158530 49920 158536 49972
rect 158588 49960 158594 49972
rect 168466 49960 168472 49972
rect 158588 49932 168472 49960
rect 158588 49920 158594 49932
rect 168466 49920 168472 49932
rect 168524 49920 168530 49972
rect 207106 49920 207112 49972
rect 207164 49960 207170 49972
rect 211982 49960 211988 49972
rect 207164 49932 211988 49960
rect 207164 49920 207170 49932
rect 211982 49920 211988 49932
rect 212040 49920 212046 49972
rect 216582 49960 216588 49972
rect 212506 49932 216588 49960
rect 158162 49852 158168 49904
rect 158220 49892 158226 49904
rect 176746 49892 176752 49904
rect 158220 49864 176752 49892
rect 158220 49852 158226 49864
rect 176746 49852 176752 49864
rect 176804 49852 176810 49904
rect 181990 49852 181996 49904
rect 182048 49892 182054 49904
rect 182174 49892 182180 49904
rect 182048 49864 182180 49892
rect 182048 49852 182054 49864
rect 182174 49852 182180 49864
rect 182232 49852 182238 49904
rect 204070 49852 204076 49904
rect 204128 49892 204134 49904
rect 211246 49892 211252 49904
rect 204128 49864 211252 49892
rect 204128 49852 204134 49864
rect 211246 49852 211252 49864
rect 211304 49852 211310 49904
rect 181806 49784 181812 49836
rect 181864 49824 181870 49836
rect 184658 49824 184664 49836
rect 181864 49796 184664 49824
rect 181864 49784 181870 49796
rect 184658 49784 184664 49796
rect 184716 49784 184722 49836
rect 201034 49784 201040 49836
rect 201092 49824 201098 49836
rect 212506 49824 212534 49932
rect 216582 49920 216588 49932
rect 216640 49920 216646 49972
rect 212902 49852 212908 49904
rect 212960 49892 212966 49904
rect 213362 49892 213368 49904
rect 212960 49864 213368 49892
rect 212960 49852 212966 49864
rect 213362 49852 213368 49864
rect 213420 49852 213426 49904
rect 201092 49796 212534 49824
rect 201092 49784 201098 49796
rect 212626 49784 212632 49836
rect 212684 49824 212690 49836
rect 220170 49824 220176 49836
rect 212684 49796 220176 49824
rect 212684 49784 212690 49796
rect 220170 49784 220176 49796
rect 220228 49784 220234 49836
rect 182174 49716 182180 49768
rect 182232 49756 182238 49768
rect 184014 49756 184020 49768
rect 182232 49728 184020 49756
rect 182232 49716 182238 49728
rect 184014 49716 184020 49728
rect 184072 49716 184078 49768
rect 204438 49716 204444 49768
rect 204496 49756 204502 49768
rect 207842 49756 207848 49768
rect 204496 49728 207848 49756
rect 204496 49716 204502 49728
rect 207842 49716 207848 49728
rect 207900 49716 207906 49768
rect 212534 49716 212540 49768
rect 212592 49756 212598 49768
rect 212718 49756 212724 49768
rect 212592 49728 212724 49756
rect 212592 49716 212598 49728
rect 212718 49716 212724 49728
rect 212776 49716 212782 49768
rect 212902 49716 212908 49768
rect 212960 49756 212966 49768
rect 256050 49756 256056 49768
rect 212960 49728 256056 49756
rect 212960 49716 212966 49728
rect 256050 49716 256056 49728
rect 256108 49716 256114 49768
rect 158622 49648 158628 49700
rect 158680 49688 158686 49700
rect 161934 49688 161940 49700
rect 158680 49660 161940 49688
rect 158680 49648 158686 49660
rect 161934 49648 161940 49660
rect 161992 49648 161998 49700
rect 187694 49648 187700 49700
rect 187752 49688 187758 49700
rect 188062 49688 188068 49700
rect 187752 49660 188068 49688
rect 187752 49648 187758 49660
rect 188062 49648 188068 49660
rect 188120 49648 188126 49700
rect 203886 49648 203892 49700
rect 203944 49688 203950 49700
rect 208026 49688 208032 49700
rect 203944 49660 208032 49688
rect 203944 49648 203950 49660
rect 208026 49648 208032 49660
rect 208084 49648 208090 49700
rect 158162 49580 158168 49632
rect 158220 49620 158226 49632
rect 159450 49620 159456 49632
rect 158220 49592 159456 49620
rect 158220 49580 158226 49592
rect 159450 49580 159456 49592
rect 159508 49580 159514 49632
rect 160830 49580 160836 49632
rect 160888 49620 160894 49632
rect 161014 49620 161020 49632
rect 160888 49592 161020 49620
rect 160888 49580 160894 49592
rect 161014 49580 161020 49592
rect 161072 49580 161078 49632
rect 175366 49580 175372 49632
rect 175424 49620 175430 49632
rect 234614 49620 234620 49632
rect 175424 49592 234620 49620
rect 175424 49580 175430 49592
rect 234614 49580 234620 49592
rect 234672 49580 234678 49632
rect 160186 49512 160192 49564
rect 160244 49552 160250 49564
rect 161106 49552 161112 49564
rect 160244 49524 161112 49552
rect 160244 49512 160250 49524
rect 161106 49512 161112 49524
rect 161164 49512 161170 49564
rect 173158 49512 173164 49564
rect 173216 49552 173222 49564
rect 177022 49552 177028 49564
rect 173216 49524 177028 49552
rect 173216 49512 173222 49524
rect 177022 49512 177028 49524
rect 177080 49512 177086 49564
rect 228358 49552 228364 49564
rect 186286 49524 228364 49552
rect 157794 49444 157800 49496
rect 157852 49484 157858 49496
rect 166994 49484 167000 49496
rect 157852 49456 167000 49484
rect 157852 49444 157858 49456
rect 166994 49444 167000 49456
rect 167052 49444 167058 49496
rect 172146 49444 172152 49496
rect 172204 49484 172210 49496
rect 186286 49484 186314 49524
rect 228358 49512 228364 49524
rect 228416 49512 228422 49564
rect 172204 49456 186314 49484
rect 172204 49444 172210 49456
rect 209682 49444 209688 49496
rect 209740 49484 209746 49496
rect 209740 49456 220124 49484
rect 209740 49444 209746 49456
rect 157978 49376 157984 49428
rect 158036 49416 158042 49428
rect 160094 49416 160100 49428
rect 158036 49388 160100 49416
rect 158036 49376 158042 49388
rect 160094 49376 160100 49388
rect 160152 49376 160158 49428
rect 178494 49416 178500 49428
rect 170876 49388 178500 49416
rect 160554 49308 160560 49360
rect 160612 49348 160618 49360
rect 161382 49348 161388 49360
rect 160612 49320 161388 49348
rect 160612 49308 160618 49320
rect 161382 49308 161388 49320
rect 161440 49308 161446 49360
rect 170876 49280 170904 49388
rect 178494 49376 178500 49388
rect 178552 49376 178558 49428
rect 186774 49376 186780 49428
rect 186832 49416 186838 49428
rect 187694 49416 187700 49428
rect 186832 49388 187700 49416
rect 186832 49376 186838 49388
rect 187694 49376 187700 49388
rect 187752 49376 187758 49428
rect 193674 49376 193680 49428
rect 193732 49416 193738 49428
rect 212902 49416 212908 49428
rect 193732 49388 212908 49416
rect 193732 49376 193738 49388
rect 212902 49376 212908 49388
rect 212960 49376 212966 49428
rect 213196 49388 215294 49416
rect 172514 49308 172520 49360
rect 172572 49348 172578 49360
rect 176930 49348 176936 49360
rect 172572 49320 176936 49348
rect 172572 49308 172578 49320
rect 176930 49308 176936 49320
rect 176988 49308 176994 49360
rect 211982 49308 211988 49360
rect 212040 49348 212046 49360
rect 213196 49348 213224 49388
rect 212040 49320 213224 49348
rect 215266 49348 215294 49388
rect 218238 49348 218244 49360
rect 215266 49320 218244 49348
rect 212040 49308 212046 49320
rect 218238 49308 218244 49320
rect 218296 49308 218302 49360
rect 220096 49348 220124 49456
rect 220170 49444 220176 49496
rect 220228 49484 220234 49496
rect 220228 49456 224954 49484
rect 220228 49444 220234 49456
rect 224926 49416 224954 49456
rect 260098 49416 260104 49428
rect 224926 49388 260104 49416
rect 260098 49376 260104 49388
rect 260156 49376 260162 49428
rect 258994 49348 259000 49360
rect 220096 49320 259000 49348
rect 258994 49308 259000 49320
rect 259052 49308 259058 49360
rect 166966 49252 170904 49280
rect 158346 49172 158352 49224
rect 158404 49212 158410 49224
rect 166966 49212 166994 49252
rect 172698 49240 172704 49292
rect 172756 49280 172762 49292
rect 177942 49280 177948 49292
rect 172756 49252 177948 49280
rect 172756 49240 172762 49252
rect 177942 49240 177948 49252
rect 178000 49240 178006 49292
rect 186774 49240 186780 49292
rect 186832 49280 186838 49292
rect 186958 49280 186964 49292
rect 186832 49252 186964 49280
rect 186832 49240 186838 49252
rect 186958 49240 186964 49252
rect 187016 49240 187022 49292
rect 203702 49240 203708 49292
rect 203760 49280 203766 49292
rect 206646 49280 206652 49292
rect 203760 49252 206652 49280
rect 203760 49240 203766 49252
rect 206646 49240 206652 49252
rect 206704 49240 206710 49292
rect 208302 49240 208308 49292
rect 208360 49280 208366 49292
rect 258626 49280 258632 49292
rect 208360 49252 258632 49280
rect 208360 49240 208366 49252
rect 258626 49240 258632 49252
rect 258684 49240 258690 49292
rect 158404 49184 166994 49212
rect 158404 49172 158410 49184
rect 167454 49172 167460 49224
rect 167512 49212 167518 49224
rect 168466 49212 168472 49224
rect 167512 49184 168472 49212
rect 167512 49172 167518 49184
rect 168466 49172 168472 49184
rect 168524 49172 168530 49224
rect 171962 49172 171968 49224
rect 172020 49212 172026 49224
rect 173802 49212 173808 49224
rect 172020 49184 173808 49212
rect 172020 49172 172026 49184
rect 173802 49172 173808 49184
rect 173860 49172 173866 49224
rect 208210 49172 208216 49224
rect 208268 49212 208274 49224
rect 258902 49212 258908 49224
rect 208268 49184 258908 49212
rect 208268 49172 208274 49184
rect 258902 49172 258908 49184
rect 258960 49172 258966 49224
rect 157702 49104 157708 49156
rect 157760 49144 157766 49156
rect 165798 49144 165804 49156
rect 157760 49116 165804 49144
rect 157760 49104 157766 49116
rect 165798 49104 165804 49116
rect 165856 49104 165862 49156
rect 179598 49104 179604 49156
rect 179656 49144 179662 49156
rect 179874 49144 179880 49156
rect 179656 49116 179880 49144
rect 179656 49104 179662 49116
rect 179874 49104 179880 49116
rect 179932 49104 179938 49156
rect 186958 49104 186964 49156
rect 187016 49144 187022 49156
rect 187142 49144 187148 49156
rect 187016 49116 187148 49144
rect 187016 49104 187022 49116
rect 187142 49104 187148 49116
rect 187200 49104 187206 49156
rect 259178 49144 259184 49156
rect 213104 49116 259184 49144
rect 157610 49036 157616 49088
rect 157668 49076 157674 49088
rect 165522 49076 165528 49088
rect 157668 49048 165528 49076
rect 157668 49036 157674 49048
rect 165522 49036 165528 49048
rect 165580 49036 165586 49088
rect 172790 49036 172796 49088
rect 172848 49076 172854 49088
rect 177850 49076 177856 49088
rect 172848 49048 177856 49076
rect 172848 49036 172854 49048
rect 177850 49036 177856 49048
rect 177908 49036 177914 49088
rect 179782 49036 179788 49088
rect 179840 49036 179846 49088
rect 188062 49036 188068 49088
rect 188120 49076 188126 49088
rect 188120 49048 200804 49076
rect 188120 49036 188126 49048
rect 161382 48968 161388 49020
rect 161440 49008 161446 49020
rect 176194 49008 176200 49020
rect 161440 48980 176200 49008
rect 161440 48968 161446 48980
rect 176194 48968 176200 48980
rect 176252 48968 176258 49020
rect 179598 48968 179604 49020
rect 179656 49008 179662 49020
rect 179800 49008 179828 49036
rect 179656 48980 179828 49008
rect 179656 48968 179662 48980
rect 187326 48968 187332 49020
rect 187384 49008 187390 49020
rect 187384 48980 195974 49008
rect 187384 48968 187390 48980
rect 173250 48900 173256 48952
rect 173308 48940 173314 48952
rect 177942 48940 177948 48952
rect 173308 48912 177948 48940
rect 173308 48900 173314 48912
rect 177942 48900 177948 48912
rect 178000 48900 178006 48952
rect 179414 48900 179420 48952
rect 179472 48940 179478 48952
rect 179782 48940 179788 48952
rect 179472 48912 179788 48940
rect 179472 48900 179478 48912
rect 179782 48900 179788 48912
rect 179840 48900 179846 48952
rect 182358 48900 182364 48952
rect 182416 48940 182422 48952
rect 184566 48940 184572 48952
rect 182416 48912 184572 48940
rect 182416 48900 182422 48912
rect 184566 48900 184572 48912
rect 184624 48900 184630 48952
rect 161566 48832 161572 48884
rect 161624 48872 161630 48884
rect 162118 48872 162124 48884
rect 161624 48844 162124 48872
rect 161624 48832 161630 48844
rect 162118 48832 162124 48844
rect 162176 48832 162182 48884
rect 177114 48832 177120 48884
rect 177172 48872 177178 48884
rect 183922 48872 183928 48884
rect 177172 48844 183928 48872
rect 177172 48832 177178 48844
rect 183922 48832 183928 48844
rect 183980 48832 183986 48884
rect 186222 48832 186228 48884
rect 186280 48872 186286 48884
rect 187326 48872 187332 48884
rect 186280 48844 187332 48872
rect 186280 48832 186286 48844
rect 187326 48832 187332 48844
rect 187384 48832 187390 48884
rect 195946 48872 195974 48980
rect 197538 48900 197544 48952
rect 197596 48940 197602 48952
rect 198090 48940 198096 48952
rect 197596 48912 198096 48940
rect 197596 48900 197602 48912
rect 198090 48900 198096 48912
rect 198148 48900 198154 48952
rect 200776 48940 200804 49048
rect 209590 49036 209596 49088
rect 209648 49076 209654 49088
rect 213104 49076 213132 49116
rect 259178 49104 259184 49116
rect 259236 49104 259242 49156
rect 259270 49076 259276 49088
rect 209648 49048 213132 49076
rect 213196 49048 259276 49076
rect 209648 49036 209654 49048
rect 211982 49008 211988 49020
rect 207952 48980 211988 49008
rect 207952 48940 207980 48980
rect 211982 48968 211988 48980
rect 212040 48968 212046 49020
rect 200776 48912 207980 48940
rect 209130 48900 209136 48952
rect 209188 48940 209194 48952
rect 209774 48940 209780 48952
rect 209188 48912 209780 48940
rect 209188 48900 209194 48912
rect 209774 48900 209780 48912
rect 209832 48900 209838 48952
rect 210234 48900 210240 48952
rect 210292 48940 210298 48952
rect 210602 48940 210608 48952
rect 210292 48912 210608 48940
rect 210292 48900 210298 48912
rect 210602 48900 210608 48912
rect 210660 48900 210666 48952
rect 210878 48872 210884 48884
rect 195946 48844 210884 48872
rect 210878 48832 210884 48844
rect 210936 48832 210942 48884
rect 179322 48804 179328 48816
rect 157306 48776 179328 48804
rect 156874 48424 156880 48476
rect 156932 48464 156938 48476
rect 157306 48464 157334 48776
rect 179322 48764 179328 48776
rect 179380 48764 179386 48816
rect 196250 48764 196256 48816
rect 196308 48804 196314 48816
rect 196526 48804 196532 48816
rect 196308 48776 196532 48804
rect 196308 48764 196314 48776
rect 196526 48764 196532 48776
rect 196584 48764 196590 48816
rect 210050 48764 210056 48816
rect 210108 48804 210114 48816
rect 210418 48804 210424 48816
rect 210108 48776 210424 48804
rect 210108 48764 210114 48776
rect 210418 48764 210424 48776
rect 210476 48764 210482 48816
rect 211522 48764 211528 48816
rect 211580 48804 211586 48816
rect 211982 48804 211988 48816
rect 211580 48776 211988 48804
rect 211580 48764 211586 48776
rect 211982 48764 211988 48776
rect 212040 48764 212046 48816
rect 161750 48696 161756 48748
rect 161808 48736 161814 48748
rect 162026 48736 162032 48748
rect 161808 48708 162032 48736
rect 161808 48696 161814 48708
rect 162026 48696 162032 48708
rect 162084 48696 162090 48748
rect 163222 48696 163228 48748
rect 163280 48736 163286 48748
rect 163590 48736 163596 48748
rect 163280 48708 163596 48736
rect 163280 48696 163286 48708
rect 163590 48696 163596 48708
rect 163648 48696 163654 48748
rect 163682 48696 163688 48748
rect 163740 48696 163746 48748
rect 169018 48696 169024 48748
rect 169076 48736 169082 48748
rect 169478 48736 169484 48748
rect 169076 48708 169484 48736
rect 169076 48696 169082 48708
rect 169478 48696 169484 48708
rect 169536 48696 169542 48748
rect 177298 48696 177304 48748
rect 177356 48736 177362 48748
rect 183370 48736 183376 48748
rect 177356 48708 183376 48736
rect 177356 48696 177362 48708
rect 183370 48696 183376 48708
rect 183428 48696 183434 48748
rect 200022 48696 200028 48748
rect 200080 48736 200086 48748
rect 204438 48736 204444 48748
rect 200080 48708 204444 48736
rect 200080 48696 200086 48708
rect 204438 48696 204444 48708
rect 204496 48696 204502 48748
rect 205726 48696 205732 48748
rect 205784 48736 205790 48748
rect 213196 48736 213224 49048
rect 259270 49036 259276 49048
rect 259328 49036 259334 49088
rect 259362 49008 259368 49020
rect 205784 48708 213224 48736
rect 213288 48980 259368 49008
rect 205784 48696 205790 48708
rect 159634 48628 159640 48680
rect 159692 48668 159698 48680
rect 162762 48668 162768 48680
rect 159692 48640 162768 48668
rect 159692 48628 159698 48640
rect 162762 48628 162768 48640
rect 162820 48628 162826 48680
rect 163130 48628 163136 48680
rect 163188 48668 163194 48680
rect 163700 48668 163728 48696
rect 178678 48668 178684 48680
rect 163188 48640 163728 48668
rect 166966 48640 178684 48668
rect 163188 48628 163194 48640
rect 161474 48560 161480 48612
rect 161532 48600 161538 48612
rect 165246 48600 165252 48612
rect 161532 48572 165252 48600
rect 161532 48560 161538 48572
rect 165246 48560 165252 48572
rect 165304 48560 165310 48612
rect 159726 48492 159732 48544
rect 159784 48532 159790 48544
rect 163038 48532 163044 48544
rect 159784 48504 163044 48532
rect 159784 48492 159790 48504
rect 163038 48492 163044 48504
rect 163096 48492 163102 48544
rect 156932 48436 157334 48464
rect 156932 48424 156938 48436
rect 158438 48424 158444 48476
rect 158496 48464 158502 48476
rect 161198 48464 161204 48476
rect 158496 48436 161204 48464
rect 158496 48424 158502 48436
rect 161198 48424 161204 48436
rect 161256 48424 161262 48476
rect 163590 48424 163596 48476
rect 163648 48464 163654 48476
rect 164510 48464 164516 48476
rect 163648 48436 164516 48464
rect 163648 48424 163654 48436
rect 164510 48424 164516 48436
rect 164568 48424 164574 48476
rect 164786 48424 164792 48476
rect 164844 48464 164850 48476
rect 165246 48464 165252 48476
rect 164844 48436 165252 48464
rect 164844 48424 164850 48436
rect 165246 48424 165252 48436
rect 165304 48424 165310 48476
rect 155218 48356 155224 48408
rect 155276 48396 155282 48408
rect 166966 48396 166994 48640
rect 178678 48628 178684 48640
rect 178736 48628 178742 48680
rect 179046 48628 179052 48680
rect 179104 48668 179110 48680
rect 183738 48668 183744 48680
rect 179104 48640 183744 48668
rect 179104 48628 179110 48640
rect 183738 48628 183744 48640
rect 183796 48628 183802 48680
rect 186682 48628 186688 48680
rect 186740 48668 186746 48680
rect 188614 48668 188620 48680
rect 186740 48640 188620 48668
rect 186740 48628 186746 48640
rect 188614 48628 188620 48640
rect 188672 48628 188678 48680
rect 197354 48628 197360 48680
rect 197412 48668 197418 48680
rect 197998 48668 198004 48680
rect 197412 48640 198004 48668
rect 197412 48628 197418 48640
rect 197998 48628 198004 48640
rect 198056 48628 198062 48680
rect 199194 48628 199200 48680
rect 199252 48668 199258 48680
rect 203978 48668 203984 48680
rect 199252 48640 203984 48668
rect 199252 48628 199258 48640
rect 203978 48628 203984 48640
rect 204036 48628 204042 48680
rect 206278 48628 206284 48680
rect 206336 48668 206342 48680
rect 213288 48668 213316 48980
rect 259362 48968 259368 48980
rect 259420 48968 259426 49020
rect 214006 48900 214012 48952
rect 214064 48940 214070 48952
rect 216122 48940 216128 48952
rect 214064 48912 216128 48940
rect 214064 48900 214070 48912
rect 216122 48900 216128 48912
rect 216180 48900 216186 48952
rect 215294 48832 215300 48884
rect 215352 48872 215358 48884
rect 215754 48872 215760 48884
rect 215352 48844 215760 48872
rect 215352 48832 215358 48844
rect 215754 48832 215760 48844
rect 215812 48832 215818 48884
rect 214098 48764 214104 48816
rect 214156 48804 214162 48816
rect 214282 48804 214288 48816
rect 214156 48776 214288 48804
rect 214156 48764 214162 48776
rect 214282 48764 214288 48776
rect 214340 48764 214346 48816
rect 214374 48764 214380 48816
rect 214432 48804 214438 48816
rect 214926 48804 214932 48816
rect 214432 48776 214932 48804
rect 214432 48764 214438 48776
rect 214926 48764 214932 48776
rect 214984 48764 214990 48816
rect 215570 48764 215576 48816
rect 215628 48804 215634 48816
rect 216030 48804 216036 48816
rect 215628 48776 216036 48804
rect 215628 48764 215634 48776
rect 216030 48764 216036 48776
rect 216088 48764 216094 48816
rect 214006 48696 214012 48748
rect 214064 48736 214070 48748
rect 214742 48736 214748 48748
rect 214064 48708 214748 48736
rect 214064 48696 214070 48708
rect 214742 48696 214748 48708
rect 214800 48696 214806 48748
rect 206336 48640 213316 48668
rect 206336 48628 206342 48640
rect 215662 48628 215668 48680
rect 215720 48668 215726 48680
rect 215938 48668 215944 48680
rect 215720 48640 215944 48668
rect 215720 48628 215726 48640
rect 215938 48628 215944 48640
rect 215996 48628 216002 48680
rect 254578 48600 254584 48612
rect 176626 48572 254584 48600
rect 172054 48492 172060 48544
rect 172112 48532 172118 48544
rect 176626 48532 176654 48572
rect 254578 48560 254584 48572
rect 254636 48560 254642 48612
rect 172112 48504 176654 48532
rect 172112 48492 172118 48504
rect 177666 48492 177672 48544
rect 177724 48532 177730 48544
rect 179782 48532 179788 48544
rect 177724 48504 179788 48532
rect 177724 48492 177730 48504
rect 179782 48492 179788 48504
rect 179840 48492 179846 48544
rect 184198 48492 184204 48544
rect 184256 48532 184262 48544
rect 185026 48532 185032 48544
rect 184256 48504 185032 48532
rect 184256 48492 184262 48504
rect 185026 48492 185032 48504
rect 185084 48492 185090 48544
rect 208302 48532 208308 48544
rect 186286 48504 208308 48532
rect 173618 48424 173624 48476
rect 173676 48464 173682 48476
rect 186286 48464 186314 48504
rect 208302 48492 208308 48504
rect 208360 48492 208366 48544
rect 210142 48492 210148 48544
rect 210200 48532 210206 48544
rect 210970 48532 210976 48544
rect 210200 48504 210976 48532
rect 210200 48492 210206 48504
rect 210970 48492 210976 48504
rect 211028 48492 211034 48544
rect 212534 48492 212540 48544
rect 212592 48532 212598 48544
rect 213178 48532 213184 48544
rect 212592 48504 213184 48532
rect 212592 48492 212598 48504
rect 213178 48492 213184 48504
rect 213236 48492 213242 48544
rect 214190 48492 214196 48544
rect 214248 48532 214254 48544
rect 214466 48532 214472 48544
rect 214248 48504 214472 48532
rect 214248 48492 214254 48504
rect 214466 48492 214472 48504
rect 214524 48492 214530 48544
rect 173676 48436 186314 48464
rect 173676 48424 173682 48436
rect 196066 48424 196072 48476
rect 196124 48464 196130 48476
rect 199838 48464 199844 48476
rect 196124 48436 199844 48464
rect 196124 48424 196130 48436
rect 199838 48424 199844 48436
rect 199896 48424 199902 48476
rect 200114 48424 200120 48476
rect 200172 48464 200178 48476
rect 203886 48464 203892 48476
rect 200172 48436 203892 48464
rect 200172 48424 200178 48436
rect 203886 48424 203892 48436
rect 203944 48424 203950 48476
rect 208118 48424 208124 48476
rect 208176 48464 208182 48476
rect 215938 48464 215944 48476
rect 208176 48436 215944 48464
rect 208176 48424 208182 48436
rect 215938 48424 215944 48436
rect 215996 48424 216002 48476
rect 155276 48368 166994 48396
rect 155276 48356 155282 48368
rect 179138 48356 179144 48408
rect 179196 48396 179202 48408
rect 179966 48396 179972 48408
rect 179196 48368 179972 48396
rect 179196 48356 179202 48368
rect 179966 48356 179972 48368
rect 180024 48356 180030 48408
rect 180518 48356 180524 48408
rect 180576 48396 180582 48408
rect 184014 48396 184020 48408
rect 180576 48368 184020 48396
rect 180576 48356 180582 48368
rect 184014 48356 184020 48368
rect 184072 48356 184078 48408
rect 198274 48356 198280 48408
rect 198332 48396 198338 48408
rect 202506 48396 202512 48408
rect 198332 48368 202512 48396
rect 198332 48356 198338 48368
rect 202506 48356 202512 48368
rect 202564 48356 202570 48408
rect 203150 48356 203156 48408
rect 203208 48396 203214 48408
rect 204622 48396 204628 48408
rect 203208 48368 204628 48396
rect 203208 48356 203214 48368
rect 204622 48356 204628 48368
rect 204680 48356 204686 48408
rect 210878 48356 210884 48408
rect 210936 48396 210942 48408
rect 216674 48396 216680 48408
rect 210936 48368 216680 48396
rect 210936 48356 210942 48368
rect 216674 48356 216680 48368
rect 216732 48356 216738 48408
rect 164418 48288 164424 48340
rect 164476 48328 164482 48340
rect 164970 48328 164976 48340
rect 164476 48300 164976 48328
rect 164476 48288 164482 48300
rect 164970 48288 164976 48300
rect 165028 48288 165034 48340
rect 179230 48288 179236 48340
rect 179288 48328 179294 48340
rect 179506 48328 179512 48340
rect 179288 48300 179512 48328
rect 179288 48288 179294 48300
rect 179506 48288 179512 48300
rect 179564 48288 179570 48340
rect 196526 48288 196532 48340
rect 196584 48328 196590 48340
rect 196986 48328 196992 48340
rect 196584 48300 196992 48328
rect 196584 48288 196590 48300
rect 196986 48288 196992 48300
rect 197044 48288 197050 48340
rect 202046 48288 202052 48340
rect 202104 48328 202110 48340
rect 203702 48328 203708 48340
rect 202104 48300 203708 48328
rect 202104 48288 202110 48300
rect 203702 48288 203708 48300
rect 203760 48288 203766 48340
rect 213178 48288 213184 48340
rect 213236 48328 213242 48340
rect 213546 48328 213552 48340
rect 213236 48300 213552 48328
rect 213236 48288 213242 48300
rect 213546 48288 213552 48300
rect 213604 48288 213610 48340
rect 214374 48288 214380 48340
rect 214432 48328 214438 48340
rect 216306 48328 216312 48340
rect 214432 48300 216312 48328
rect 214432 48288 214438 48300
rect 216306 48288 216312 48300
rect 216364 48288 216370 48340
rect 178402 48260 178408 48272
rect 157306 48232 178408 48260
rect 156966 48084 156972 48136
rect 157024 48124 157030 48136
rect 157306 48124 157334 48232
rect 178402 48220 178408 48232
rect 178460 48220 178466 48272
rect 251818 48260 251824 48272
rect 181456 48232 251824 48260
rect 162118 48152 162124 48204
rect 162176 48192 162182 48204
rect 162486 48192 162492 48204
rect 162176 48164 162492 48192
rect 162176 48152 162182 48164
rect 162486 48152 162492 48164
rect 162544 48152 162550 48204
rect 162854 48152 162860 48204
rect 162912 48192 162918 48204
rect 164234 48192 164240 48204
rect 162912 48164 164240 48192
rect 162912 48152 162918 48164
rect 164234 48152 164240 48164
rect 164292 48152 164298 48204
rect 164786 48152 164792 48204
rect 164844 48192 164850 48204
rect 165614 48192 165620 48204
rect 164844 48164 165620 48192
rect 164844 48152 164850 48164
rect 165614 48152 165620 48164
rect 165672 48152 165678 48204
rect 175182 48152 175188 48204
rect 175240 48192 175246 48204
rect 181456 48192 181484 48232
rect 251818 48220 251824 48232
rect 251876 48220 251882 48272
rect 243630 48192 243636 48204
rect 175240 48164 181484 48192
rect 186286 48164 243636 48192
rect 175240 48152 175246 48164
rect 157024 48096 157334 48124
rect 157024 48084 157030 48096
rect 161658 48084 161664 48136
rect 161716 48124 161722 48136
rect 162394 48124 162400 48136
rect 161716 48096 162400 48124
rect 161716 48084 161722 48096
rect 162394 48084 162400 48096
rect 162452 48084 162458 48136
rect 165062 48084 165068 48136
rect 165120 48124 165126 48136
rect 165338 48124 165344 48136
rect 165120 48096 165344 48124
rect 165120 48084 165126 48096
rect 165338 48084 165344 48096
rect 165396 48084 165402 48136
rect 174722 48084 174728 48136
rect 174780 48124 174786 48136
rect 186286 48124 186314 48164
rect 243630 48152 243636 48164
rect 243688 48152 243694 48204
rect 174780 48096 186314 48124
rect 174780 48084 174786 48096
rect 201494 48084 201500 48136
rect 201552 48124 201558 48136
rect 253658 48124 253664 48136
rect 201552 48096 253664 48124
rect 201552 48084 201558 48096
rect 253658 48084 253664 48096
rect 253716 48084 253722 48136
rect 156782 48016 156788 48068
rect 156840 48056 156846 48068
rect 178218 48056 178224 48068
rect 156840 48028 178224 48056
rect 156840 48016 156846 48028
rect 178218 48016 178224 48028
rect 178276 48016 178282 48068
rect 180794 48016 180800 48068
rect 180852 48056 180858 48068
rect 183830 48056 183836 48068
rect 180852 48028 183836 48056
rect 180852 48016 180858 48028
rect 183830 48016 183836 48028
rect 183888 48016 183894 48068
rect 190638 48016 190644 48068
rect 190696 48056 190702 48068
rect 190822 48056 190828 48068
rect 190696 48028 190828 48056
rect 190696 48016 190702 48028
rect 190822 48016 190828 48028
rect 190880 48016 190886 48068
rect 190914 48016 190920 48068
rect 190972 48056 190978 48068
rect 191374 48056 191380 48068
rect 190972 48028 191380 48056
rect 190972 48016 190978 48028
rect 191374 48016 191380 48028
rect 191432 48016 191438 48068
rect 196158 48016 196164 48068
rect 196216 48056 196222 48068
rect 196434 48056 196440 48068
rect 196216 48028 196440 48056
rect 196216 48016 196222 48028
rect 196434 48016 196440 48028
rect 196492 48016 196498 48068
rect 205634 48016 205640 48068
rect 205692 48056 205698 48068
rect 259086 48056 259092 48068
rect 205692 48028 259092 48056
rect 205692 48016 205698 48028
rect 259086 48016 259092 48028
rect 259144 48016 259150 48068
rect 146938 47948 146944 48000
rect 146996 47988 147002 48000
rect 176838 47988 176844 48000
rect 146996 47960 176844 47988
rect 146996 47948 147002 47960
rect 176838 47948 176844 47960
rect 176896 47948 176902 48000
rect 179598 47948 179604 48000
rect 179656 47988 179662 48000
rect 180610 47988 180616 48000
rect 179656 47960 180616 47988
rect 179656 47948 179662 47960
rect 180610 47948 180616 47960
rect 180668 47948 180674 48000
rect 189902 47948 189908 48000
rect 189960 47988 189966 48000
rect 244274 47988 244280 48000
rect 189960 47960 244280 47988
rect 189960 47948 189966 47960
rect 244274 47948 244280 47960
rect 244332 47948 244338 48000
rect 164694 47880 164700 47932
rect 164752 47920 164758 47932
rect 165430 47920 165436 47932
rect 164752 47892 165436 47920
rect 164752 47880 164758 47892
rect 165430 47880 165436 47892
rect 165488 47880 165494 47932
rect 169110 47880 169116 47932
rect 169168 47920 169174 47932
rect 169754 47920 169760 47932
rect 169168 47892 169760 47920
rect 169168 47880 169174 47892
rect 169754 47880 169760 47892
rect 169812 47880 169818 47932
rect 179690 47880 179696 47932
rect 179748 47920 179754 47932
rect 180058 47920 180064 47932
rect 179748 47892 180064 47920
rect 179748 47880 179754 47892
rect 180058 47880 180064 47892
rect 180116 47880 180122 47932
rect 190362 47880 190368 47932
rect 190420 47920 190426 47932
rect 248414 47920 248420 47932
rect 190420 47892 248420 47920
rect 190420 47880 190426 47892
rect 248414 47880 248420 47892
rect 248472 47880 248478 47932
rect 190454 47812 190460 47864
rect 190512 47852 190518 47864
rect 251174 47852 251180 47864
rect 190512 47824 251180 47852
rect 190512 47812 190518 47824
rect 251174 47812 251180 47824
rect 251232 47812 251238 47864
rect 159358 47744 159364 47796
rect 159416 47784 159422 47796
rect 169662 47784 169668 47796
rect 159416 47756 169668 47784
rect 159416 47744 159422 47756
rect 169662 47744 169668 47756
rect 169720 47744 169726 47796
rect 195698 47744 195704 47796
rect 195756 47784 195762 47796
rect 256418 47784 256424 47796
rect 195756 47756 256424 47784
rect 195756 47744 195762 47756
rect 256418 47744 256424 47756
rect 256476 47744 256482 47796
rect 134518 47676 134524 47728
rect 134576 47716 134582 47728
rect 160830 47716 160836 47728
rect 134576 47688 160836 47716
rect 134576 47676 134582 47688
rect 160830 47676 160836 47688
rect 160888 47676 160894 47728
rect 191926 47676 191932 47728
rect 191984 47716 191990 47728
rect 255958 47716 255964 47728
rect 191984 47688 255964 47716
rect 191984 47676 191990 47688
rect 255958 47676 255964 47688
rect 256016 47676 256022 47728
rect 134610 47608 134616 47660
rect 134668 47648 134674 47660
rect 168282 47648 168288 47660
rect 134668 47620 168288 47648
rect 134668 47608 134674 47620
rect 168282 47608 168288 47620
rect 168340 47608 168346 47660
rect 192018 47608 192024 47660
rect 192076 47648 192082 47660
rect 256510 47648 256516 47660
rect 192076 47620 256516 47648
rect 192076 47608 192082 47620
rect 256510 47608 256516 47620
rect 256568 47608 256574 47660
rect 133138 47540 133144 47592
rect 133196 47580 133202 47592
rect 166718 47580 166724 47592
rect 133196 47552 166724 47580
rect 133196 47540 133202 47552
rect 166718 47540 166724 47552
rect 166776 47540 166782 47592
rect 167270 47540 167276 47592
rect 167328 47580 167334 47592
rect 167638 47580 167644 47592
rect 167328 47552 167644 47580
rect 167328 47540 167334 47552
rect 167638 47540 167644 47552
rect 167696 47540 167702 47592
rect 173250 47540 173256 47592
rect 173308 47580 173314 47592
rect 182634 47580 182640 47592
rect 173308 47552 182640 47580
rect 173308 47540 173314 47552
rect 182634 47540 182640 47552
rect 182692 47540 182698 47592
rect 191558 47540 191564 47592
rect 191616 47580 191622 47592
rect 255314 47580 255320 47592
rect 191616 47552 255320 47580
rect 191616 47540 191622 47552
rect 255314 47540 255320 47552
rect 255372 47540 255378 47592
rect 152458 47472 152464 47524
rect 152516 47512 152522 47524
rect 177758 47512 177764 47524
rect 152516 47484 177764 47512
rect 152516 47472 152522 47484
rect 177758 47472 177764 47484
rect 177816 47472 177822 47524
rect 193214 47472 193220 47524
rect 193272 47512 193278 47524
rect 193858 47512 193864 47524
rect 193272 47484 193864 47512
rect 193272 47472 193278 47484
rect 193858 47472 193864 47484
rect 193916 47472 193922 47524
rect 203058 47472 203064 47524
rect 203116 47512 203122 47524
rect 253750 47512 253756 47524
rect 203116 47484 253756 47512
rect 203116 47472 203122 47484
rect 253750 47472 253756 47484
rect 253808 47472 253814 47524
rect 136542 47404 136548 47456
rect 136600 47444 136606 47456
rect 143074 47444 143080 47456
rect 136600 47416 143080 47444
rect 136600 47404 136606 47416
rect 143074 47404 143080 47416
rect 143132 47404 143138 47456
rect 159542 47404 159548 47456
rect 159600 47444 159606 47456
rect 160278 47444 160284 47456
rect 159600 47416 160284 47444
rect 159600 47404 159606 47416
rect 160278 47404 160284 47416
rect 160336 47404 160342 47456
rect 163222 47404 163228 47456
rect 163280 47444 163286 47456
rect 164142 47444 164148 47456
rect 163280 47416 164148 47444
rect 163280 47404 163286 47416
rect 164142 47404 164148 47416
rect 164200 47404 164206 47456
rect 167454 47404 167460 47456
rect 167512 47444 167518 47456
rect 167730 47444 167736 47456
rect 167512 47416 167736 47444
rect 167512 47404 167518 47416
rect 167730 47404 167736 47416
rect 167788 47404 167794 47456
rect 176654 47404 176660 47456
rect 176712 47444 176718 47456
rect 181806 47444 181812 47456
rect 176712 47416 181812 47444
rect 176712 47404 176718 47416
rect 181806 47404 181812 47416
rect 181864 47404 181870 47456
rect 189350 47404 189356 47456
rect 189408 47444 189414 47456
rect 190362 47444 190368 47456
rect 189408 47416 190368 47444
rect 189408 47404 189414 47416
rect 190362 47404 190368 47416
rect 190420 47404 190426 47456
rect 193674 47404 193680 47456
rect 193732 47444 193738 47456
rect 194594 47444 194600 47456
rect 193732 47416 194600 47444
rect 193732 47404 193738 47416
rect 194594 47404 194600 47416
rect 194652 47404 194658 47456
rect 194778 47404 194784 47456
rect 194836 47444 194842 47456
rect 195514 47444 195520 47456
rect 194836 47416 195520 47444
rect 194836 47404 194842 47416
rect 195514 47404 195520 47416
rect 195572 47404 195578 47456
rect 196158 47404 196164 47456
rect 196216 47444 196222 47456
rect 197078 47444 197084 47456
rect 196216 47416 197084 47444
rect 196216 47404 196222 47416
rect 197078 47404 197084 47416
rect 197136 47404 197142 47456
rect 205818 47404 205824 47456
rect 205876 47444 205882 47456
rect 224218 47444 224224 47456
rect 205876 47416 224224 47444
rect 205876 47404 205882 47416
rect 224218 47404 224224 47416
rect 224276 47404 224282 47456
rect 175458 47336 175464 47388
rect 175516 47376 175522 47388
rect 218146 47376 218152 47388
rect 175516 47348 218152 47376
rect 175516 47336 175522 47348
rect 218146 47336 218152 47348
rect 218204 47336 218210 47388
rect 166994 47268 167000 47320
rect 167052 47308 167058 47320
rect 167822 47308 167828 47320
rect 167052 47280 167828 47308
rect 167052 47268 167058 47280
rect 167822 47268 167828 47280
rect 167880 47268 167886 47320
rect 178862 47268 178868 47320
rect 178920 47308 178926 47320
rect 184382 47308 184388 47320
rect 178920 47280 184388 47308
rect 178920 47268 178926 47280
rect 184382 47268 184388 47280
rect 184440 47268 184446 47320
rect 189442 47268 189448 47320
rect 189500 47308 189506 47320
rect 190178 47308 190184 47320
rect 189500 47280 190184 47308
rect 189500 47268 189506 47280
rect 190178 47268 190184 47280
rect 190236 47268 190242 47320
rect 177758 47200 177764 47252
rect 177816 47240 177822 47252
rect 181530 47240 181536 47252
rect 177816 47212 181536 47240
rect 177816 47200 177822 47212
rect 181530 47200 181536 47212
rect 181588 47200 181594 47252
rect 177482 47132 177488 47184
rect 177540 47172 177546 47184
rect 180886 47172 180892 47184
rect 177540 47144 180892 47172
rect 177540 47132 177546 47144
rect 180886 47132 180892 47144
rect 180944 47132 180950 47184
rect 181254 47132 181260 47184
rect 181312 47172 181318 47184
rect 181438 47172 181444 47184
rect 181312 47144 181444 47172
rect 181312 47132 181318 47144
rect 181438 47132 181444 47144
rect 181496 47132 181502 47184
rect 184382 47132 184388 47184
rect 184440 47172 184446 47184
rect 184842 47172 184848 47184
rect 184440 47144 184848 47172
rect 184440 47132 184446 47144
rect 184842 47132 184848 47144
rect 184900 47132 184906 47184
rect 178678 47064 178684 47116
rect 178736 47104 178742 47116
rect 183278 47104 183284 47116
rect 178736 47076 183284 47104
rect 178736 47064 178742 47076
rect 183278 47064 183284 47076
rect 183336 47064 183342 47116
rect 198826 47064 198832 47116
rect 198884 47104 198890 47116
rect 199194 47104 199200 47116
rect 198884 47076 199200 47104
rect 198884 47064 198890 47076
rect 199194 47064 199200 47076
rect 199252 47064 199258 47116
rect 178770 46996 178776 47048
rect 178828 47036 178834 47048
rect 181898 47036 181904 47048
rect 178828 47008 181904 47036
rect 178828 46996 178834 47008
rect 181898 46996 181904 47008
rect 181956 46996 181962 47048
rect 159450 46928 159456 46980
rect 159508 46968 159514 46980
rect 163406 46968 163412 46980
rect 159508 46940 163412 46968
rect 159508 46928 159514 46940
rect 163406 46928 163412 46940
rect 163464 46928 163470 46980
rect 168558 46928 168564 46980
rect 168616 46968 168622 46980
rect 169202 46968 169208 46980
rect 168616 46940 169208 46968
rect 168616 46928 168622 46940
rect 169202 46928 169208 46940
rect 169260 46928 169266 46980
rect 177574 46928 177580 46980
rect 177632 46968 177638 46980
rect 180334 46968 180340 46980
rect 177632 46940 180340 46968
rect 177632 46928 177638 46940
rect 180334 46928 180340 46940
rect 180392 46928 180398 46980
rect 183554 46928 183560 46980
rect 183612 46968 183618 46980
rect 184934 46968 184940 46980
rect 183612 46940 184940 46968
rect 183612 46928 183618 46940
rect 184934 46928 184940 46940
rect 184992 46928 184998 46980
rect 185854 46928 185860 46980
rect 185912 46968 185918 46980
rect 186038 46968 186044 46980
rect 185912 46940 186044 46968
rect 185912 46928 185918 46940
rect 186038 46928 186044 46940
rect 186096 46928 186102 46980
rect 186958 46928 186964 46980
rect 187016 46968 187022 46980
rect 190086 46968 190092 46980
rect 187016 46940 190092 46968
rect 187016 46928 187022 46940
rect 190086 46928 190092 46940
rect 190144 46928 190150 46980
rect 204622 46928 204628 46980
rect 204680 46968 204686 46980
rect 205174 46968 205180 46980
rect 204680 46940 205180 46968
rect 204680 46928 204686 46940
rect 205174 46928 205180 46940
rect 205232 46928 205238 46980
rect 172974 46860 172980 46912
rect 173032 46900 173038 46912
rect 247678 46900 247684 46912
rect 173032 46872 247684 46900
rect 173032 46860 173038 46872
rect 247678 46860 247684 46872
rect 247736 46860 247742 46912
rect 167362 46792 167368 46844
rect 167420 46832 167426 46844
rect 168098 46832 168104 46844
rect 167420 46804 168104 46832
rect 167420 46792 167426 46804
rect 168098 46792 168104 46804
rect 168156 46792 168162 46844
rect 173526 46792 173532 46844
rect 173584 46832 173590 46844
rect 240870 46832 240876 46844
rect 173584 46804 240876 46832
rect 173584 46792 173590 46804
rect 240870 46792 240876 46804
rect 240928 46792 240934 46844
rect 151262 46724 151268 46776
rect 151320 46764 151326 46776
rect 178586 46764 178592 46776
rect 151320 46736 178592 46764
rect 151320 46724 151326 46736
rect 178586 46724 178592 46736
rect 178644 46724 178650 46776
rect 204346 46724 204352 46776
rect 204404 46764 204410 46776
rect 204622 46764 204628 46776
rect 204404 46736 204628 46764
rect 204404 46724 204410 46736
rect 204622 46724 204628 46736
rect 204680 46724 204686 46776
rect 153838 46656 153844 46708
rect 153896 46696 153902 46708
rect 177206 46696 177212 46708
rect 153896 46668 177212 46696
rect 153896 46656 153902 46668
rect 177206 46656 177212 46668
rect 177264 46656 177270 46708
rect 188430 46656 188436 46708
rect 188488 46696 188494 46708
rect 188488 46668 195974 46696
rect 188488 46656 188494 46668
rect 151170 46588 151176 46640
rect 151228 46628 151234 46640
rect 177390 46628 177396 46640
rect 151228 46600 177396 46628
rect 151228 46588 151234 46600
rect 177390 46588 177396 46600
rect 177448 46588 177454 46640
rect 189534 46588 189540 46640
rect 189592 46628 189598 46640
rect 189592 46600 195836 46628
rect 189592 46588 189598 46600
rect 161842 46520 161848 46572
rect 161900 46560 161906 46572
rect 162210 46560 162216 46572
rect 161900 46532 162216 46560
rect 161900 46520 161906 46532
rect 162210 46520 162216 46532
rect 162268 46520 162274 46572
rect 191006 46520 191012 46572
rect 191064 46560 191070 46572
rect 191064 46532 195744 46560
rect 191064 46520 191070 46532
rect 138658 46452 138664 46504
rect 138716 46492 138722 46504
rect 159910 46492 159916 46504
rect 138716 46464 159916 46492
rect 138716 46452 138722 46464
rect 159910 46452 159916 46464
rect 159968 46452 159974 46504
rect 185210 46452 185216 46504
rect 185268 46492 185274 46504
rect 185854 46492 185860 46504
rect 185268 46464 185860 46492
rect 185268 46452 185274 46464
rect 185854 46452 185860 46464
rect 185912 46452 185918 46504
rect 153194 46384 153200 46436
rect 153252 46424 153258 46436
rect 182910 46424 182916 46436
rect 153252 46396 182916 46424
rect 153252 46384 153258 46396
rect 182910 46384 182916 46396
rect 182968 46384 182974 46436
rect 186774 46384 186780 46436
rect 186832 46424 186838 46436
rect 191006 46424 191012 46436
rect 186832 46396 191012 46424
rect 186832 46384 186838 46396
rect 191006 46384 191012 46396
rect 191064 46384 191070 46436
rect 134702 46316 134708 46368
rect 134760 46356 134766 46368
rect 168374 46356 168380 46368
rect 134760 46328 168380 46356
rect 134760 46316 134766 46328
rect 168374 46316 168380 46328
rect 168432 46316 168438 46368
rect 171318 46316 171324 46368
rect 171376 46356 171382 46368
rect 171502 46356 171508 46368
rect 171376 46328 171508 46356
rect 171376 46316 171382 46328
rect 171502 46316 171508 46328
rect 171560 46316 171566 46368
rect 175274 46316 175280 46368
rect 175332 46356 175338 46368
rect 182358 46356 182364 46368
rect 175332 46328 182364 46356
rect 175332 46316 175338 46328
rect 182358 46316 182364 46328
rect 182416 46316 182422 46368
rect 185210 46316 185216 46368
rect 185268 46356 185274 46368
rect 185762 46356 185768 46368
rect 185268 46328 185768 46356
rect 185268 46316 185274 46328
rect 185762 46316 185768 46328
rect 185820 46316 185826 46368
rect 190454 46316 190460 46368
rect 190512 46356 190518 46368
rect 191190 46356 191196 46368
rect 190512 46328 191196 46356
rect 190512 46316 190518 46328
rect 191190 46316 191196 46328
rect 191248 46316 191254 46368
rect 143534 46248 143540 46300
rect 143592 46288 143598 46300
rect 182082 46288 182088 46300
rect 143592 46260 182088 46288
rect 143592 46248 143598 46260
rect 182082 46248 182088 46260
rect 182140 46248 182146 46300
rect 182910 46248 182916 46300
rect 182968 46288 182974 46300
rect 183462 46288 183468 46300
rect 182968 46260 183468 46288
rect 182968 46248 182974 46260
rect 183462 46248 183468 46260
rect 183520 46248 183526 46300
rect 186590 46248 186596 46300
rect 186648 46288 186654 46300
rect 188522 46288 188528 46300
rect 186648 46260 188528 46288
rect 186648 46248 186654 46260
rect 188522 46248 188528 46260
rect 188580 46248 188586 46300
rect 190730 46248 190736 46300
rect 190788 46288 190794 46300
rect 191282 46288 191288 46300
rect 190788 46260 191288 46288
rect 190788 46248 190794 46260
rect 191282 46248 191288 46260
rect 191340 46248 191346 46300
rect 135990 46180 135996 46232
rect 136048 46220 136054 46232
rect 180242 46220 180248 46232
rect 136048 46192 180248 46220
rect 136048 46180 136054 46192
rect 180242 46180 180248 46192
rect 180300 46180 180306 46232
rect 185302 46180 185308 46232
rect 185360 46220 185366 46232
rect 185762 46220 185768 46232
rect 185360 46192 185768 46220
rect 185360 46180 185366 46192
rect 185762 46180 185768 46192
rect 185820 46180 185826 46232
rect 188062 46180 188068 46232
rect 188120 46220 188126 46232
rect 188706 46220 188712 46232
rect 188120 46192 188712 46220
rect 188120 46180 188126 46192
rect 188706 46180 188712 46192
rect 188764 46180 188770 46232
rect 192478 46180 192484 46232
rect 192536 46220 192542 46232
rect 192754 46220 192760 46232
rect 192536 46192 192760 46220
rect 192536 46180 192542 46192
rect 192754 46180 192760 46192
rect 192812 46180 192818 46232
rect 195716 46220 195744 46532
rect 195808 46288 195836 46600
rect 195946 46356 195974 46668
rect 201494 46656 201500 46708
rect 201552 46696 201558 46708
rect 201770 46696 201776 46708
rect 201552 46668 201776 46696
rect 201552 46656 201558 46668
rect 201770 46656 201776 46668
rect 201828 46656 201834 46708
rect 201402 46588 201408 46640
rect 201460 46628 201466 46640
rect 201862 46628 201868 46640
rect 201460 46600 201868 46628
rect 201460 46588 201466 46600
rect 201862 46588 201868 46600
rect 201920 46588 201926 46640
rect 211062 46520 211068 46572
rect 211120 46560 211126 46572
rect 211706 46560 211712 46572
rect 211120 46532 211712 46560
rect 211120 46520 211126 46532
rect 211706 46520 211712 46532
rect 211764 46520 211770 46572
rect 204438 46452 204444 46504
rect 204496 46492 204502 46504
rect 205266 46492 205272 46504
rect 204496 46464 205272 46492
rect 204496 46452 204502 46464
rect 205266 46452 205272 46464
rect 205324 46452 205330 46504
rect 211338 46452 211344 46504
rect 211396 46492 211402 46504
rect 211798 46492 211804 46504
rect 211396 46464 211804 46492
rect 211396 46452 211402 46464
rect 211798 46452 211804 46464
rect 211856 46452 211862 46504
rect 201586 46384 201592 46436
rect 201644 46424 201650 46436
rect 202322 46424 202328 46436
rect 201644 46396 202328 46424
rect 201644 46384 201650 46396
rect 202322 46384 202328 46396
rect 202380 46384 202386 46436
rect 204346 46384 204352 46436
rect 204404 46424 204410 46436
rect 204990 46424 204996 46436
rect 204404 46396 204996 46424
rect 204404 46384 204410 46396
rect 204990 46384 204996 46396
rect 205048 46384 205054 46436
rect 211154 46384 211160 46436
rect 211212 46424 211218 46436
rect 211706 46424 211712 46436
rect 211212 46396 211712 46424
rect 211212 46384 211218 46396
rect 211706 46384 211712 46396
rect 211764 46384 211770 46436
rect 212626 46384 212632 46436
rect 212684 46424 212690 46436
rect 212810 46424 212816 46436
rect 212684 46396 212816 46424
rect 212684 46384 212690 46396
rect 212810 46384 212816 46396
rect 212868 46384 212874 46436
rect 227714 46356 227720 46368
rect 195946 46328 227720 46356
rect 227714 46316 227720 46328
rect 227772 46316 227778 46368
rect 237374 46288 237380 46300
rect 195808 46260 237380 46288
rect 237374 46248 237380 46260
rect 237432 46248 237438 46300
rect 259454 46220 259460 46232
rect 195716 46192 259460 46220
rect 259454 46180 259460 46192
rect 259512 46180 259518 46232
rect 161934 46112 161940 46164
rect 161992 46152 161998 46164
rect 162578 46152 162584 46164
rect 161992 46124 162584 46152
rect 161992 46112 161998 46124
rect 162578 46112 162584 46124
rect 162636 46112 162642 46164
rect 166350 46112 166356 46164
rect 166408 46152 166414 46164
rect 166902 46152 166908 46164
rect 166408 46124 166908 46152
rect 166408 46112 166414 46124
rect 166902 46112 166908 46124
rect 166960 46112 166966 46164
rect 169754 46112 169760 46164
rect 169812 46152 169818 46164
rect 170030 46152 170036 46164
rect 169812 46124 170036 46152
rect 169812 46112 169818 46124
rect 170030 46112 170036 46124
rect 170088 46112 170094 46164
rect 171502 46112 171508 46164
rect 171560 46152 171566 46164
rect 171686 46152 171692 46164
rect 171560 46124 171692 46152
rect 171560 46112 171566 46124
rect 171686 46112 171692 46124
rect 171744 46112 171750 46164
rect 177482 46112 177488 46164
rect 177540 46152 177546 46164
rect 177758 46152 177764 46164
rect 177540 46124 177764 46152
rect 177540 46112 177546 46124
rect 177758 46112 177764 46124
rect 177816 46112 177822 46164
rect 197354 46112 197360 46164
rect 197412 46152 197418 46164
rect 198366 46152 198372 46164
rect 197412 46124 198372 46152
rect 197412 46112 197418 46124
rect 198366 46112 198372 46124
rect 198424 46112 198430 46164
rect 201678 46112 201684 46164
rect 201736 46152 201742 46164
rect 202046 46152 202052 46164
rect 201736 46124 202052 46152
rect 201736 46112 201742 46124
rect 202046 46112 202052 46124
rect 202104 46112 202110 46164
rect 203058 46112 203064 46164
rect 203116 46152 203122 46164
rect 203426 46152 203432 46164
rect 203116 46124 203432 46152
rect 203116 46112 203122 46124
rect 203426 46112 203432 46124
rect 203484 46112 203490 46164
rect 204438 46112 204444 46164
rect 204496 46152 204502 46164
rect 204714 46152 204720 46164
rect 204496 46124 204720 46152
rect 204496 46112 204502 46124
rect 204714 46112 204720 46124
rect 204772 46112 204778 46164
rect 205726 46112 205732 46164
rect 205784 46152 205790 46164
rect 206462 46152 206468 46164
rect 205784 46124 206468 46152
rect 205784 46112 205790 46124
rect 206462 46112 206468 46124
rect 206520 46112 206526 46164
rect 207106 46112 207112 46164
rect 207164 46152 207170 46164
rect 207934 46152 207940 46164
rect 207164 46124 207940 46152
rect 207164 46112 207170 46124
rect 207934 46112 207940 46124
rect 207992 46112 207998 46164
rect 210418 46112 210424 46164
rect 210476 46152 210482 46164
rect 210694 46152 210700 46164
rect 210476 46124 210700 46152
rect 210476 46112 210482 46124
rect 210694 46112 210700 46124
rect 210752 46112 210758 46164
rect 211798 46112 211804 46164
rect 211856 46152 211862 46164
rect 212074 46152 212080 46164
rect 211856 46124 212080 46152
rect 211856 46112 211862 46124
rect 212074 46112 212080 46124
rect 212132 46112 212138 46164
rect 212442 46112 212448 46164
rect 212500 46152 212506 46164
rect 212810 46152 212816 46164
rect 212500 46124 212816 46152
rect 212500 46112 212506 46124
rect 212810 46112 212816 46124
rect 212868 46112 212874 46164
rect 170122 46044 170128 46096
rect 170180 46084 170186 46096
rect 170950 46084 170956 46096
rect 170180 46056 170956 46084
rect 170180 46044 170186 46056
rect 170950 46044 170956 46056
rect 171008 46044 171014 46096
rect 185302 46044 185308 46096
rect 185360 46084 185366 46096
rect 185946 46084 185952 46096
rect 185360 46056 185952 46084
rect 185360 46044 185366 46056
rect 185946 46044 185952 46056
rect 186004 46044 186010 46096
rect 189258 46044 189264 46096
rect 189316 46084 189322 46096
rect 189994 46084 190000 46096
rect 189316 46056 190000 46084
rect 189316 46044 189322 46056
rect 189994 46044 190000 46056
rect 190052 46044 190058 46096
rect 193306 46044 193312 46096
rect 193364 46084 193370 46096
rect 193950 46084 193956 46096
rect 193364 46056 193956 46084
rect 193364 46044 193370 46056
rect 193950 46044 193956 46056
rect 194008 46044 194014 46096
rect 199102 46044 199108 46096
rect 199160 46084 199166 46096
rect 199562 46084 199568 46096
rect 199160 46056 199568 46084
rect 199160 46044 199166 46056
rect 199562 46044 199568 46056
rect 199620 46044 199626 46096
rect 200206 46044 200212 46096
rect 200264 46084 200270 46096
rect 201310 46084 201316 46096
rect 200264 46056 201316 46084
rect 200264 46044 200270 46056
rect 201310 46044 201316 46056
rect 201368 46044 201374 46096
rect 201494 46044 201500 46096
rect 201552 46084 201558 46096
rect 202230 46084 202236 46096
rect 201552 46056 202236 46084
rect 201552 46044 201558 46056
rect 202230 46044 202236 46056
rect 202288 46044 202294 46096
rect 202874 46044 202880 46096
rect 202932 46084 202938 46096
rect 203518 46084 203524 46096
rect 202932 46056 203524 46084
rect 202932 46044 202938 46056
rect 203518 46044 203524 46056
rect 203576 46044 203582 46096
rect 204254 46044 204260 46096
rect 204312 46084 204318 46096
rect 204806 46084 204812 46096
rect 204312 46056 204812 46084
rect 204312 46044 204318 46056
rect 204806 46044 204812 46056
rect 204864 46044 204870 46096
rect 205818 46044 205824 46096
rect 205876 46084 205882 46096
rect 206554 46084 206560 46096
rect 205876 46056 206560 46084
rect 205876 46044 205882 46056
rect 206554 46044 206560 46056
rect 206612 46044 206618 46096
rect 168926 45976 168932 46028
rect 168984 46016 168990 46028
rect 169570 46016 169576 46028
rect 168984 45988 169576 46016
rect 168984 45976 168990 45988
rect 169570 45976 169576 45988
rect 169628 45976 169634 46028
rect 170030 45976 170036 46028
rect 170088 46016 170094 46028
rect 170674 46016 170680 46028
rect 170088 45988 170680 46016
rect 170088 45976 170094 45988
rect 170674 45976 170680 45988
rect 170732 45976 170738 46028
rect 171134 45976 171140 46028
rect 171192 46016 171198 46028
rect 171686 46016 171692 46028
rect 171192 45988 171692 46016
rect 171192 45976 171198 45988
rect 171686 45976 171692 45988
rect 171744 45976 171750 46028
rect 198826 45976 198832 46028
rect 198884 46016 198890 46028
rect 199470 46016 199476 46028
rect 198884 45988 199476 46016
rect 198884 45976 198890 45988
rect 199470 45976 199476 45988
rect 199528 45976 199534 46028
rect 200298 45976 200304 46028
rect 200356 46016 200362 46028
rect 200666 46016 200672 46028
rect 200356 45988 200672 46016
rect 200356 45976 200362 45988
rect 200666 45976 200672 45988
rect 200724 45976 200730 46028
rect 200758 45976 200764 46028
rect 200816 46016 200822 46028
rect 201126 46016 201132 46028
rect 200816 45988 201132 46016
rect 200816 45976 200822 45988
rect 201126 45976 201132 45988
rect 201184 45976 201190 46028
rect 201678 45976 201684 46028
rect 201736 46016 201742 46028
rect 202414 46016 202420 46028
rect 201736 45988 202420 46016
rect 201736 45976 201742 45988
rect 202414 45976 202420 45988
rect 202472 45976 202478 46028
rect 204714 45976 204720 46028
rect 204772 46016 204778 46028
rect 205082 46016 205088 46028
rect 204772 45988 205088 46016
rect 204772 45976 204778 45988
rect 205082 45976 205088 45988
rect 205140 45976 205146 46028
rect 193306 45908 193312 45960
rect 193364 45948 193370 45960
rect 194134 45948 194140 45960
rect 193364 45920 194140 45948
rect 193364 45908 193370 45920
rect 194134 45908 194140 45920
rect 194192 45908 194198 45960
rect 207290 45908 207296 45960
rect 207348 45948 207354 45960
rect 207750 45948 207756 45960
rect 207348 45920 207756 45948
rect 207348 45908 207354 45920
rect 207750 45908 207756 45920
rect 207808 45908 207814 45960
rect 167730 45840 167736 45892
rect 167788 45880 167794 45892
rect 168190 45880 168196 45892
rect 167788 45852 168196 45880
rect 167788 45840 167794 45852
rect 168190 45840 168196 45852
rect 168248 45840 168254 45892
rect 198734 45840 198740 45892
rect 198792 45880 198798 45892
rect 199470 45880 199476 45892
rect 198792 45852 199476 45880
rect 198792 45840 198798 45852
rect 199470 45840 199476 45852
rect 199528 45840 199534 45892
rect 200298 45840 200304 45892
rect 200356 45880 200362 45892
rect 201218 45880 201224 45892
rect 200356 45852 201224 45880
rect 200356 45840 200362 45852
rect 201218 45840 201224 45852
rect 201276 45840 201282 45892
rect 211338 45772 211344 45824
rect 211396 45812 211402 45824
rect 212166 45812 212172 45824
rect 211396 45784 212172 45812
rect 211396 45772 211402 45784
rect 212166 45772 212172 45784
rect 212224 45772 212230 45824
rect 198734 45704 198740 45756
rect 198792 45744 198798 45756
rect 199654 45744 199660 45756
rect 198792 45716 199660 45744
rect 198792 45704 198798 45716
rect 199654 45704 199660 45716
rect 199712 45704 199718 45756
rect 135622 45500 135628 45552
rect 135680 45540 135686 45552
rect 138750 45540 138756 45552
rect 135680 45512 138756 45540
rect 135680 45500 135686 45512
rect 138750 45500 138756 45512
rect 138808 45500 138814 45552
rect 158714 45432 158720 45484
rect 158772 45472 158778 45484
rect 160002 45472 160008 45484
rect 158772 45444 160008 45472
rect 158772 45432 158778 45444
rect 160002 45432 160008 45444
rect 160060 45432 160066 45484
rect 185578 45228 185584 45280
rect 185636 45268 185642 45280
rect 189718 45268 189724 45280
rect 185636 45240 189724 45268
rect 185636 45228 185642 45240
rect 189718 45228 189724 45240
rect 189776 45228 189782 45280
rect 162946 45160 162952 45212
rect 163004 45200 163010 45212
rect 164050 45200 164056 45212
rect 163004 45172 164056 45200
rect 163004 45160 163010 45172
rect 164050 45160 164056 45172
rect 164108 45160 164114 45212
rect 168374 45024 168380 45076
rect 168432 45064 168438 45076
rect 177114 45064 177120 45076
rect 168432 45036 177120 45064
rect 168432 45024 168438 45036
rect 177114 45024 177120 45036
rect 177172 45024 177178 45076
rect 183094 45064 183100 45076
rect 177316 45036 183100 45064
rect 155954 44956 155960 45008
rect 156012 44996 156018 45008
rect 177316 44996 177344 45036
rect 183094 45024 183100 45036
rect 183152 45024 183158 45076
rect 181990 44996 181996 45008
rect 156012 44968 177344 44996
rect 177408 44968 181996 44996
rect 156012 44956 156018 44968
rect 143626 44888 143632 44940
rect 143684 44928 143690 44940
rect 177408 44928 177436 44968
rect 181990 44956 181996 44968
rect 182048 44956 182054 45008
rect 188430 44956 188436 45008
rect 188488 44996 188494 45008
rect 226334 44996 226340 45008
rect 188488 44968 226340 44996
rect 188488 44956 188494 44968
rect 226334 44956 226340 44968
rect 226392 44956 226398 45008
rect 143684 44900 177436 44928
rect 143684 44888 143690 44900
rect 178034 44888 178040 44940
rect 178092 44928 178098 44940
rect 184658 44928 184664 44940
rect 178092 44900 184664 44928
rect 178092 44888 178098 44900
rect 184658 44888 184664 44900
rect 184716 44888 184722 44940
rect 190270 44888 190276 44940
rect 190328 44928 190334 44940
rect 249794 44928 249800 44940
rect 190328 44900 249800 44928
rect 190328 44888 190334 44900
rect 249794 44888 249800 44900
rect 249852 44888 249858 44940
rect 139394 44820 139400 44872
rect 139452 44860 139458 44872
rect 181622 44860 181628 44872
rect 139452 44832 181628 44860
rect 139452 44820 139458 44832
rect 181622 44820 181628 44832
rect 181680 44820 181686 44872
rect 190914 44820 190920 44872
rect 190972 44860 190978 44872
rect 253934 44860 253940 44872
rect 190972 44832 253940 44860
rect 190972 44820 190978 44832
rect 253934 44820 253940 44832
rect 253992 44820 253998 44872
rect 203150 44412 203156 44464
rect 203208 44452 203214 44464
rect 203610 44452 203616 44464
rect 203208 44424 203616 44452
rect 203208 44412 203214 44424
rect 203610 44412 203616 44424
rect 203668 44412 203674 44464
rect 171134 44140 171140 44192
rect 171192 44180 171198 44192
rect 180518 44180 180524 44192
rect 171192 44152 180524 44180
rect 171192 44140 171198 44152
rect 180518 44140 180524 44152
rect 180576 44140 180582 44192
rect 203702 44140 203708 44192
rect 203760 44180 203766 44192
rect 203978 44180 203984 44192
rect 203760 44152 203984 44180
rect 203760 44140 203766 44152
rect 203978 44140 203984 44152
rect 204036 44140 204042 44192
rect 187602 44072 187608 44124
rect 187660 44112 187666 44124
rect 191098 44112 191104 44124
rect 187660 44084 191104 44112
rect 187660 44072 187666 44084
rect 191098 44072 191104 44084
rect 191156 44072 191162 44124
rect 208762 44004 208768 44056
rect 208820 44044 208826 44056
rect 209222 44044 209228 44056
rect 208820 44016 209228 44044
rect 208820 44004 208826 44016
rect 209222 44004 209228 44016
rect 209280 44004 209286 44056
rect 174814 43868 174820 43920
rect 174872 43908 174878 43920
rect 182818 43908 182824 43920
rect 174872 43880 182824 43908
rect 174872 43868 174878 43880
rect 182818 43868 182824 43880
rect 182876 43868 182882 43920
rect 208762 43868 208768 43920
rect 208820 43908 208826 43920
rect 209314 43908 209320 43920
rect 208820 43880 209320 43908
rect 208820 43868 208826 43880
rect 209314 43868 209320 43880
rect 209372 43868 209378 43920
rect 174630 43800 174636 43852
rect 174688 43840 174694 43852
rect 174688 43812 183554 43840
rect 174688 43800 174694 43812
rect 183186 43772 183192 43784
rect 173866 43744 183192 43772
rect 157334 43528 157340 43580
rect 157392 43568 157398 43580
rect 173866 43568 173894 43744
rect 183186 43732 183192 43744
rect 183244 43732 183250 43784
rect 183526 43704 183554 43812
rect 184106 43704 184112 43716
rect 183526 43676 184112 43704
rect 184106 43664 184112 43676
rect 184164 43664 184170 43716
rect 190362 43664 190368 43716
rect 190420 43704 190426 43716
rect 190420 43676 195974 43704
rect 190420 43664 190426 43676
rect 190178 43596 190184 43648
rect 190236 43636 190242 43648
rect 195946 43636 195974 43676
rect 235994 43636 236000 43648
rect 190236 43608 194364 43636
rect 195946 43608 236000 43636
rect 190236 43596 190242 43608
rect 157392 43540 173894 43568
rect 157392 43528 157398 43540
rect 189902 43528 189908 43580
rect 189960 43568 189966 43580
rect 194336 43568 194364 43608
rect 235994 43596 236000 43608
rect 236052 43596 236058 43648
rect 240134 43568 240140 43580
rect 189960 43540 194272 43568
rect 194336 43540 240140 43568
rect 189960 43528 189966 43540
rect 136542 43460 136548 43512
rect 136600 43500 136606 43512
rect 140130 43500 140136 43512
rect 136600 43472 140136 43500
rect 136600 43460 136606 43472
rect 140130 43460 140136 43472
rect 140188 43460 140194 43512
rect 151814 43460 151820 43512
rect 151872 43500 151878 43512
rect 174814 43500 174820 43512
rect 151872 43472 174820 43500
rect 151872 43460 151878 43472
rect 174814 43460 174820 43472
rect 174872 43460 174878 43512
rect 176746 43460 176752 43512
rect 176804 43500 176810 43512
rect 184566 43500 184572 43512
rect 176804 43472 184572 43500
rect 176804 43460 176810 43472
rect 184566 43460 184572 43472
rect 184624 43460 184630 43512
rect 191374 43460 191380 43512
rect 191432 43500 191438 43512
rect 194244 43500 194272 43540
rect 240134 43528 240140 43540
rect 240192 43528 240198 43580
rect 242986 43500 242992 43512
rect 191432 43472 194180 43500
rect 194244 43472 242992 43500
rect 191432 43460 191438 43472
rect 136634 43392 136640 43444
rect 136692 43432 136698 43444
rect 180886 43432 180892 43444
rect 136692 43404 180892 43432
rect 136692 43392 136698 43404
rect 180886 43392 180892 43404
rect 180944 43392 180950 43444
rect 194152 43432 194180 43472
rect 242986 43460 242992 43472
rect 243044 43460 243050 43512
rect 258074 43432 258080 43444
rect 194152 43404 258080 43432
rect 258074 43392 258080 43404
rect 258132 43392 258138 43444
rect 197078 43324 197084 43376
rect 197136 43364 197142 43376
rect 197538 43364 197544 43376
rect 197136 43336 197544 43364
rect 197136 43324 197142 43336
rect 197538 43324 197544 43336
rect 197596 43324 197602 43376
rect 201402 43324 201408 43376
rect 201460 43364 201466 43376
rect 201770 43364 201776 43376
rect 201460 43336 201776 43364
rect 201460 43324 201466 43336
rect 201770 43324 201776 43336
rect 201828 43324 201834 43376
rect 211062 43324 211068 43376
rect 211120 43364 211126 43376
rect 211522 43364 211528 43376
rect 211120 43336 211528 43364
rect 211120 43324 211126 43336
rect 211522 43324 211528 43336
rect 211580 43324 211586 43376
rect 160922 43256 160928 43308
rect 160980 43296 160986 43308
rect 161290 43296 161296 43308
rect 160980 43268 161296 43296
rect 160980 43256 160986 43268
rect 161290 43256 161296 43268
rect 161348 43256 161354 43308
rect 192018 42984 192024 43036
rect 192076 43024 192082 43036
rect 192294 43024 192300 43036
rect 192076 42996 192300 43024
rect 192076 42984 192082 42996
rect 192294 42984 192300 42996
rect 192352 42984 192358 43036
rect 212994 42984 213000 43036
rect 213052 43024 213058 43036
rect 213822 43024 213828 43036
rect 213052 42996 213828 43024
rect 213052 42984 213058 42996
rect 213822 42984 213828 42996
rect 213880 42984 213886 43036
rect 163314 42848 163320 42900
rect 163372 42888 163378 42900
rect 163958 42888 163964 42900
rect 163372 42860 163964 42888
rect 163372 42848 163378 42860
rect 163958 42848 163964 42860
rect 164016 42848 164022 42900
rect 192294 42848 192300 42900
rect 192352 42888 192358 42900
rect 192662 42888 192668 42900
rect 192352 42860 192668 42888
rect 192352 42848 192358 42860
rect 192662 42848 192668 42860
rect 192720 42848 192726 42900
rect 186038 42780 186044 42832
rect 186096 42820 186102 42832
rect 189902 42820 189908 42832
rect 186096 42792 189908 42820
rect 186096 42780 186102 42792
rect 189902 42780 189908 42792
rect 189960 42780 189966 42832
rect 165982 42576 165988 42628
rect 166040 42616 166046 42628
rect 166258 42616 166264 42628
rect 166040 42588 166264 42616
rect 166040 42576 166046 42588
rect 166258 42576 166264 42588
rect 166316 42576 166322 42628
rect 165890 42440 165896 42492
rect 165948 42480 165954 42492
rect 166810 42480 166816 42492
rect 165948 42452 166816 42480
rect 165948 42440 165954 42452
rect 166810 42440 166816 42452
rect 166868 42440 166874 42492
rect 170490 42032 170496 42084
rect 170548 42072 170554 42084
rect 580902 42072 580908 42084
rect 170548 42044 580908 42072
rect 170548 42032 170554 42044
rect 580902 42032 580908 42044
rect 580960 42032 580966 42084
rect 170582 41964 170588 42016
rect 170640 42004 170646 42016
rect 580718 42004 580724 42016
rect 170640 41976 580724 42004
rect 170640 41964 170646 41976
rect 580718 41964 580724 41976
rect 580776 41964 580782 42016
rect 171686 41896 171692 41948
rect 171744 41936 171750 41948
rect 580442 41936 580448 41948
rect 171744 41908 580448 41936
rect 171744 41896 171750 41908
rect 580442 41896 580448 41908
rect 580500 41896 580506 41948
rect 173802 41828 173808 41880
rect 173860 41868 173866 41880
rect 580534 41868 580540 41880
rect 173860 41840 580540 41868
rect 173860 41828 173866 41840
rect 580534 41828 580540 41840
rect 580592 41828 580598 41880
rect 166258 41624 166264 41676
rect 166316 41664 166322 41676
rect 166626 41664 166632 41676
rect 166316 41636 166632 41664
rect 166316 41624 166322 41636
rect 166626 41624 166632 41636
rect 166684 41624 166690 41676
rect 172514 41420 172520 41472
rect 172572 41460 172578 41472
rect 173342 41460 173348 41472
rect 172572 41432 173348 41460
rect 172572 41420 172578 41432
rect 173342 41420 173348 41432
rect 173400 41420 173406 41472
rect 170306 41352 170312 41404
rect 170364 41392 170370 41404
rect 580166 41392 580172 41404
rect 170364 41364 580172 41392
rect 170364 41352 170370 41364
rect 580166 41352 580172 41364
rect 580224 41352 580230 41404
rect 136082 41284 136088 41336
rect 136140 41324 136146 41336
rect 138842 41324 138848 41336
rect 136140 41296 138848 41324
rect 136140 41284 136146 41296
rect 138842 41284 138848 41296
rect 138900 41284 138906 41336
rect 171594 41284 171600 41336
rect 171652 41324 171658 41336
rect 580350 41324 580356 41336
rect 171652 41296 580356 41324
rect 171652 41284 171658 41296
rect 580350 41284 580356 41296
rect 580408 41284 580414 41336
rect 171502 41216 171508 41268
rect 171560 41256 171566 41268
rect 580258 41256 580264 41268
rect 171560 41228 580264 41256
rect 171560 41216 171566 41228
rect 580258 41216 580264 41228
rect 580316 41216 580322 41268
rect 172146 41148 172152 41200
rect 172204 41188 172210 41200
rect 580810 41188 580816 41200
rect 172204 41160 580816 41188
rect 172204 41148 172210 41160
rect 580810 41148 580816 41160
rect 580868 41148 580874 41200
rect 170398 41080 170404 41132
rect 170456 41120 170462 41132
rect 550174 41120 550180 41132
rect 170456 41092 550180 41120
rect 170456 41080 170462 41092
rect 550174 41080 550180 41092
rect 550232 41080 550238 41132
rect 171686 41012 171692 41064
rect 171744 41052 171750 41064
rect 551462 41052 551468 41064
rect 171744 41024 551468 41052
rect 171744 41012 171750 41024
rect 551462 41012 551468 41024
rect 551520 41012 551526 41064
rect 193950 40808 193956 40860
rect 194008 40848 194014 40860
rect 287054 40848 287060 40860
rect 194008 40820 287060 40848
rect 194008 40808 194014 40820
rect 287054 40808 287060 40820
rect 287112 40808 287118 40860
rect 198182 40740 198188 40792
rect 198240 40780 198246 40792
rect 350534 40780 350540 40792
rect 198240 40752 350540 40780
rect 198240 40740 198246 40752
rect 350534 40740 350540 40752
rect 350592 40740 350598 40792
rect 200942 40672 200948 40724
rect 201000 40712 201006 40724
rect 382274 40712 382280 40724
rect 201000 40684 382280 40712
rect 201000 40672 201006 40684
rect 382274 40672 382280 40684
rect 382332 40672 382338 40724
rect 170030 39992 170036 40044
rect 170088 40032 170094 40044
rect 580074 40032 580080 40044
rect 170088 40004 580080 40032
rect 170088 39992 170094 40004
rect 580074 39992 580080 40004
rect 580132 39992 580138 40044
rect 170214 39924 170220 39976
rect 170272 39964 170278 39976
rect 551738 39964 551744 39976
rect 170272 39936 551744 39964
rect 170272 39924 170278 39936
rect 551738 39924 551744 39936
rect 551796 39924 551802 39976
rect 170122 39856 170128 39908
rect 170180 39896 170186 39908
rect 551646 39896 551652 39908
rect 170180 39868 551652 39896
rect 170180 39856 170186 39868
rect 551646 39856 551652 39868
rect 551704 39856 551710 39908
rect 171226 39788 171232 39840
rect 171284 39828 171290 39840
rect 551554 39828 551560 39840
rect 171284 39800 551560 39828
rect 171284 39788 171290 39800
rect 551554 39788 551560 39800
rect 551612 39788 551618 39840
rect 171318 39720 171324 39772
rect 171376 39760 171382 39772
rect 551278 39760 551284 39772
rect 171376 39732 551284 39760
rect 171376 39720 171382 39732
rect 551278 39720 551284 39732
rect 551336 39720 551342 39772
rect 171410 39652 171416 39704
rect 171468 39692 171474 39704
rect 551370 39692 551376 39704
rect 171468 39664 551376 39692
rect 171468 39652 171474 39664
rect 551370 39652 551376 39664
rect 551428 39652 551434 39704
rect 198090 39516 198096 39568
rect 198148 39556 198154 39568
rect 347774 39556 347780 39568
rect 198148 39528 347780 39556
rect 198148 39516 198154 39528
rect 347774 39516 347780 39528
rect 347832 39516 347838 39568
rect 199470 39448 199476 39500
rect 199528 39488 199534 39500
rect 357434 39488 357440 39500
rect 199528 39460 357440 39488
rect 199528 39448 199534 39460
rect 357434 39448 357440 39460
rect 357492 39448 357498 39500
rect 203702 39380 203708 39432
rect 203760 39420 203766 39432
rect 365714 39420 365720 39432
rect 203760 39392 365720 39420
rect 203760 39380 203766 39392
rect 365714 39380 365720 39392
rect 365772 39380 365778 39432
rect 199378 39312 199384 39364
rect 199436 39352 199442 39364
rect 361574 39352 361580 39364
rect 199436 39324 361580 39352
rect 199436 39312 199442 39324
rect 361574 39312 361580 39324
rect 361632 39312 361638 39364
rect 172514 38564 172520 38616
rect 172572 38604 172578 38616
rect 574738 38604 574744 38616
rect 172572 38576 574744 38604
rect 172572 38564 172578 38576
rect 574738 38564 574744 38576
rect 574796 38564 574802 38616
rect 172606 38496 172612 38548
rect 172664 38536 172670 38548
rect 573358 38536 573364 38548
rect 172664 38508 573364 38536
rect 172664 38496 172670 38508
rect 573358 38496 573364 38508
rect 573416 38496 573422 38548
rect 196802 38292 196808 38344
rect 196860 38332 196866 38344
rect 332594 38332 332600 38344
rect 196860 38304 332600 38332
rect 196860 38292 196866 38304
rect 332594 38292 332600 38304
rect 332652 38292 332658 38344
rect 202138 38224 202144 38276
rect 202196 38264 202202 38276
rect 400214 38264 400220 38276
rect 202196 38236 400220 38264
rect 202196 38224 202202 38236
rect 400214 38224 400220 38236
rect 400272 38224 400278 38276
rect 209222 38156 209228 38208
rect 209280 38196 209286 38208
rect 462958 38196 462964 38208
rect 209280 38168 462964 38196
rect 209280 38156 209286 38168
rect 462958 38156 462964 38168
rect 463016 38156 463022 38208
rect 207658 38088 207664 38140
rect 207716 38128 207722 38140
rect 474734 38128 474740 38140
rect 207716 38100 474740 38128
rect 207716 38088 207722 38100
rect 474734 38088 474740 38100
rect 474792 38088 474798 38140
rect 136542 38020 136548 38072
rect 136600 38060 136606 38072
rect 144270 38060 144276 38072
rect 136600 38032 144276 38060
rect 136600 38020 136606 38032
rect 144270 38020 144276 38032
rect 144328 38020 144334 38072
rect 210602 38020 210608 38072
rect 210660 38060 210666 38072
rect 505094 38060 505100 38072
rect 210660 38032 505100 38060
rect 210660 38020 210666 38032
rect 505094 38020 505100 38032
rect 505152 38020 505158 38072
rect 210510 37952 210516 38004
rect 210568 37992 210574 38004
rect 507854 37992 507860 38004
rect 210568 37964 507860 37992
rect 210568 37952 210574 37964
rect 507854 37952 507860 37964
rect 507912 37952 507918 38004
rect 140774 37884 140780 37936
rect 140832 37924 140838 37936
rect 181346 37924 181352 37936
rect 140832 37896 181352 37924
rect 140832 37884 140838 37896
rect 181346 37884 181352 37896
rect 181404 37884 181410 37936
rect 213362 37884 213368 37936
rect 213420 37924 213426 37936
rect 539594 37924 539600 37936
rect 213420 37896 539600 37924
rect 213420 37884 213426 37896
rect 539594 37884 539600 37896
rect 539652 37884 539658 37936
rect 200850 37068 200856 37120
rect 200908 37108 200914 37120
rect 385034 37108 385040 37120
rect 200908 37080 385040 37108
rect 200908 37068 200914 37080
rect 385034 37068 385040 37080
rect 385092 37068 385098 37120
rect 211982 37000 211988 37052
rect 212040 37040 212046 37052
rect 450538 37040 450544 37052
rect 212040 37012 450544 37040
rect 212040 37000 212046 37012
rect 450538 37000 450544 37012
rect 450596 37000 450602 37052
rect 211890 36932 211896 36984
rect 211948 36972 211954 36984
rect 479518 36972 479524 36984
rect 211948 36944 479524 36972
rect 211948 36932 211954 36944
rect 479518 36932 479524 36944
rect 479576 36932 479582 36984
rect 213270 36864 213276 36916
rect 213328 36904 213334 36916
rect 543734 36904 543740 36916
rect 213328 36876 543740 36904
rect 213328 36864 213334 36876
rect 543734 36864 543740 36876
rect 543792 36864 543798 36916
rect 213178 36796 213184 36848
rect 213236 36836 213242 36848
rect 547874 36836 547880 36848
rect 213236 36808 547880 36836
rect 213236 36796 213242 36808
rect 547874 36796 547880 36808
rect 547932 36796 547938 36848
rect 216030 36728 216036 36780
rect 216088 36768 216094 36780
rect 554774 36768 554780 36780
rect 216088 36740 554780 36768
rect 216088 36728 216094 36740
rect 554774 36728 554780 36740
rect 554832 36728 554838 36780
rect 154574 36660 154580 36712
rect 154632 36700 154638 36712
rect 182450 36700 182456 36712
rect 154632 36672 182456 36700
rect 154632 36660 154638 36672
rect 182450 36660 182456 36672
rect 182508 36660 182514 36712
rect 214742 36660 214748 36712
rect 214800 36700 214806 36712
rect 557534 36700 557540 36712
rect 214800 36672 557540 36700
rect 214800 36660 214806 36672
rect 557534 36660 557540 36672
rect 557592 36660 557598 36712
rect 169938 36592 169944 36644
rect 169996 36632 170002 36644
rect 580350 36632 580356 36644
rect 169996 36604 580356 36632
rect 169996 36592 170002 36604
rect 580350 36592 580356 36604
rect 580408 36592 580414 36644
rect 169754 36524 169760 36576
rect 169812 36564 169818 36576
rect 580258 36564 580264 36576
rect 169812 36536 580264 36564
rect 169812 36524 169818 36536
rect 580258 36524 580264 36536
rect 580316 36524 580322 36576
rect 136542 35844 136548 35896
rect 136600 35884 136606 35896
rect 147030 35884 147036 35896
rect 136600 35856 147036 35884
rect 136600 35844 136606 35856
rect 147030 35844 147036 35856
rect 147088 35844 147094 35896
rect 193858 35436 193864 35488
rect 193916 35476 193922 35488
rect 298094 35476 298100 35488
rect 193916 35448 298100 35476
rect 193916 35436 193922 35448
rect 298094 35436 298100 35448
rect 298152 35436 298158 35488
rect 199286 35368 199292 35420
rect 199344 35408 199350 35420
rect 364334 35408 364340 35420
rect 199344 35380 364340 35408
rect 199344 35368 199350 35380
rect 364334 35368 364340 35380
rect 364392 35368 364398 35420
rect 209038 35300 209044 35352
rect 209096 35340 209102 35352
rect 489914 35340 489920 35352
rect 209096 35312 489920 35340
rect 209096 35300 209102 35312
rect 489914 35300 489920 35312
rect 489972 35300 489978 35352
rect 209130 35232 209136 35284
rect 209188 35272 209194 35284
rect 494054 35272 494060 35284
rect 209188 35244 494060 35272
rect 209188 35232 209194 35244
rect 494054 35232 494060 35244
rect 494112 35232 494118 35284
rect 138014 35164 138020 35216
rect 138072 35204 138078 35216
rect 181714 35204 181720 35216
rect 138072 35176 181720 35204
rect 138072 35164 138078 35176
rect 181714 35164 181720 35176
rect 181772 35164 181778 35216
rect 214650 35164 214656 35216
rect 214708 35204 214714 35216
rect 561674 35204 561680 35216
rect 214708 35176 561680 35204
rect 214708 35164 214714 35176
rect 561674 35164 561680 35176
rect 561732 35164 561738 35216
rect 199562 33872 199568 33924
rect 199620 33912 199626 33924
rect 324314 33912 324320 33924
rect 199620 33884 324320 33912
rect 199620 33872 199626 33884
rect 324314 33872 324320 33884
rect 324372 33872 324378 33924
rect 196710 33804 196716 33856
rect 196768 33844 196774 33856
rect 324406 33844 324412 33856
rect 196768 33816 324412 33844
rect 196768 33804 196774 33816
rect 324406 33804 324412 33816
rect 324464 33804 324470 33856
rect 169754 33736 169760 33788
rect 169812 33776 169818 33788
rect 184474 33776 184480 33788
rect 169812 33748 184480 33776
rect 169812 33736 169818 33748
rect 184474 33736 184480 33748
rect 184532 33736 184538 33788
rect 214558 33736 214564 33788
rect 214616 33776 214622 33788
rect 564434 33776 564440 33788
rect 214616 33748 564440 33776
rect 214616 33736 214622 33748
rect 564434 33736 564440 33748
rect 564492 33736 564498 33788
rect 136542 32988 136548 33040
rect 136600 33028 136606 33040
rect 141510 33028 141516 33040
rect 136600 33000 141516 33028
rect 136600 32988 136606 33000
rect 141510 32988 141516 33000
rect 141568 32988 141574 33040
rect 205266 32512 205272 32564
rect 205324 32552 205330 32564
rect 372614 32552 372620 32564
rect 205324 32524 372620 32552
rect 205324 32512 205330 32524
rect 372614 32512 372620 32524
rect 372672 32512 372678 32564
rect 210418 32444 210424 32496
rect 210476 32484 210482 32496
rect 511994 32484 512000 32496
rect 210476 32456 512000 32484
rect 210476 32444 210482 32456
rect 511994 32444 512000 32456
rect 512052 32444 512058 32496
rect 188246 32376 188252 32428
rect 188304 32416 188310 32428
rect 213178 32416 213184 32428
rect 188304 32388 213184 32416
rect 188304 32376 188310 32388
rect 213178 32376 213184 32388
rect 213236 32376 213242 32428
rect 215846 32376 215852 32428
rect 215904 32416 215910 32428
rect 576854 32416 576860 32428
rect 215904 32388 576860 32416
rect 215904 32376 215910 32388
rect 576854 32376 576860 32388
rect 576912 32376 576918 32428
rect 195422 31288 195428 31340
rect 195480 31328 195486 31340
rect 311894 31328 311900 31340
rect 195480 31300 311900 31328
rect 195480 31288 195486 31300
rect 311894 31288 311900 31300
rect 311952 31288 311958 31340
rect 196618 31220 196624 31272
rect 196676 31260 196682 31272
rect 331214 31260 331220 31272
rect 196676 31232 331220 31260
rect 196676 31220 196682 31232
rect 331214 31220 331220 31232
rect 331272 31220 331278 31272
rect 207934 31152 207940 31204
rect 207992 31192 207998 31204
rect 425054 31192 425060 31204
rect 207992 31164 425060 31192
rect 207992 31152 207998 31164
rect 425054 31152 425060 31164
rect 425112 31152 425118 31204
rect 214466 31084 214472 31136
rect 214524 31124 214530 31136
rect 487798 31124 487804 31136
rect 214524 31096 487804 31124
rect 214524 31084 214530 31096
rect 487798 31084 487804 31096
rect 487856 31084 487862 31136
rect 211798 31016 211804 31068
rect 211856 31056 211862 31068
rect 529934 31056 529940 31068
rect 211856 31028 529940 31056
rect 211856 31016 211862 31028
rect 529934 31016 529940 31028
rect 529992 31016 529998 31068
rect 195330 29928 195336 29980
rect 195388 29968 195394 29980
rect 313274 29968 313280 29980
rect 195388 29940 313280 29968
rect 195388 29928 195394 29940
rect 313274 29928 313280 29940
rect 313332 29928 313338 29980
rect 197998 29860 198004 29912
rect 198056 29900 198062 29912
rect 340874 29900 340880 29912
rect 198056 29872 340880 29900
rect 198056 29860 198062 29872
rect 340874 29860 340880 29872
rect 340932 29860 340938 29912
rect 202046 29792 202052 29844
rect 202104 29832 202110 29844
rect 394694 29832 394700 29844
rect 202104 29804 394700 29832
rect 202104 29792 202110 29804
rect 394694 29792 394700 29804
rect 394752 29792 394758 29844
rect 213086 29724 213092 29776
rect 213144 29764 213150 29776
rect 538214 29764 538220 29776
rect 213144 29736 538220 29764
rect 213144 29724 213150 29736
rect 538214 29724 538220 29736
rect 538272 29724 538278 29776
rect 215754 29656 215760 29708
rect 215812 29696 215818 29708
rect 572714 29696 572720 29708
rect 215812 29668 572720 29696
rect 215812 29656 215818 29668
rect 572714 29656 572720 29668
rect 572772 29656 572778 29708
rect 179414 29588 179420 29640
rect 179472 29628 179478 29640
rect 579614 29628 579620 29640
rect 179472 29600 579620 29628
rect 179472 29588 179478 29600
rect 579614 29588 579620 29600
rect 579672 29588 579678 29640
rect 135438 29044 135444 29096
rect 135496 29084 135502 29096
rect 142982 29084 142988 29096
rect 135496 29056 142988 29084
rect 135496 29044 135502 29056
rect 142982 29044 142988 29056
rect 143040 29044 143046 29096
rect 192478 28568 192484 28620
rect 192536 28608 192542 28620
rect 281534 28608 281540 28620
rect 192536 28580 281540 28608
rect 192536 28568 192542 28580
rect 281534 28568 281540 28580
rect 281592 28568 281598 28620
rect 195238 28500 195244 28552
rect 195296 28540 195302 28552
rect 307754 28540 307760 28552
rect 195296 28512 307760 28540
rect 195296 28500 195302 28512
rect 307754 28500 307760 28512
rect 307812 28500 307818 28552
rect 195146 28432 195152 28484
rect 195204 28472 195210 28484
rect 309134 28472 309140 28484
rect 195204 28444 309140 28472
rect 195204 28432 195210 28444
rect 309134 28432 309140 28444
rect 309192 28432 309198 28484
rect 199194 28364 199200 28416
rect 199252 28404 199258 28416
rect 358814 28404 358820 28416
rect 199252 28376 358820 28404
rect 199252 28364 199258 28376
rect 358814 28364 358820 28376
rect 358872 28364 358878 28416
rect 200758 28296 200764 28348
rect 200816 28336 200822 28348
rect 386414 28336 386420 28348
rect 200816 28308 386420 28336
rect 200816 28296 200822 28308
rect 386414 28296 386420 28308
rect 386472 28296 386478 28348
rect 136542 28228 136548 28280
rect 136600 28268 136606 28280
rect 148410 28268 148416 28280
rect 136600 28240 148416 28268
rect 136600 28228 136606 28240
rect 148410 28228 148416 28240
rect 148468 28228 148474 28280
rect 214374 28228 214380 28280
rect 214432 28268 214438 28280
rect 558914 28268 558920 28280
rect 214432 28240 558920 28268
rect 214432 28228 214438 28240
rect 558914 28228 558920 28240
rect 558972 28228 558978 28280
rect 193766 27208 193772 27260
rect 193824 27248 193830 27260
rect 292666 27248 292672 27260
rect 193824 27220 292672 27248
rect 193824 27208 193830 27220
rect 292666 27208 292672 27220
rect 292724 27208 292730 27260
rect 197906 27140 197912 27192
rect 197964 27180 197970 27192
rect 345014 27180 345020 27192
rect 197964 27152 345020 27180
rect 197964 27140 197970 27152
rect 345014 27140 345020 27152
rect 345072 27140 345078 27192
rect 200666 27072 200672 27124
rect 200724 27112 200730 27124
rect 378134 27112 378140 27124
rect 200724 27084 378140 27112
rect 200724 27072 200730 27084
rect 378134 27072 378140 27084
rect 378192 27072 378198 27124
rect 203334 27004 203340 27056
rect 203392 27044 203398 27056
rect 415394 27044 415400 27056
rect 203392 27016 415400 27044
rect 203392 27004 203398 27016
rect 415394 27004 415400 27016
rect 415452 27004 415458 27056
rect 151906 26936 151912 26988
rect 151964 26976 151970 26988
rect 183002 26976 183008 26988
rect 151964 26948 183008 26976
rect 151964 26936 151970 26948
rect 183002 26936 183008 26948
rect 183060 26936 183066 26988
rect 214282 26936 214288 26988
rect 214340 26976 214346 26988
rect 560294 26976 560300 26988
rect 214340 26948 560300 26976
rect 214340 26936 214346 26948
rect 560294 26936 560300 26948
rect 560352 26936 560358 26988
rect 135254 26868 135260 26920
rect 135312 26908 135318 26920
rect 181530 26908 181536 26920
rect 135312 26880 181536 26908
rect 135312 26868 135318 26880
rect 181530 26868 181536 26880
rect 181588 26868 181594 26920
rect 215662 26868 215668 26920
rect 215720 26908 215726 26920
rect 572806 26908 572812 26920
rect 215720 26880 572812 26908
rect 215720 26868 215726 26880
rect 572806 26868 572812 26880
rect 572864 26868 572870 26920
rect 3418 25712 3424 25764
rect 3476 25752 3482 25764
rect 179874 25752 179880 25764
rect 3476 25724 179880 25752
rect 3476 25712 3482 25724
rect 179874 25712 179880 25724
rect 179932 25712 179938 25764
rect 196526 25712 196532 25764
rect 196584 25752 196590 25764
rect 333974 25752 333980 25764
rect 196584 25724 333980 25752
rect 196584 25712 196590 25724
rect 333974 25712 333980 25724
rect 334032 25712 334038 25764
rect 3510 25644 3516 25696
rect 3568 25684 3574 25696
rect 179782 25684 179788 25696
rect 3568 25656 179788 25684
rect 3568 25644 3574 25656
rect 179782 25644 179788 25656
rect 179840 25644 179846 25696
rect 185394 25644 185400 25696
rect 185452 25684 185458 25696
rect 186774 25684 186780 25696
rect 185452 25656 186780 25684
rect 185452 25644 185458 25656
rect 186774 25644 186780 25656
rect 186832 25644 186838 25696
rect 199102 25644 199108 25696
rect 199160 25684 199166 25696
rect 368474 25684 368480 25696
rect 199160 25656 368480 25684
rect 199160 25644 199166 25656
rect 368474 25644 368480 25656
rect 368532 25644 368538 25696
rect 3786 25576 3792 25628
rect 3844 25616 3850 25628
rect 179690 25616 179696 25628
rect 3844 25588 179696 25616
rect 3844 25576 3850 25588
rect 179690 25576 179696 25588
rect 179748 25576 179754 25628
rect 200574 25576 200580 25628
rect 200632 25616 200638 25628
rect 383654 25616 383660 25628
rect 200632 25588 383660 25616
rect 200632 25576 200638 25588
rect 383654 25576 383660 25588
rect 383712 25576 383718 25628
rect 3694 25508 3700 25560
rect 3752 25548 3758 25560
rect 179230 25548 179236 25560
rect 3752 25520 179236 25548
rect 3752 25508 3758 25520
rect 179230 25508 179236 25520
rect 179288 25508 179294 25560
rect 212994 25508 213000 25560
rect 213052 25548 213058 25560
rect 545114 25548 545120 25560
rect 213052 25520 545120 25548
rect 213052 25508 213058 25520
rect 545114 25508 545120 25520
rect 545172 25508 545178 25560
rect 3602 25440 3608 25492
rect 3660 25480 3666 25492
rect 179138 25480 179144 25492
rect 3660 25452 179144 25480
rect 3660 25440 3666 25452
rect 179138 25440 179144 25452
rect 179196 25440 179202 25492
rect 24118 25372 24124 25424
rect 24176 25412 24182 25424
rect 179966 25412 179972 25424
rect 24176 25384 179972 25412
rect 24176 25372 24182 25384
rect 179966 25372 179972 25384
rect 180024 25372 180030 25424
rect 89714 24760 89720 24812
rect 89772 24800 89778 24812
rect 157794 24800 157800 24812
rect 89772 24772 157800 24800
rect 89772 24760 89778 24772
rect 157794 24760 157800 24772
rect 157852 24760 157858 24812
rect 95234 24692 95240 24744
rect 95292 24732 95298 24744
rect 168282 24732 168288 24744
rect 95292 24704 168288 24732
rect 95292 24692 95298 24704
rect 168282 24692 168288 24704
rect 168340 24692 168346 24744
rect 81434 24624 81440 24676
rect 81492 24664 81498 24676
rect 166902 24664 166908 24676
rect 81492 24636 166908 24664
rect 81492 24624 81498 24636
rect 166902 24624 166908 24636
rect 166960 24624 166966 24676
rect 71774 24556 71780 24608
rect 71832 24596 71838 24608
rect 157610 24596 157616 24608
rect 71832 24568 157616 24596
rect 71832 24556 71838 24568
rect 157610 24556 157616 24568
rect 157668 24556 157674 24608
rect 64874 24488 64880 24540
rect 64932 24528 64938 24540
rect 165246 24528 165252 24540
rect 64932 24500 165252 24528
rect 64932 24488 64938 24500
rect 165246 24488 165252 24500
rect 165304 24488 165310 24540
rect 60734 24420 60740 24472
rect 60792 24460 60798 24472
rect 164970 24460 164976 24472
rect 60792 24432 164976 24460
rect 60792 24420 60798 24432
rect 164970 24420 164976 24432
rect 165028 24420 165034 24472
rect 195054 24420 195060 24472
rect 195112 24460 195118 24472
rect 316034 24460 316040 24472
rect 195112 24432 316040 24460
rect 195112 24420 195118 24432
rect 316034 24420 316040 24432
rect 316092 24420 316098 24472
rect 57974 24352 57980 24404
rect 58032 24392 58038 24404
rect 163590 24392 163596 24404
rect 58032 24364 163596 24392
rect 58032 24352 58038 24364
rect 163590 24352 163596 24364
rect 163648 24352 163654 24404
rect 199010 24352 199016 24404
rect 199068 24392 199074 24404
rect 362954 24392 362960 24404
rect 199068 24364 362960 24392
rect 199068 24352 199074 24364
rect 362954 24352 362960 24364
rect 363012 24352 363018 24404
rect 46934 24284 46940 24336
rect 46992 24324 46998 24336
rect 158622 24324 158628 24336
rect 46992 24296 158628 24324
rect 46992 24284 46998 24296
rect 158622 24284 158628 24296
rect 158680 24284 158686 24336
rect 200482 24284 200488 24336
rect 200540 24324 200546 24336
rect 382366 24324 382372 24336
rect 200540 24296 382372 24324
rect 200540 24284 200546 24296
rect 382366 24284 382372 24296
rect 382424 24284 382430 24336
rect 45554 24216 45560 24268
rect 45612 24256 45618 24268
rect 159634 24256 159640 24268
rect 45612 24228 159640 24256
rect 45612 24216 45618 24228
rect 159634 24216 159640 24228
rect 159692 24216 159698 24268
rect 208946 24216 208952 24268
rect 209004 24256 209010 24268
rect 488534 24256 488540 24268
rect 209004 24228 488540 24256
rect 209004 24216 209010 24228
rect 488534 24216 488540 24228
rect 488592 24216 488598 24268
rect 38654 24148 38660 24200
rect 38712 24188 38718 24200
rect 159726 24188 159732 24200
rect 38712 24160 159732 24188
rect 38712 24148 38718 24160
rect 159726 24148 159732 24160
rect 159784 24148 159790 24200
rect 214098 24148 214104 24200
rect 214156 24188 214162 24200
rect 556246 24188 556252 24200
rect 214156 24160 556252 24188
rect 214156 24148 214162 24160
rect 556246 24148 556252 24160
rect 556304 24148 556310 24200
rect 35894 24080 35900 24132
rect 35952 24120 35958 24132
rect 162578 24120 162584 24132
rect 35952 24092 162584 24120
rect 35952 24080 35958 24092
rect 162578 24080 162584 24092
rect 162636 24080 162642 24132
rect 214190 24080 214196 24132
rect 214248 24120 214254 24132
rect 563054 24120 563060 24132
rect 214248 24092 563060 24120
rect 214248 24080 214254 24092
rect 563054 24080 563060 24092
rect 563112 24080 563118 24132
rect 107654 24012 107660 24064
rect 107712 24052 107718 24064
rect 158530 24052 158536 24064
rect 107712 24024 158536 24052
rect 107712 24012 107718 24024
rect 158530 24012 158536 24024
rect 158588 24012 158594 24064
rect 120074 23944 120080 23996
rect 120132 23984 120138 23996
rect 169018 23984 169024 23996
rect 120132 23956 169024 23984
rect 120132 23944 120138 23956
rect 169018 23944 169024 23956
rect 169076 23944 169082 23996
rect 110414 23876 110420 23928
rect 110472 23916 110478 23928
rect 157702 23916 157708 23928
rect 110472 23888 157708 23916
rect 110472 23876 110478 23888
rect 157702 23876 157708 23888
rect 157760 23876 157766 23928
rect 193674 23332 193680 23384
rect 193732 23372 193738 23384
rect 299474 23372 299480 23384
rect 193732 23344 299480 23372
rect 193732 23332 193738 23344
rect 299474 23332 299480 23344
rect 299532 23332 299538 23384
rect 196434 23264 196440 23316
rect 196492 23304 196498 23316
rect 325694 23304 325700 23316
rect 196492 23276 325700 23304
rect 196492 23264 196498 23276
rect 325694 23264 325700 23276
rect 325752 23264 325758 23316
rect 197814 23196 197820 23248
rect 197872 23236 197878 23248
rect 349154 23236 349160 23248
rect 197872 23208 349160 23236
rect 197872 23196 197878 23208
rect 349154 23196 349160 23208
rect 349212 23196 349218 23248
rect 201862 23128 201868 23180
rect 201920 23168 201926 23180
rect 396074 23168 396080 23180
rect 201920 23140 396080 23168
rect 201920 23128 201926 23140
rect 396074 23128 396080 23140
rect 396132 23128 396138 23180
rect 201954 23060 201960 23112
rect 202012 23100 202018 23112
rect 398834 23100 398840 23112
rect 202012 23072 398840 23100
rect 202012 23060 202018 23072
rect 398834 23060 398840 23072
rect 398892 23060 398898 23112
rect 204806 22992 204812 23044
rect 204864 23032 204870 23044
rect 440326 23032 440332 23044
rect 204864 23004 440332 23032
rect 204864 22992 204870 23004
rect 440326 22992 440332 23004
rect 440384 22992 440390 23044
rect 85574 22924 85580 22976
rect 85632 22964 85638 22976
rect 166258 22964 166264 22976
rect 85632 22936 166264 22964
rect 85632 22924 85638 22936
rect 166258 22924 166264 22936
rect 166316 22924 166322 22976
rect 210234 22924 210240 22976
rect 210292 22964 210298 22976
rect 503714 22964 503720 22976
rect 210292 22936 503720 22964
rect 210292 22924 210298 22936
rect 503714 22924 503720 22936
rect 503772 22924 503778 22976
rect 31754 22856 31760 22908
rect 31812 22896 31818 22908
rect 162118 22896 162124 22908
rect 31812 22868 162124 22896
rect 31812 22856 31818 22868
rect 162118 22856 162124 22868
rect 162176 22856 162182 22908
rect 210326 22856 210332 22908
rect 210384 22896 210390 22908
rect 506474 22896 506480 22908
rect 210384 22868 506480 22896
rect 210384 22856 210390 22868
rect 506474 22856 506480 22868
rect 506532 22856 506538 22908
rect 13814 22788 13820 22840
rect 13872 22828 13878 22840
rect 160554 22828 160560 22840
rect 13872 22800 160560 22828
rect 13872 22788 13878 22800
rect 160554 22788 160560 22800
rect 160612 22788 160618 22840
rect 211706 22788 211712 22840
rect 211764 22828 211770 22840
rect 517514 22828 517520 22840
rect 211764 22800 517520 22828
rect 211764 22788 211770 22800
rect 517514 22788 517520 22800
rect 517572 22788 517578 22840
rect 9674 22720 9680 22772
rect 9732 22760 9738 22772
rect 160646 22760 160652 22772
rect 9732 22732 160652 22760
rect 9732 22720 9738 22732
rect 160646 22720 160652 22732
rect 160704 22720 160710 22772
rect 179414 22720 179420 22772
rect 179472 22760 179478 22772
rect 184382 22760 184388 22772
rect 179472 22732 184388 22760
rect 179472 22720 179478 22732
rect 184382 22720 184388 22732
rect 184440 22720 184446 22772
rect 185302 22720 185308 22772
rect 185360 22760 185366 22772
rect 193674 22760 193680 22772
rect 185360 22732 193680 22760
rect 185360 22720 185366 22732
rect 193674 22720 193680 22732
rect 193732 22720 193738 22772
rect 214006 22720 214012 22772
rect 214064 22760 214070 22772
rect 564526 22760 564532 22772
rect 214064 22732 564532 22760
rect 214064 22720 214070 22732
rect 564526 22720 564532 22732
rect 564584 22720 564590 22772
rect 121454 21700 121460 21752
rect 121512 21740 121518 21752
rect 169110 21740 169116 21752
rect 121512 21712 169116 21740
rect 121512 21700 121518 21712
rect 169110 21700 169116 21712
rect 169168 21700 169174 21752
rect 78674 21632 78680 21684
rect 78732 21672 78738 21684
rect 166166 21672 166172 21684
rect 78732 21644 166172 21672
rect 78732 21632 78738 21644
rect 166166 21632 166172 21644
rect 166224 21632 166230 21684
rect 190822 21632 190828 21684
rect 190880 21672 190886 21684
rect 260834 21672 260840 21684
rect 190880 21644 260840 21672
rect 190880 21632 190886 21644
rect 260834 21632 260840 21644
rect 260892 21632 260898 21684
rect 53834 21564 53840 21616
rect 53892 21604 53898 21616
rect 162854 21604 162860 21616
rect 53892 21576 162860 21604
rect 53892 21564 53898 21576
rect 162854 21564 162860 21576
rect 162912 21564 162918 21616
rect 258626 21564 258632 21616
rect 258684 21604 258690 21616
rect 471974 21604 471980 21616
rect 258684 21576 471980 21604
rect 258684 21564 258690 21576
rect 471974 21564 471980 21576
rect 472032 21564 472038 21616
rect 49694 21496 49700 21548
rect 49752 21536 49758 21548
rect 163406 21536 163412 21548
rect 49752 21508 163412 21536
rect 49752 21496 49758 21508
rect 163406 21496 163412 21508
rect 163464 21496 163470 21548
rect 204714 21496 204720 21548
rect 204772 21536 204778 21548
rect 441614 21536 441620 21548
rect 204772 21508 441620 21536
rect 204772 21496 204778 21508
rect 441614 21496 441620 21508
rect 441672 21496 441678 21548
rect 15194 21428 15200 21480
rect 15252 21468 15258 21480
rect 158438 21468 158444 21480
rect 15252 21440 158444 21468
rect 15252 21428 15258 21440
rect 158438 21428 158444 21440
rect 158496 21428 158502 21480
rect 211614 21428 211620 21480
rect 211672 21468 211678 21480
rect 520274 21468 520280 21480
rect 211672 21440 520280 21468
rect 211672 21428 211678 21440
rect 520274 21428 520280 21440
rect 520332 21428 520338 21480
rect 4154 21360 4160 21412
rect 4212 21400 4218 21412
rect 159542 21400 159548 21412
rect 4212 21372 159548 21400
rect 4212 21360 4218 21372
rect 159542 21360 159548 21372
rect 159600 21360 159606 21412
rect 212902 21360 212908 21412
rect 212960 21400 212966 21412
rect 540974 21400 540980 21412
rect 212960 21372 540980 21400
rect 212960 21360 212966 21372
rect 540974 21360 540980 21372
rect 541032 21360 541038 21412
rect 3418 20612 3424 20664
rect 3476 20652 3482 20664
rect 177574 20652 177580 20664
rect 3476 20624 177580 20652
rect 3476 20612 3482 20624
rect 177574 20612 177580 20624
rect 177632 20612 177638 20664
rect 190638 20544 190644 20596
rect 190696 20584 190702 20596
rect 262214 20584 262220 20596
rect 190696 20556 262220 20584
rect 190696 20544 190702 20556
rect 262214 20544 262220 20556
rect 262272 20544 262278 20596
rect 169846 20476 169852 20528
rect 169904 20516 169910 20528
rect 269758 20516 269764 20528
rect 169904 20488 269764 20516
rect 169904 20476 169910 20488
rect 269758 20476 269764 20488
rect 269816 20476 269822 20528
rect 253750 20408 253756 20460
rect 253808 20448 253814 20460
rect 411254 20448 411260 20460
rect 253808 20420 411260 20448
rect 253808 20408 253814 20420
rect 411254 20408 411260 20420
rect 411312 20408 411318 20460
rect 200390 20340 200396 20392
rect 200448 20380 200454 20392
rect 379514 20380 379520 20392
rect 200448 20352 379520 20380
rect 200448 20340 200454 20352
rect 379514 20340 379520 20352
rect 379572 20340 379578 20392
rect 259362 20272 259368 20324
rect 259420 20312 259426 20324
rect 454034 20312 454040 20324
rect 259420 20284 454040 20312
rect 259420 20272 259426 20284
rect 454034 20272 454040 20284
rect 454092 20272 454098 20324
rect 122834 20204 122840 20256
rect 122892 20244 122898 20256
rect 168926 20244 168932 20256
rect 122892 20216 168932 20244
rect 122892 20204 122898 20216
rect 168926 20204 168932 20216
rect 168984 20204 168990 20256
rect 203518 20204 203524 20256
rect 203576 20244 203582 20256
rect 404354 20244 404360 20256
rect 203576 20216 404360 20244
rect 203576 20204 203582 20216
rect 404354 20204 404360 20216
rect 404412 20204 404418 20256
rect 102134 20136 102140 20188
rect 102192 20176 102198 20188
rect 167638 20176 167644 20188
rect 102192 20148 167644 20176
rect 102192 20136 102198 20148
rect 167638 20136 167644 20148
rect 167696 20136 167702 20188
rect 205174 20136 205180 20188
rect 205232 20176 205238 20188
rect 415486 20176 415492 20188
rect 205232 20148 415492 20176
rect 205232 20136 205238 20148
rect 415486 20136 415492 20148
rect 415544 20136 415550 20188
rect 82814 20068 82820 20120
rect 82872 20108 82878 20120
rect 166074 20108 166080 20120
rect 82872 20080 166080 20108
rect 82872 20068 82878 20080
rect 166074 20068 166080 20080
rect 166132 20068 166138 20120
rect 203242 20068 203248 20120
rect 203300 20108 203306 20120
rect 422294 20108 422300 20120
rect 203300 20080 422300 20108
rect 203300 20068 203306 20080
rect 422294 20068 422300 20080
rect 422352 20068 422358 20120
rect 67634 20000 67640 20052
rect 67692 20040 67698 20052
rect 164878 20040 164884 20052
rect 67692 20012 164884 20040
rect 67692 20000 67698 20012
rect 164878 20000 164884 20012
rect 164936 20000 164942 20052
rect 204622 20000 204628 20052
rect 204680 20040 204686 20052
rect 429194 20040 429200 20052
rect 204680 20012 429200 20040
rect 204680 20000 204686 20012
rect 429194 20000 429200 20012
rect 429252 20000 429258 20052
rect 34514 19932 34520 19984
rect 34572 19972 34578 19984
rect 162026 19972 162032 19984
rect 34572 19944 162032 19972
rect 34572 19932 34578 19944
rect 162026 19932 162032 19944
rect 162084 19932 162090 19984
rect 186682 19932 186688 19984
rect 186740 19972 186746 19984
rect 203518 19972 203524 19984
rect 186740 19944 203524 19972
rect 186740 19932 186746 19944
rect 203518 19932 203524 19944
rect 203576 19932 203582 19984
rect 206278 19932 206284 19984
rect 206336 19972 206342 19984
rect 456794 19972 456800 19984
rect 206336 19944 456800 19972
rect 206336 19932 206342 19944
rect 456794 19932 456800 19944
rect 456852 19932 456858 19984
rect 192202 19184 192208 19236
rect 192260 19224 192266 19236
rect 273254 19224 273260 19236
rect 192260 19196 273260 19224
rect 192260 19184 192266 19196
rect 273254 19184 273260 19196
rect 273312 19184 273318 19236
rect 192386 19116 192392 19168
rect 192444 19156 192450 19168
rect 276014 19156 276020 19168
rect 192444 19128 276020 19156
rect 192444 19116 192450 19128
rect 276014 19116 276020 19128
rect 276072 19116 276078 19168
rect 192294 19048 192300 19100
rect 192352 19088 192358 19100
rect 280154 19088 280160 19100
rect 192352 19060 280160 19088
rect 192352 19048 192358 19060
rect 280154 19048 280160 19060
rect 280212 19048 280218 19100
rect 193582 18980 193588 19032
rect 193640 19020 193646 19032
rect 291194 19020 291200 19032
rect 193640 18992 291200 19020
rect 193640 18980 193646 18992
rect 291194 18980 291200 18992
rect 291252 18980 291258 19032
rect 193490 18912 193496 18964
rect 193548 18952 193554 18964
rect 293954 18952 293960 18964
rect 193548 18924 293960 18952
rect 193548 18912 193554 18924
rect 293954 18912 293960 18924
rect 294012 18912 294018 18964
rect 194962 18844 194968 18896
rect 195020 18884 195026 18896
rect 304994 18884 305000 18896
rect 195020 18856 305000 18884
rect 195020 18844 195026 18856
rect 304994 18844 305000 18856
rect 305052 18844 305058 18896
rect 69014 18776 69020 18828
rect 69072 18816 69078 18828
rect 164694 18816 164700 18828
rect 69072 18788 164700 18816
rect 69072 18776 69078 18788
rect 164694 18776 164700 18788
rect 164752 18776 164758 18828
rect 196342 18776 196348 18828
rect 196400 18816 196406 18828
rect 329834 18816 329840 18828
rect 196400 18788 329840 18816
rect 196400 18776 196406 18788
rect 329834 18776 329840 18788
rect 329892 18776 329898 18828
rect 69106 18708 69112 18760
rect 69164 18748 69170 18760
rect 164786 18748 164792 18760
rect 69164 18720 164792 18748
rect 69164 18708 69170 18720
rect 164786 18708 164792 18720
rect 164844 18708 164850 18760
rect 206646 18708 206652 18760
rect 206704 18748 206710 18760
rect 418154 18748 418160 18760
rect 206704 18720 418160 18748
rect 206704 18708 206710 18720
rect 418154 18708 418160 18720
rect 418212 18708 418218 18760
rect 11054 18640 11060 18692
rect 11112 18680 11118 18692
rect 160370 18680 160376 18692
rect 11112 18652 160376 18680
rect 11112 18640 11118 18652
rect 160370 18640 160376 18652
rect 160428 18640 160434 18692
rect 215938 18640 215944 18692
rect 215996 18680 216002 18692
rect 436094 18680 436100 18692
rect 215996 18652 436100 18680
rect 215996 18640 216002 18652
rect 436094 18640 436100 18652
rect 436152 18640 436158 18692
rect 6914 18572 6920 18624
rect 6972 18612 6978 18624
rect 160462 18612 160468 18624
rect 6972 18584 160468 18612
rect 6972 18572 6978 18584
rect 160462 18572 160468 18584
rect 160520 18572 160526 18624
rect 260190 18572 260196 18624
rect 260248 18612 260254 18624
rect 536834 18612 536840 18624
rect 260248 18584 536840 18612
rect 260248 18572 260254 18584
rect 536834 18572 536840 18584
rect 536892 18572 536898 18624
rect 255866 17892 255872 17944
rect 255924 17932 255930 17944
rect 397454 17932 397460 17944
rect 255924 17904 397460 17932
rect 255924 17892 255930 17904
rect 397454 17892 397460 17904
rect 397512 17892 397518 17944
rect 210142 17824 210148 17876
rect 210200 17864 210206 17876
rect 468478 17864 468484 17876
rect 210200 17836 468484 17864
rect 210200 17824 210206 17836
rect 468478 17824 468484 17836
rect 468536 17824 468542 17876
rect 207382 17756 207388 17808
rect 207440 17796 207446 17808
rect 466454 17796 466460 17808
rect 207440 17768 466460 17796
rect 207440 17756 207446 17768
rect 466454 17756 466460 17768
rect 466512 17756 466518 17808
rect 207566 17688 207572 17740
rect 207624 17728 207630 17740
rect 470594 17728 470600 17740
rect 207624 17700 470600 17728
rect 207624 17688 207630 17700
rect 470594 17688 470600 17700
rect 470652 17688 470658 17740
rect 207474 17620 207480 17672
rect 207532 17660 207538 17672
rect 473354 17660 473360 17672
rect 207532 17632 473360 17660
rect 207532 17620 207538 17632
rect 473354 17620 473360 17632
rect 473412 17620 473418 17672
rect 211430 17552 211436 17604
rect 211488 17592 211494 17604
rect 521654 17592 521660 17604
rect 211488 17564 521660 17592
rect 211488 17552 211494 17564
rect 521654 17552 521660 17564
rect 521712 17552 521718 17604
rect 126974 17484 126980 17536
rect 127032 17524 127038 17536
rect 180242 17524 180248 17536
rect 127032 17496 180248 17524
rect 127032 17484 127038 17496
rect 180242 17484 180248 17496
rect 180300 17484 180306 17536
rect 211522 17484 211528 17536
rect 211580 17524 211586 17536
rect 524414 17524 524420 17536
rect 211580 17496 524420 17524
rect 211580 17484 211586 17496
rect 524414 17484 524420 17496
rect 524472 17484 524478 17536
rect 125594 17416 125600 17468
rect 125652 17456 125658 17468
rect 179598 17456 179604 17468
rect 125652 17428 179604 17456
rect 125652 17416 125658 17428
rect 179598 17416 179604 17428
rect 179656 17416 179662 17468
rect 211338 17416 211344 17468
rect 211396 17456 211402 17468
rect 528554 17456 528560 17468
rect 211396 17428 528560 17456
rect 211396 17416 211402 17428
rect 528554 17416 528560 17428
rect 528612 17416 528618 17468
rect 60826 17348 60832 17400
rect 60884 17388 60890 17400
rect 164602 17388 164608 17400
rect 60884 17360 164608 17388
rect 60884 17348 60890 17360
rect 164602 17348 164608 17360
rect 164660 17348 164666 17400
rect 212718 17348 212724 17400
rect 212776 17388 212782 17400
rect 535454 17388 535460 17400
rect 212776 17360 535460 17388
rect 212776 17348 212782 17360
rect 535454 17348 535460 17360
rect 535512 17348 535518 17400
rect 51074 17280 51080 17332
rect 51132 17320 51138 17332
rect 163314 17320 163320 17332
rect 51132 17292 163320 17320
rect 51132 17280 51138 17292
rect 163314 17280 163320 17292
rect 163372 17280 163378 17332
rect 212626 17280 212632 17332
rect 212684 17320 212690 17332
rect 539686 17320 539692 17332
rect 212684 17292 539692 17320
rect 212684 17280 212690 17292
rect 539686 17280 539692 17292
rect 539744 17280 539750 17332
rect 33134 17212 33140 17264
rect 33192 17252 33198 17264
rect 161934 17252 161940 17264
rect 33192 17224 161940 17252
rect 33192 17212 33198 17224
rect 161934 17212 161940 17224
rect 161992 17212 161998 17264
rect 212810 17212 212816 17264
rect 212868 17252 212874 17264
rect 546494 17252 546500 17264
rect 212868 17224 546500 17252
rect 212868 17212 212874 17224
rect 546494 17212 546500 17224
rect 546552 17212 546558 17264
rect 194870 17144 194876 17196
rect 194928 17184 194934 17196
rect 316126 17184 316132 17196
rect 194928 17156 316132 17184
rect 194928 17144 194934 17156
rect 316126 17144 316132 17156
rect 316184 17144 316190 17196
rect 202966 16328 202972 16380
rect 203024 16368 203030 16380
rect 414290 16368 414296 16380
rect 203024 16340 414296 16368
rect 203024 16328 203030 16340
rect 414290 16328 414296 16340
rect 414348 16328 414354 16380
rect 203058 16260 203064 16312
rect 203116 16300 203122 16312
rect 417418 16300 417424 16312
rect 203116 16272 417424 16300
rect 203116 16260 203122 16272
rect 417418 16260 417424 16272
rect 417476 16260 417482 16312
rect 116394 16192 116400 16244
rect 116452 16232 116458 16244
rect 168834 16232 168840 16244
rect 116452 16204 168840 16232
rect 116452 16192 116458 16204
rect 168834 16192 168840 16204
rect 168892 16192 168898 16244
rect 203150 16192 203156 16244
rect 203208 16232 203214 16244
rect 420914 16232 420920 16244
rect 203208 16204 420920 16232
rect 203208 16192 203214 16204
rect 420914 16192 420920 16204
rect 420972 16192 420978 16244
rect 104066 16124 104072 16176
rect 104124 16164 104130 16176
rect 167362 16164 167368 16176
rect 104124 16136 167368 16164
rect 104124 16124 104130 16136
rect 167362 16124 167368 16136
rect 167420 16124 167426 16176
rect 204530 16124 204536 16176
rect 204588 16164 204594 16176
rect 432046 16164 432052 16176
rect 204588 16136 432052 16164
rect 204588 16124 204594 16136
rect 432046 16124 432052 16136
rect 432104 16124 432110 16176
rect 102226 16056 102232 16108
rect 102284 16096 102290 16108
rect 167454 16096 167460 16108
rect 102284 16068 167460 16096
rect 102284 16056 102290 16068
rect 167454 16056 167460 16068
rect 167512 16056 167518 16108
rect 204438 16056 204444 16108
rect 204496 16096 204502 16108
rect 435082 16096 435088 16108
rect 204496 16068 435088 16096
rect 204496 16056 204502 16068
rect 435082 16056 435088 16068
rect 435140 16056 435146 16108
rect 98178 15988 98184 16040
rect 98236 16028 98242 16040
rect 167546 16028 167552 16040
rect 98236 16000 167552 16028
rect 98236 15988 98242 16000
rect 167546 15988 167552 16000
rect 167604 15988 167610 16040
rect 204346 15988 204352 16040
rect 204404 16028 204410 16040
rect 439130 16028 439136 16040
rect 204404 16000 439136 16028
rect 204404 15988 204410 16000
rect 439130 15988 439136 16000
rect 439188 15988 439194 16040
rect 28442 15920 28448 15972
rect 28500 15960 28506 15972
rect 161842 15960 161848 15972
rect 28500 15932 161848 15960
rect 28500 15920 28506 15932
rect 161842 15920 161848 15932
rect 161900 15920 161906 15972
rect 208854 15920 208860 15972
rect 208912 15960 208918 15972
rect 490006 15960 490012 15972
rect 208912 15932 490012 15960
rect 208912 15920 208918 15932
rect 490006 15920 490012 15932
rect 490064 15920 490070 15972
rect 2866 15852 2872 15904
rect 2924 15892 2930 15904
rect 158714 15892 158720 15904
rect 2924 15864 158720 15892
rect 2924 15852 2930 15864
rect 158714 15852 158720 15864
rect 158772 15852 158778 15904
rect 189258 15852 189264 15904
rect 189316 15892 189322 15904
rect 203978 15892 203984 15904
rect 189316 15864 203984 15892
rect 189316 15852 189322 15864
rect 203978 15852 203984 15864
rect 204036 15852 204042 15904
rect 210050 15852 210056 15904
rect 210108 15892 210114 15904
rect 507210 15892 507216 15904
rect 210108 15864 507216 15892
rect 210108 15852 210114 15864
rect 507210 15852 507216 15864
rect 507268 15852 507274 15904
rect 202414 15104 202420 15156
rect 202472 15144 202478 15156
rect 339494 15144 339500 15156
rect 202472 15116 339500 15144
rect 202472 15104 202478 15116
rect 339494 15104 339500 15116
rect 339552 15104 339558 15156
rect 196158 15036 196164 15088
rect 196216 15076 196222 15088
rect 336274 15076 336280 15088
rect 196216 15048 336280 15076
rect 196216 15036 196222 15048
rect 336274 15036 336280 15048
rect 336332 15036 336338 15088
rect 197630 14968 197636 15020
rect 197688 15008 197694 15020
rect 342898 15008 342904 15020
rect 197688 14980 342904 15008
rect 197688 14968 197694 14980
rect 342898 14968 342904 14980
rect 342956 14968 342962 15020
rect 197722 14900 197728 14952
rect 197780 14940 197786 14952
rect 346946 14940 346952 14952
rect 197780 14912 346952 14940
rect 197780 14900 197786 14912
rect 346946 14900 346952 14912
rect 347004 14900 347010 14952
rect 259270 14832 259276 14884
rect 259328 14872 259334 14884
rect 447410 14872 447416 14884
rect 259328 14844 447416 14872
rect 259328 14832 259334 14844
rect 447410 14832 447416 14844
rect 447468 14832 447474 14884
rect 206186 14764 206192 14816
rect 206244 14804 206250 14816
rect 453298 14804 453304 14816
rect 206244 14776 453304 14804
rect 206244 14764 206250 14776
rect 453298 14764 453304 14776
rect 453356 14764 453362 14816
rect 206094 14696 206100 14748
rect 206152 14736 206158 14748
rect 456886 14736 456892 14748
rect 206152 14708 456892 14736
rect 206152 14696 206158 14708
rect 456886 14696 456892 14708
rect 456944 14696 456950 14748
rect 114002 14628 114008 14680
rect 114060 14668 114066 14680
rect 168742 14668 168748 14680
rect 114060 14640 168748 14668
rect 114060 14628 114066 14640
rect 168742 14628 168748 14640
rect 168800 14628 168806 14680
rect 207198 14628 207204 14680
rect 207256 14668 207262 14680
rect 469858 14668 469864 14680
rect 207256 14640 469864 14668
rect 207256 14628 207262 14640
rect 469858 14628 469864 14640
rect 469916 14628 469922 14680
rect 87506 14560 87512 14612
rect 87564 14600 87570 14612
rect 165890 14600 165896 14612
rect 87564 14572 165896 14600
rect 87564 14560 87570 14572
rect 165890 14560 165896 14572
rect 165948 14560 165954 14612
rect 207290 14560 207296 14612
rect 207348 14600 207354 14612
rect 473446 14600 473452 14612
rect 207348 14572 473452 14600
rect 207348 14560 207354 14572
rect 473446 14560 473452 14572
rect 473504 14560 473510 14612
rect 80882 14492 80888 14544
rect 80940 14532 80946 14544
rect 165982 14532 165988 14544
rect 80940 14504 165988 14532
rect 80940 14492 80946 14504
rect 165982 14492 165988 14504
rect 166040 14492 166046 14544
rect 207106 14492 207112 14544
rect 207164 14532 207170 14544
rect 476482 14532 476488 14544
rect 207164 14504 476488 14532
rect 207164 14492 207170 14504
rect 476482 14492 476488 14504
rect 476540 14492 476546 14544
rect 13538 14424 13544 14476
rect 13596 14464 13602 14476
rect 160278 14464 160284 14476
rect 13596 14436 160284 14464
rect 13596 14424 13602 14436
rect 160278 14424 160284 14436
rect 160336 14424 160342 14476
rect 212534 14424 212540 14476
rect 212592 14464 212598 14476
rect 542722 14464 542728 14476
rect 212592 14436 542728 14464
rect 212592 14424 212598 14436
rect 542722 14424 542728 14436
rect 542780 14424 542786 14476
rect 197170 14356 197176 14408
rect 197228 14396 197234 14408
rect 332686 14396 332692 14408
rect 197228 14368 332692 14396
rect 197228 14356 197234 14368
rect 332686 14356 332692 14368
rect 332744 14356 332750 14408
rect 196250 14288 196256 14340
rect 196308 14328 196314 14340
rect 328730 14328 328736 14340
rect 196308 14300 328736 14328
rect 196308 14288 196314 14300
rect 328730 14288 328736 14300
rect 328788 14288 328794 14340
rect 114738 13268 114744 13320
rect 114796 13308 114802 13320
rect 168650 13308 168656 13320
rect 114796 13280 168656 13308
rect 114796 13268 114802 13280
rect 168650 13268 168656 13280
rect 168708 13268 168714 13320
rect 192110 13268 192116 13320
rect 192168 13308 192174 13320
rect 272426 13308 272432 13320
rect 192168 13280 272432 13308
rect 192168 13268 192174 13280
rect 272426 13268 272432 13280
rect 272484 13268 272490 13320
rect 63218 13200 63224 13252
rect 63276 13240 63282 13252
rect 164510 13240 164516 13252
rect 63276 13212 164516 13240
rect 63276 13200 63282 13212
rect 164510 13200 164516 13212
rect 164568 13200 164574 13252
rect 259178 13200 259184 13252
rect 259236 13240 259242 13252
rect 465166 13240 465172 13252
rect 259236 13212 465172 13240
rect 259236 13200 259242 13212
rect 465166 13200 465172 13212
rect 465224 13200 465230 13252
rect 30098 13132 30104 13184
rect 30156 13172 30162 13184
rect 161658 13172 161664 13184
rect 30156 13144 161664 13172
rect 30156 13132 30162 13144
rect 161658 13132 161664 13144
rect 161716 13132 161722 13184
rect 209958 13132 209964 13184
rect 210016 13172 210022 13184
rect 500586 13172 500592 13184
rect 210016 13144 500592 13172
rect 210016 13132 210022 13144
rect 500586 13132 500592 13144
rect 500644 13132 500650 13184
rect 26234 13064 26240 13116
rect 26292 13104 26298 13116
rect 161750 13104 161756 13116
rect 26292 13076 161756 13104
rect 26292 13064 26298 13076
rect 161750 13064 161756 13076
rect 161808 13064 161814 13116
rect 215570 13064 215576 13116
rect 215628 13104 215634 13116
rect 578602 13104 578608 13116
rect 215628 13076 578608 13104
rect 215628 13064 215634 13076
rect 578602 13064 578608 13076
rect 578660 13064 578666 13116
rect 185210 12384 185216 12436
rect 185268 12424 185274 12436
rect 192018 12424 192024 12436
rect 185268 12396 192024 12424
rect 185268 12384 185274 12396
rect 192018 12384 192024 12396
rect 192076 12384 192082 12436
rect 253658 12384 253664 12436
rect 253716 12424 253722 12436
rect 394234 12424 394240 12436
rect 253716 12396 394240 12424
rect 253716 12384 253722 12396
rect 394234 12384 394240 12396
rect 394292 12384 394298 12436
rect 203794 12316 203800 12368
rect 203852 12356 203858 12368
rect 376018 12356 376024 12368
rect 203852 12328 376024 12356
rect 203852 12316 203858 12328
rect 376018 12316 376024 12328
rect 376076 12316 376082 12368
rect 200298 12248 200304 12300
rect 200356 12288 200362 12300
rect 389450 12288 389456 12300
rect 200356 12260 389456 12288
rect 200356 12248 200362 12260
rect 389450 12248 389456 12260
rect 389508 12248 389514 12300
rect 205910 12180 205916 12232
rect 205968 12220 205974 12232
rect 448606 12220 448612 12232
rect 205968 12192 448612 12220
rect 205968 12180 205974 12192
rect 448606 12180 448612 12192
rect 448664 12180 448670 12232
rect 206002 12112 206008 12164
rect 206060 12152 206066 12164
rect 451642 12152 451648 12164
rect 206060 12124 451648 12152
rect 206060 12112 206066 12124
rect 451642 12112 451648 12124
rect 451700 12112 451706 12164
rect 205726 12044 205732 12096
rect 205784 12084 205790 12096
rect 455690 12084 455696 12096
rect 205784 12056 455696 12084
rect 205784 12044 205790 12056
rect 455690 12044 455696 12056
rect 455748 12044 455754 12096
rect 128906 11976 128912 12028
rect 128964 12016 128970 12028
rect 178954 12016 178960 12028
rect 128964 11988 178960 12016
rect 128964 11976 128970 11988
rect 178954 11976 178960 11988
rect 179012 11976 179018 12028
rect 205818 11976 205824 12028
rect 205876 12016 205882 12028
rect 459186 12016 459192 12028
rect 205876 11988 459192 12016
rect 205876 11976 205882 11988
rect 459186 11976 459192 11988
rect 459244 11976 459250 12028
rect 99834 11908 99840 11960
rect 99892 11948 99898 11960
rect 167270 11948 167276 11960
rect 99892 11920 167276 11948
rect 99892 11908 99898 11920
rect 167270 11908 167276 11920
rect 167328 11908 167334 11960
rect 207014 11908 207020 11960
rect 207072 11948 207078 11960
rect 465810 11948 465816 11960
rect 207072 11920 465816 11948
rect 207072 11908 207078 11920
rect 465810 11908 465816 11920
rect 465868 11908 465874 11960
rect 77386 11840 77392 11892
rect 77444 11880 77450 11892
rect 165798 11880 165804 11892
rect 77444 11852 165804 11880
rect 77444 11840 77450 11852
rect 165798 11840 165804 11852
rect 165856 11840 165862 11892
rect 208762 11840 208768 11892
rect 208820 11880 208826 11892
rect 493042 11880 493048 11892
rect 208820 11852 493048 11880
rect 208820 11840 208826 11852
rect 493042 11840 493048 11852
rect 493100 11840 493106 11892
rect 53282 11772 53288 11824
rect 53340 11812 53346 11824
rect 163222 11812 163228 11824
rect 53340 11784 163228 11812
rect 53340 11772 53346 11784
rect 163222 11772 163228 11784
rect 163280 11772 163286 11824
rect 166074 11772 166080 11824
rect 166132 11812 166138 11824
rect 179046 11812 179052 11824
rect 166132 11784 179052 11812
rect 166132 11772 166138 11784
rect 179046 11772 179052 11784
rect 179104 11772 179110 11824
rect 211246 11772 211252 11824
rect 211304 11812 211310 11824
rect 523770 11812 523776 11824
rect 211304 11784 523776 11812
rect 211304 11772 211310 11784
rect 523770 11772 523776 11784
rect 523828 11772 523834 11824
rect 8754 11704 8760 11756
rect 8812 11744 8818 11756
rect 161014 11744 161020 11756
rect 8812 11716 161020 11744
rect 8812 11704 8818 11716
rect 161014 11704 161020 11716
rect 161072 11704 161078 11756
rect 176654 11704 176660 11756
rect 176712 11744 176718 11756
rect 177850 11744 177856 11756
rect 176712 11716 177856 11744
rect 176712 11704 176718 11716
rect 177850 11704 177856 11716
rect 177908 11704 177914 11756
rect 211154 11704 211160 11756
rect 211212 11744 211218 11756
rect 527818 11744 527824 11756
rect 211212 11716 527824 11744
rect 211212 11704 211218 11716
rect 527818 11704 527824 11716
rect 527876 11704 527882 11756
rect 143534 11636 143540 11688
rect 143592 11676 143598 11688
rect 144730 11676 144736 11688
rect 143592 11648 144736 11676
rect 143592 11636 143598 11648
rect 144730 11636 144736 11648
rect 144788 11636 144794 11688
rect 192110 11636 192116 11688
rect 192168 11676 192174 11688
rect 276106 11676 276112 11688
rect 192168 11648 276112 11676
rect 192168 11636 192174 11648
rect 276106 11636 276112 11648
rect 276164 11636 276170 11688
rect 182358 11432 182364 11484
rect 182416 11472 182422 11484
rect 184198 11472 184204 11484
rect 182416 11444 184204 11472
rect 182416 11432 182422 11444
rect 184198 11432 184204 11444
rect 184256 11432 184262 11484
rect 192754 10548 192760 10600
rect 192812 10588 192818 10600
rect 279050 10588 279056 10600
rect 192812 10560 279056 10588
rect 192812 10548 192818 10560
rect 279050 10548 279056 10560
rect 279108 10548 279114 10600
rect 118786 10480 118792 10532
rect 118844 10520 118850 10532
rect 168558 10520 168564 10532
rect 118844 10492 168564 10520
rect 118844 10480 118850 10492
rect 168558 10480 168564 10492
rect 168616 10480 168622 10532
rect 194502 10480 194508 10532
rect 194560 10520 194566 10532
rect 297266 10520 297272 10532
rect 194560 10492 297272 10520
rect 194560 10480 194566 10492
rect 297266 10480 297272 10492
rect 297324 10480 297330 10532
rect 100754 10412 100760 10464
rect 100812 10452 100818 10464
rect 167178 10452 167184 10464
rect 100812 10424 167184 10452
rect 100812 10412 100818 10424
rect 167178 10412 167184 10424
rect 167236 10412 167242 10464
rect 201770 10412 201776 10464
rect 201828 10452 201834 10464
rect 398926 10452 398932 10464
rect 201828 10424 398932 10452
rect 201828 10412 201834 10424
rect 398926 10412 398932 10424
rect 398984 10412 398990 10464
rect 97442 10344 97448 10396
rect 97500 10384 97506 10396
rect 167822 10384 167828 10396
rect 97500 10356 167828 10384
rect 97500 10344 97506 10356
rect 167822 10344 167828 10356
rect 167880 10344 167886 10396
rect 187142 10344 187148 10396
rect 187200 10384 187206 10396
rect 194594 10384 194600 10396
rect 187200 10356 194600 10384
rect 187200 10344 187206 10356
rect 194594 10344 194600 10356
rect 194652 10344 194658 10396
rect 208670 10344 208676 10396
rect 208728 10384 208734 10396
rect 486418 10384 486424 10396
rect 208728 10356 486424 10384
rect 208728 10344 208734 10356
rect 486418 10344 486424 10356
rect 486476 10344 486482 10396
rect 86402 10276 86408 10328
rect 86460 10316 86466 10328
rect 166442 10316 166448 10328
rect 86460 10288 166448 10316
rect 86460 10276 86466 10288
rect 166442 10276 166448 10288
rect 166500 10276 166506 10328
rect 186590 10276 186596 10328
rect 186648 10316 186654 10328
rect 206186 10316 206192 10328
rect 186648 10288 206192 10316
rect 186648 10276 186654 10288
rect 206186 10276 206192 10288
rect 206244 10276 206250 10328
rect 215478 10276 215484 10328
rect 215536 10316 215542 10328
rect 575106 10316 575112 10328
rect 215536 10288 575112 10316
rect 215536 10276 215542 10288
rect 575106 10276 575112 10288
rect 575164 10276 575170 10328
rect 197538 9596 197544 9648
rect 197596 9636 197602 9648
rect 344554 9636 344560 9648
rect 197596 9608 344560 9636
rect 197596 9596 197602 9608
rect 344554 9596 344560 9608
rect 344612 9596 344618 9648
rect 253474 9528 253480 9580
rect 253532 9568 253538 9580
rect 413094 9568 413100 9580
rect 253532 9540 413100 9568
rect 253532 9528 253538 9540
rect 413094 9528 413100 9540
rect 413152 9528 413158 9580
rect 198918 9460 198924 9512
rect 198976 9500 198982 9512
rect 361114 9500 361120 9512
rect 198976 9472 361120 9500
rect 198976 9460 198982 9472
rect 361114 9460 361120 9472
rect 361172 9460 361178 9512
rect 188154 9392 188160 9444
rect 188212 9432 188218 9444
rect 220446 9432 220452 9444
rect 188212 9404 220452 9432
rect 188212 9392 188218 9404
rect 220446 9392 220452 9404
rect 220504 9392 220510 9444
rect 253566 9392 253572 9444
rect 253624 9432 253630 9444
rect 430850 9432 430856 9444
rect 253624 9404 430856 9432
rect 253624 9392 253630 9404
rect 430850 9392 430856 9404
rect 430908 9392 430914 9444
rect 189166 9324 189172 9376
rect 189224 9364 189230 9376
rect 241698 9364 241704 9376
rect 189224 9336 241704 9364
rect 189224 9324 189230 9336
rect 241698 9324 241704 9336
rect 241756 9324 241762 9376
rect 253198 9324 253204 9376
rect 253256 9364 253262 9376
rect 434438 9364 434444 9376
rect 253256 9336 434444 9364
rect 253256 9324 253262 9336
rect 434438 9324 434444 9336
rect 434496 9324 434502 9376
rect 200114 9256 200120 9308
rect 200172 9296 200178 9308
rect 388254 9296 388260 9308
rect 200172 9268 388260 9296
rect 200172 9256 200178 9268
rect 388254 9256 388260 9268
rect 388312 9256 388318 9308
rect 200206 9188 200212 9240
rect 200264 9228 200270 9240
rect 391842 9228 391848 9240
rect 200264 9200 391848 9228
rect 200264 9188 200270 9200
rect 391842 9188 391848 9200
rect 391900 9188 391906 9240
rect 202874 9120 202880 9172
rect 202932 9160 202938 9172
rect 420178 9160 420184 9172
rect 202932 9132 420184 9160
rect 202932 9120 202938 9132
rect 420178 9120 420184 9132
rect 420236 9120 420242 9172
rect 119890 9052 119896 9104
rect 119948 9092 119954 9104
rect 169202 9092 169208 9104
rect 119948 9064 169208 9092
rect 119948 9052 119954 9064
rect 169202 9052 169208 9064
rect 169260 9052 169266 9104
rect 206738 9052 206744 9104
rect 206796 9092 206802 9104
rect 460382 9092 460388 9104
rect 206796 9064 460388 9092
rect 206796 9052 206802 9064
rect 460382 9052 460388 9064
rect 460440 9052 460446 9104
rect 71498 8984 71504 9036
rect 71556 9024 71562 9036
rect 161474 9024 161480 9036
rect 71556 8996 161480 9024
rect 71556 8984 71562 8996
rect 161474 8984 161480 8996
rect 161532 8984 161538 9036
rect 208578 8984 208584 9036
rect 208636 9024 208642 9036
rect 482830 9024 482836 9036
rect 208636 8996 482836 9024
rect 208636 8984 208642 8996
rect 482830 8984 482836 8996
rect 482888 8984 482894 9036
rect 45462 8916 45468 8968
rect 45520 8956 45526 8968
rect 163130 8956 163136 8968
rect 45520 8928 163136 8956
rect 45520 8916 45526 8928
rect 163130 8916 163136 8928
rect 163188 8916 163194 8968
rect 208486 8916 208492 8968
rect 208544 8956 208550 8968
rect 485222 8956 485228 8968
rect 208544 8928 485228 8956
rect 208544 8916 208550 8928
rect 485222 8916 485228 8928
rect 485280 8916 485286 8968
rect 253290 8848 253296 8900
rect 253348 8888 253354 8900
rect 381170 8888 381176 8900
rect 253348 8860 381176 8888
rect 253348 8848 253354 8860
rect 381170 8848 381176 8860
rect 381228 8848 381234 8900
rect 194778 7964 194784 8016
rect 194836 8004 194842 8016
rect 315022 8004 315028 8016
rect 194836 7976 315028 8004
rect 194836 7964 194842 7976
rect 315022 7964 315028 7976
rect 315080 7964 315086 8016
rect 197446 7896 197452 7948
rect 197504 7936 197510 7948
rect 350442 7936 350448 7948
rect 197504 7908 350448 7936
rect 197504 7896 197510 7908
rect 350442 7896 350448 7908
rect 350500 7896 350506 7948
rect 84470 7828 84476 7880
rect 84528 7868 84534 7880
rect 166350 7868 166356 7880
rect 84528 7840 166356 7868
rect 84528 7828 84534 7840
rect 166350 7828 166356 7840
rect 166408 7828 166414 7880
rect 197354 7828 197360 7880
rect 197412 7868 197418 7880
rect 352834 7868 352840 7880
rect 197412 7840 352840 7868
rect 197412 7828 197418 7840
rect 352834 7828 352840 7840
rect 352892 7828 352898 7880
rect 64322 7760 64328 7812
rect 64380 7800 64386 7812
rect 164418 7800 164424 7812
rect 64380 7772 164424 7800
rect 64380 7760 64386 7772
rect 164418 7760 164424 7772
rect 164476 7760 164482 7812
rect 198826 7760 198832 7812
rect 198884 7800 198890 7812
rect 367002 7800 367008 7812
rect 198884 7772 367008 7800
rect 198884 7760 198890 7772
rect 367002 7760 367008 7772
rect 367060 7760 367066 7812
rect 59630 7692 59636 7744
rect 59688 7732 59694 7744
rect 165430 7732 165436 7744
rect 59688 7704 165436 7732
rect 59688 7692 59694 7704
rect 165430 7692 165436 7704
rect 165488 7692 165494 7744
rect 201678 7692 201684 7744
rect 201736 7732 201742 7744
rect 406010 7732 406016 7744
rect 201736 7704 406016 7732
rect 201736 7692 201742 7704
rect 406010 7692 406016 7704
rect 406068 7692 406074 7744
rect 48958 7624 48964 7676
rect 49016 7664 49022 7676
rect 163038 7664 163044 7676
rect 49016 7636 163044 7664
rect 49016 7624 49022 7636
rect 163038 7624 163044 7636
rect 163096 7624 163102 7676
rect 209866 7624 209872 7676
rect 209924 7664 209930 7676
rect 510062 7664 510068 7676
rect 209924 7636 510068 7664
rect 209924 7624 209930 7636
rect 510062 7624 510068 7636
rect 510120 7624 510126 7676
rect 27706 7556 27712 7608
rect 27764 7596 27770 7608
rect 161566 7596 161572 7608
rect 27764 7568 161572 7596
rect 27764 7556 27770 7568
rect 161566 7556 161572 7568
rect 161624 7556 161630 7608
rect 215386 7556 215392 7608
rect 215444 7596 215450 7608
rect 571518 7596 571524 7608
rect 215444 7568 571524 7596
rect 215444 7556 215450 7568
rect 571518 7556 571524 7568
rect 571576 7556 571582 7608
rect 3418 6808 3424 6860
rect 3476 6848 3482 6860
rect 135990 6848 135996 6860
rect 3476 6820 135996 6848
rect 3476 6808 3482 6820
rect 135990 6808 135996 6820
rect 136048 6808 136054 6860
rect 187786 6808 187792 6860
rect 187844 6848 187850 6860
rect 216858 6848 216864 6860
rect 187844 6820 216864 6848
rect 187844 6808 187850 6820
rect 216858 6808 216864 6820
rect 216916 6808 216922 6860
rect 269758 6808 269764 6860
rect 269816 6848 269822 6860
rect 580166 6848 580172 6860
rect 269816 6820 580172 6848
rect 269816 6808 269822 6820
rect 580166 6808 580172 6820
rect 580224 6808 580230 6860
rect 187878 6740 187884 6792
rect 187936 6780 187942 6792
rect 222746 6780 222752 6792
rect 187936 6752 222752 6780
rect 187936 6740 187942 6752
rect 222746 6740 222752 6752
rect 222804 6740 222810 6792
rect 256234 6740 256240 6792
rect 256292 6780 256298 6792
rect 327994 6780 328000 6792
rect 256292 6752 328000 6780
rect 256292 6740 256298 6752
rect 327994 6740 328000 6752
rect 328052 6740 328058 6792
rect 191834 6672 191840 6724
rect 191892 6712 191898 6724
rect 270034 6712 270040 6724
rect 191892 6684 270040 6712
rect 191892 6672 191898 6684
rect 270034 6672 270040 6684
rect 270092 6672 270098 6724
rect 187970 6604 187976 6656
rect 188028 6644 188034 6656
rect 226426 6644 226432 6656
rect 188028 6616 226432 6644
rect 188028 6604 188034 6616
rect 226426 6604 226432 6616
rect 226484 6604 226490 6656
rect 256602 6604 256608 6656
rect 256660 6644 256666 6656
rect 342162 6644 342168 6656
rect 256660 6616 342168 6644
rect 256660 6604 256666 6616
rect 342162 6604 342168 6616
rect 342220 6604 342226 6656
rect 193306 6536 193312 6588
rect 193364 6576 193370 6588
rect 299658 6576 299664 6588
rect 193364 6548 299664 6576
rect 193364 6536 193370 6548
rect 299658 6536 299664 6548
rect 299716 6536 299722 6588
rect 194686 6468 194692 6520
rect 194744 6508 194750 6520
rect 311434 6508 311440 6520
rect 194744 6480 311440 6508
rect 194744 6468 194750 6480
rect 311434 6468 311440 6480
rect 311492 6468 311498 6520
rect 188062 6400 188068 6452
rect 188120 6440 188126 6452
rect 229830 6440 229836 6452
rect 188120 6412 229836 6440
rect 188120 6400 188126 6412
rect 229830 6400 229836 6412
rect 229888 6400 229894 6452
rect 256326 6400 256332 6452
rect 256384 6440 256390 6452
rect 377674 6440 377680 6452
rect 256384 6412 377680 6440
rect 256384 6400 256390 6412
rect 377674 6400 377680 6412
rect 377732 6400 377738 6452
rect 162486 6332 162492 6384
rect 162544 6372 162550 6384
rect 182910 6372 182916 6384
rect 162544 6344 182916 6372
rect 162544 6332 162550 6344
rect 182910 6332 182916 6344
rect 182968 6332 182974 6384
rect 201586 6332 201592 6384
rect 201644 6372 201650 6384
rect 403618 6372 403624 6384
rect 201644 6344 403624 6372
rect 201644 6332 201650 6344
rect 403618 6332 403624 6344
rect 403676 6332 403682 6384
rect 105722 6264 105728 6316
rect 105780 6304 105786 6316
rect 167730 6304 167736 6316
rect 105780 6276 167736 6304
rect 105780 6264 105786 6276
rect 167730 6264 167736 6276
rect 167788 6264 167794 6316
rect 204254 6264 204260 6316
rect 204312 6304 204318 6316
rect 437934 6304 437940 6316
rect 204312 6276 437940 6304
rect 204312 6264 204318 6276
rect 437934 6264 437940 6276
rect 437992 6264 437998 6316
rect 66714 6196 66720 6248
rect 66772 6236 66778 6248
rect 165062 6236 165068 6248
rect 66772 6208 165068 6236
rect 66772 6196 66778 6208
rect 165062 6196 165068 6208
rect 165120 6196 165126 6248
rect 209774 6196 209780 6248
rect 209832 6236 209838 6248
rect 502978 6236 502984 6248
rect 209832 6208 502984 6236
rect 209832 6196 209838 6208
rect 502978 6196 502984 6208
rect 503036 6196 503042 6248
rect 52546 6128 52552 6180
rect 52604 6168 52610 6180
rect 162946 6168 162952 6180
rect 52604 6140 162952 6168
rect 52604 6128 52610 6140
rect 162946 6128 162952 6140
rect 163004 6128 163010 6180
rect 213914 6128 213920 6180
rect 213972 6168 213978 6180
rect 553762 6168 553768 6180
rect 213972 6140 553768 6168
rect 213972 6128 213978 6140
rect 553762 6128 553768 6140
rect 553820 6128 553826 6180
rect 256142 6060 256148 6112
rect 256200 6100 256206 6112
rect 306742 6100 306748 6112
rect 256200 6072 306748 6100
rect 256200 6060 256206 6072
rect 306742 6060 306748 6072
rect 306800 6060 306806 6112
rect 253382 5992 253388 6044
rect 253440 6032 253446 6044
rect 290182 6032 290188 6044
rect 253440 6004 290188 6032
rect 253440 5992 253446 6004
rect 290182 5992 290188 6004
rect 290240 5992 290246 6044
rect 185118 5516 185124 5568
rect 185176 5556 185182 5568
rect 188522 5556 188528 5568
rect 185176 5528 188528 5556
rect 185176 5516 185182 5528
rect 188522 5516 188528 5528
rect 188580 5516 188586 5568
rect 195606 5108 195612 5160
rect 195664 5148 195670 5160
rect 307938 5148 307944 5160
rect 195664 5120 307944 5148
rect 195664 5108 195670 5120
rect 307938 5108 307944 5120
rect 307996 5108 308002 5160
rect 195974 5040 195980 5092
rect 196032 5080 196038 5092
rect 323302 5080 323308 5092
rect 196032 5052 323308 5080
rect 196032 5040 196038 5052
rect 323302 5040 323308 5052
rect 323360 5040 323366 5092
rect 18230 4972 18236 5024
rect 18288 5012 18294 5024
rect 160922 5012 160928 5024
rect 18288 4984 160928 5012
rect 18288 4972 18294 4984
rect 160922 4972 160928 4984
rect 160980 4972 160986 5024
rect 198734 4972 198740 5024
rect 198792 5012 198798 5024
rect 368198 5012 368204 5024
rect 198792 4984 368204 5012
rect 198792 4972 198798 4984
rect 368198 4972 368204 4984
rect 368256 4972 368262 5024
rect 44266 4904 44272 4956
rect 44324 4944 44330 4956
rect 163590 4944 163596 4956
rect 44324 4916 163596 4944
rect 44324 4904 44330 4916
rect 163590 4904 163596 4916
rect 163648 4904 163654 4956
rect 201494 4904 201500 4956
rect 201552 4944 201558 4956
rect 402514 4944 402520 4956
rect 201552 4916 402520 4944
rect 201552 4904 201558 4916
rect 402514 4904 402520 4916
rect 402572 4904 402578 4956
rect 492306 4944 492312 4956
rect 470566 4916 492312 4944
rect 31294 4836 31300 4888
rect 31352 4876 31358 4888
rect 162302 4876 162308 4888
rect 31352 4848 162308 4876
rect 31352 4836 31358 4848
rect 162302 4836 162308 4848
rect 162360 4836 162366 4888
rect 208394 4836 208400 4888
rect 208452 4876 208458 4888
rect 470566 4876 470594 4916
rect 492306 4904 492312 4916
rect 492364 4904 492370 4956
rect 208452 4848 470594 4876
rect 208452 4836 208458 4848
rect 160094 4768 160100 4820
rect 160152 4808 160158 4820
rect 182726 4808 182732 4820
rect 160152 4780 182732 4808
rect 160152 4768 160158 4780
rect 182726 4768 182732 4780
rect 182784 4768 182790 4820
rect 215294 4768 215300 4820
rect 215352 4808 215358 4820
rect 576302 4808 576308 4820
rect 215352 4780 576308 4808
rect 215352 4768 215358 4780
rect 576302 4768 576308 4780
rect 576360 4768 576366 4820
rect 276014 4156 276020 4208
rect 276072 4196 276078 4208
rect 276750 4196 276756 4208
rect 276072 4168 276756 4196
rect 276072 4156 276078 4168
rect 276750 4156 276756 4168
rect 276808 4156 276814 4208
rect 284294 4156 284300 4208
rect 284352 4196 284358 4208
rect 285030 4196 285036 4208
rect 284352 4168 285036 4196
rect 284352 4156 284358 4168
rect 285030 4156 285036 4168
rect 285088 4156 285094 4208
rect 124674 4088 124680 4140
rect 124732 4128 124738 4140
rect 159358 4128 159364 4140
rect 124732 4100 159364 4128
rect 124732 4088 124738 4100
rect 159358 4088 159364 4100
rect 159416 4088 159422 4140
rect 168466 4088 168472 4140
rect 168524 4128 168530 4140
rect 173158 4128 173164 4140
rect 168524 4100 173164 4128
rect 168524 4088 168530 4100
rect 173158 4088 173164 4100
rect 173216 4088 173222 4140
rect 189718 4088 189724 4140
rect 189776 4128 189782 4140
rect 190822 4128 190828 4140
rect 189776 4100 190828 4128
rect 189776 4088 189782 4100
rect 190822 4088 190828 4100
rect 190880 4088 190886 4140
rect 193214 4088 193220 4140
rect 193272 4128 193278 4140
rect 296070 4128 296076 4140
rect 193272 4100 296076 4128
rect 193272 4088 193278 4100
rect 296070 4088 296076 4100
rect 296128 4088 296134 4140
rect 92750 4020 92756 4072
rect 92808 4060 92814 4072
rect 134794 4060 134800 4072
rect 92808 4032 134800 4060
rect 92808 4020 92814 4032
rect 134794 4020 134800 4032
rect 134852 4020 134858 4072
rect 189994 4020 190000 4072
rect 190052 4060 190058 4072
rect 201494 4060 201500 4072
rect 190052 4032 201500 4060
rect 190052 4020 190058 4032
rect 201494 4020 201500 4032
rect 201552 4020 201558 4072
rect 259086 4020 259092 4072
rect 259144 4060 259150 4072
rect 440234 4060 440240 4072
rect 259144 4032 440240 4060
rect 259144 4020 259150 4032
rect 440234 4020 440240 4032
rect 440292 4020 440298 4072
rect 89162 3952 89168 4004
rect 89220 3992 89226 4004
rect 133138 3992 133144 4004
rect 89220 3964 133144 3992
rect 89220 3952 89226 3964
rect 133138 3952 133144 3964
rect 133196 3952 133202 4004
rect 191190 3952 191196 4004
rect 191248 3992 191254 4004
rect 205082 3992 205088 4004
rect 191248 3964 205088 3992
rect 191248 3952 191254 3964
rect 205082 3952 205088 3964
rect 205140 3952 205146 4004
rect 258810 3952 258816 4004
rect 258868 3992 258874 4004
rect 448514 3992 448520 4004
rect 258868 3964 448520 3992
rect 258868 3952 258874 3964
rect 448514 3952 448520 3964
rect 448572 3952 448578 4004
rect 462958 3952 462964 4004
rect 463016 3992 463022 4004
rect 487614 3992 487620 4004
rect 463016 3964 487620 3992
rect 463016 3952 463022 3964
rect 487614 3952 487620 3964
rect 487672 3952 487678 4004
rect 57238 3884 57244 3936
rect 57296 3924 57302 3936
rect 133230 3924 133236 3936
rect 57296 3896 133236 3924
rect 57296 3884 57302 3896
rect 133230 3884 133236 3896
rect 133288 3884 133294 3936
rect 134150 3884 134156 3936
rect 134208 3924 134214 3936
rect 177390 3924 177396 3936
rect 134208 3896 177396 3924
rect 134208 3884 134214 3896
rect 177390 3884 177396 3896
rect 177448 3884 177454 3936
rect 186406 3884 186412 3936
rect 186464 3924 186470 3936
rect 200298 3924 200304 3936
rect 186464 3896 200304 3924
rect 186464 3884 186470 3896
rect 200298 3884 200304 3896
rect 200356 3884 200362 3936
rect 213178 3884 213184 3936
rect 213236 3924 213242 3936
rect 225138 3924 225144 3936
rect 213236 3896 225144 3924
rect 213236 3884 213242 3896
rect 225138 3884 225144 3896
rect 225196 3884 225202 3936
rect 260098 3884 260104 3936
rect 260156 3924 260162 3936
rect 461578 3924 461584 3936
rect 260156 3896 461584 3924
rect 260156 3884 260162 3896
rect 461578 3884 461584 3896
rect 461636 3884 461642 3936
rect 468478 3884 468484 3936
rect 468536 3924 468542 3936
rect 511258 3924 511264 3936
rect 468536 3896 511264 3924
rect 468536 3884 468542 3896
rect 511258 3884 511264 3896
rect 511316 3884 511322 3936
rect 25314 3816 25320 3868
rect 25372 3856 25378 3868
rect 137278 3856 137284 3868
rect 25372 3828 137284 3856
rect 25372 3816 25378 3828
rect 137278 3816 137284 3828
rect 137336 3816 137342 3868
rect 150618 3816 150624 3868
rect 150676 3856 150682 3868
rect 173250 3856 173256 3868
rect 150676 3828 173256 3856
rect 150676 3816 150682 3828
rect 173250 3816 173256 3828
rect 173308 3816 173314 3868
rect 186314 3816 186320 3868
rect 186372 3856 186378 3868
rect 210970 3856 210976 3868
rect 186372 3828 210976 3856
rect 186372 3816 186378 3828
rect 210970 3816 210976 3828
rect 211028 3816 211034 3868
rect 258902 3816 258908 3868
rect 258960 3856 258966 3868
rect 480530 3856 480536 3868
rect 258960 3828 480536 3856
rect 258960 3816 258966 3828
rect 480530 3816 480536 3828
rect 480588 3816 480594 3868
rect 43070 3748 43076 3800
rect 43128 3788 43134 3800
rect 159450 3788 159456 3800
rect 43128 3760 159456 3788
rect 43128 3748 43134 3760
rect 159450 3748 159456 3760
rect 159508 3748 159514 3800
rect 186498 3748 186504 3800
rect 186556 3788 186562 3800
rect 207382 3788 207388 3800
rect 186556 3760 207388 3788
rect 186556 3748 186562 3760
rect 207382 3748 207388 3760
rect 207440 3748 207446 3800
rect 207842 3748 207848 3800
rect 207900 3788 207906 3800
rect 433242 3788 433248 3800
rect 207900 3760 433248 3788
rect 207900 3748 207906 3760
rect 433242 3748 433248 3760
rect 433300 3748 433306 3800
rect 479518 3748 479524 3800
rect 479576 3788 479582 3800
rect 526622 3788 526628 3800
rect 479576 3760 526628 3788
rect 479576 3748 479582 3760
rect 526622 3748 526628 3760
rect 526680 3748 526686 3800
rect 11146 3680 11152 3732
rect 11204 3720 11210 3732
rect 134518 3720 134524 3732
rect 11204 3692 134524 3720
rect 11204 3680 11210 3692
rect 134518 3680 134524 3692
rect 134576 3680 134582 3732
rect 136450 3680 136456 3732
rect 136508 3720 136514 3732
rect 177482 3720 177488 3732
rect 136508 3692 177488 3720
rect 136508 3680 136514 3692
rect 177482 3680 177488 3692
rect 177540 3680 177546 3732
rect 188614 3680 188620 3732
rect 188672 3720 188678 3732
rect 203886 3720 203892 3732
rect 188672 3692 203892 3720
rect 188672 3680 188678 3692
rect 203886 3680 203892 3692
rect 203944 3680 203950 3732
rect 203978 3680 203984 3732
rect 204036 3720 204042 3732
rect 246390 3720 246396 3732
rect 204036 3692 246396 3720
rect 204036 3680 204042 3692
rect 246390 3680 246396 3692
rect 246448 3680 246454 3732
rect 258994 3680 259000 3732
rect 259052 3720 259058 3732
rect 484026 3720 484032 3732
rect 259052 3692 484032 3720
rect 259052 3680 259058 3692
rect 484026 3680 484032 3692
rect 484084 3680 484090 3732
rect 6454 3612 6460 3664
rect 6512 3652 6518 3664
rect 138658 3652 138664 3664
rect 6512 3624 138664 3652
rect 6512 3612 6518 3624
rect 138658 3612 138664 3624
rect 138716 3612 138722 3664
rect 142430 3612 142436 3664
rect 142488 3652 142494 3664
rect 178770 3652 178776 3664
rect 142488 3624 178776 3652
rect 142488 3612 142494 3624
rect 178770 3612 178776 3624
rect 178828 3612 178834 3664
rect 188798 3612 188804 3664
rect 188856 3652 188862 3664
rect 219250 3652 219256 3664
rect 188856 3624 219256 3652
rect 188856 3612 188862 3624
rect 219250 3612 219256 3624
rect 219308 3612 219314 3664
rect 224218 3612 224224 3664
rect 224276 3652 224282 3664
rect 450078 3652 450084 3664
rect 224276 3624 450084 3652
rect 224276 3612 224282 3624
rect 450078 3612 450084 3624
rect 450136 3612 450142 3664
rect 450538 3612 450544 3664
rect 450596 3652 450602 3664
rect 523034 3652 523040 3664
rect 450596 3624 523040 3652
rect 450596 3612 450602 3624
rect 523034 3612 523040 3624
rect 523092 3612 523098 3664
rect 24210 3544 24216 3596
rect 24268 3584 24274 3596
rect 158162 3584 158168 3596
rect 24268 3556 158168 3584
rect 24268 3544 24274 3556
rect 158162 3544 158168 3556
rect 158220 3544 158226 3596
rect 164878 3544 164884 3596
rect 164936 3584 164942 3596
rect 174538 3584 174544 3596
rect 164936 3556 174544 3584
rect 164936 3544 164942 3556
rect 174538 3544 174544 3556
rect 174596 3544 174602 3596
rect 184934 3544 184940 3596
rect 184992 3584 184998 3596
rect 185854 3584 185860 3596
rect 184992 3556 185860 3584
rect 184992 3544 184998 3556
rect 185854 3544 185860 3556
rect 185912 3544 185918 3596
rect 189074 3544 189080 3596
rect 189132 3584 189138 3596
rect 234614 3584 234620 3596
rect 189132 3556 234620 3584
rect 189132 3544 189138 3556
rect 234614 3544 234620 3556
rect 234672 3544 234678 3596
rect 258718 3544 258724 3596
rect 258776 3584 258782 3596
rect 501782 3584 501788 3596
rect 258776 3556 501788 3584
rect 258776 3544 258782 3556
rect 501782 3544 501788 3556
rect 501840 3544 501846 3596
rect 514754 3544 514760 3596
rect 514812 3584 514818 3596
rect 515582 3584 515588 3596
rect 514812 3556 515588 3584
rect 514812 3544 514818 3556
rect 515582 3544 515588 3556
rect 515640 3544 515646 3596
rect 531314 3544 531320 3596
rect 531372 3584 531378 3596
rect 532142 3584 532148 3596
rect 531372 3556 532148 3584
rect 531372 3544 531378 3556
rect 532142 3544 532148 3556
rect 532200 3544 532206 3596
rect 539594 3544 539600 3596
rect 539652 3584 539658 3596
rect 540422 3584 540428 3596
rect 539652 3556 540428 3584
rect 539652 3544 539658 3556
rect 540422 3544 540428 3556
rect 540480 3544 540486 3596
rect 17034 3476 17040 3528
rect 17092 3516 17098 3528
rect 18598 3516 18604 3528
rect 17092 3488 18604 3516
rect 17092 3476 17098 3488
rect 18598 3476 18604 3488
rect 18656 3476 18662 3528
rect 19426 3476 19432 3528
rect 19484 3516 19490 3528
rect 158070 3516 158076 3528
rect 19484 3488 158076 3516
rect 19484 3476 19490 3488
rect 158070 3476 158076 3488
rect 158128 3476 158134 3528
rect 161290 3476 161296 3528
rect 161348 3516 161354 3528
rect 161348 3488 173112 3516
rect 161348 3476 161354 3488
rect 566 3408 572 3460
rect 624 3448 630 3460
rect 157978 3448 157984 3460
rect 624 3420 157984 3448
rect 624 3408 630 3420
rect 157978 3408 157984 3420
rect 158036 3408 158042 3460
rect 158898 3408 158904 3460
rect 158956 3448 158962 3460
rect 158956 3420 161474 3448
rect 158956 3408 158962 3420
rect 60734 3340 60740 3392
rect 60792 3380 60798 3392
rect 61654 3380 61660 3392
rect 60792 3352 61660 3380
rect 60792 3340 60798 3352
rect 61654 3340 61660 3352
rect 61712 3340 61718 3392
rect 77294 3340 77300 3392
rect 77352 3380 77358 3392
rect 78214 3380 78220 3392
rect 77352 3352 78220 3380
rect 77352 3340 77358 3352
rect 78214 3340 78220 3352
rect 78272 3340 78278 3392
rect 102134 3340 102140 3392
rect 102192 3380 102198 3392
rect 103330 3380 103336 3392
rect 102192 3352 103336 3380
rect 102192 3340 102198 3352
rect 103330 3340 103336 3352
rect 103388 3340 103394 3392
rect 106918 3340 106924 3392
rect 106976 3380 106982 3392
rect 134610 3380 134616 3392
rect 106976 3352 134616 3380
rect 106976 3340 106982 3352
rect 134610 3340 134616 3352
rect 134668 3340 134674 3392
rect 117590 3272 117596 3324
rect 117648 3312 117654 3324
rect 134702 3312 134708 3324
rect 117648 3284 134708 3312
rect 117648 3272 117654 3284
rect 134702 3272 134708 3284
rect 134760 3272 134766 3324
rect 161446 3312 161474 3420
rect 168374 3408 168380 3460
rect 168432 3448 168438 3460
rect 169570 3448 169576 3460
rect 168432 3420 169576 3448
rect 168432 3408 168438 3420
rect 169570 3408 169576 3420
rect 169628 3408 169634 3460
rect 173084 3380 173112 3488
rect 173158 3476 173164 3528
rect 173216 3516 173222 3528
rect 174630 3516 174636 3528
rect 173216 3488 174636 3516
rect 173216 3476 173222 3488
rect 174630 3476 174636 3488
rect 174688 3476 174694 3528
rect 189810 3476 189816 3528
rect 189868 3516 189874 3528
rect 189868 3488 211752 3516
rect 189868 3476 189874 3488
rect 174262 3408 174268 3460
rect 174320 3448 174326 3460
rect 178862 3448 178868 3460
rect 174320 3420 178868 3448
rect 174320 3408 174326 3420
rect 178862 3408 178868 3420
rect 178920 3408 178926 3460
rect 191466 3408 191472 3460
rect 191524 3448 191530 3460
rect 211724 3448 211752 3488
rect 211798 3476 211804 3528
rect 211856 3516 211862 3528
rect 213362 3516 213368 3528
rect 211856 3488 213368 3516
rect 211856 3476 211862 3488
rect 213362 3476 213368 3488
rect 213420 3476 213426 3528
rect 217318 3476 217324 3528
rect 217376 3516 217382 3528
rect 217376 3488 473216 3516
rect 217376 3476 217382 3488
rect 215662 3448 215668 3460
rect 191524 3420 209774 3448
rect 211724 3420 215668 3448
rect 191524 3408 191530 3420
rect 177298 3380 177304 3392
rect 173084 3352 177304 3380
rect 177298 3340 177304 3352
rect 177356 3340 177362 3392
rect 188430 3340 188436 3392
rect 188488 3380 188494 3392
rect 188488 3352 190454 3380
rect 188488 3340 188494 3352
rect 178678 3312 178684 3324
rect 161446 3284 178684 3312
rect 178678 3272 178684 3284
rect 178736 3272 178742 3324
rect 184842 3272 184848 3324
rect 184900 3312 184906 3324
rect 189718 3312 189724 3324
rect 184900 3284 189724 3312
rect 184900 3272 184906 3284
rect 189718 3272 189724 3284
rect 189776 3272 189782 3324
rect 190426 3312 190454 3352
rect 191098 3340 191104 3392
rect 191156 3380 191162 3392
rect 202690 3380 202696 3392
rect 191156 3352 202696 3380
rect 191156 3340 191162 3352
rect 202690 3340 202696 3352
rect 202748 3340 202754 3392
rect 199102 3312 199108 3324
rect 190426 3284 199108 3312
rect 199102 3272 199108 3284
rect 199160 3272 199166 3324
rect 190086 3204 190092 3256
rect 190144 3244 190150 3256
rect 197906 3244 197912 3256
rect 190144 3216 197912 3244
rect 190144 3204 190150 3216
rect 197906 3204 197912 3216
rect 197964 3204 197970 3256
rect 209746 3244 209774 3420
rect 215662 3408 215668 3420
rect 215720 3408 215726 3460
rect 226334 3408 226340 3460
rect 226392 3448 226398 3460
rect 227530 3448 227536 3460
rect 226392 3420 227536 3448
rect 226392 3408 226398 3420
rect 227530 3408 227536 3420
rect 227588 3408 227594 3460
rect 229066 3420 238754 3448
rect 210418 3340 210424 3392
rect 210476 3380 210482 3392
rect 212166 3380 212172 3392
rect 210476 3352 212172 3380
rect 210476 3340 210482 3352
rect 212166 3340 212172 3352
rect 212224 3340 212230 3392
rect 229066 3244 229094 3420
rect 238726 3380 238754 3420
rect 251174 3408 251180 3460
rect 251232 3448 251238 3460
rect 252370 3448 252376 3460
rect 251232 3420 252376 3448
rect 251232 3408 251238 3420
rect 252370 3408 252376 3420
rect 252428 3408 252434 3460
rect 256050 3408 256056 3460
rect 256108 3448 256114 3460
rect 256108 3420 258074 3448
rect 256108 3408 256114 3420
rect 257062 3380 257068 3392
rect 238726 3352 257068 3380
rect 257062 3340 257068 3352
rect 257120 3340 257126 3392
rect 258046 3380 258074 3420
rect 271138 3408 271144 3460
rect 271196 3448 271202 3460
rect 271196 3420 470594 3448
rect 271196 3408 271202 3420
rect 292574 3380 292580 3392
rect 258046 3352 292580 3380
rect 292574 3340 292580 3352
rect 292632 3340 292638 3392
rect 299474 3340 299480 3392
rect 299532 3380 299538 3392
rect 300762 3380 300768 3392
rect 299532 3352 300768 3380
rect 299532 3340 299538 3352
rect 300762 3340 300768 3352
rect 300820 3340 300826 3392
rect 307754 3340 307760 3392
rect 307812 3380 307818 3392
rect 309042 3380 309048 3392
rect 307812 3352 309048 3380
rect 307812 3340 307818 3352
rect 309042 3340 309048 3352
rect 309100 3340 309106 3392
rect 316034 3340 316040 3392
rect 316092 3380 316098 3392
rect 317322 3380 317328 3392
rect 316092 3352 317328 3380
rect 316092 3340 316098 3352
rect 317322 3340 317328 3352
rect 317380 3340 317386 3392
rect 324406 3340 324412 3392
rect 324464 3380 324470 3392
rect 325602 3380 325608 3392
rect 324464 3352 325608 3380
rect 324464 3340 324470 3352
rect 325602 3340 325608 3352
rect 325660 3340 325666 3392
rect 332594 3340 332600 3392
rect 332652 3380 332658 3392
rect 333882 3380 333888 3392
rect 332652 3352 333888 3380
rect 332652 3340 332658 3352
rect 333882 3340 333888 3352
rect 333940 3340 333946 3392
rect 357434 3340 357440 3392
rect 357492 3380 357498 3392
rect 358722 3380 358728 3392
rect 357492 3352 358728 3380
rect 357492 3340 357498 3352
rect 358722 3340 358728 3352
rect 358780 3340 358786 3392
rect 373994 3340 374000 3392
rect 374052 3380 374058 3392
rect 375282 3380 375288 3392
rect 374052 3352 375288 3380
rect 374052 3340 374058 3352
rect 375282 3340 375288 3352
rect 375340 3340 375346 3392
rect 382274 3340 382280 3392
rect 382332 3380 382338 3392
rect 383562 3380 383568 3392
rect 382332 3352 383568 3380
rect 382332 3340 382338 3352
rect 383562 3340 383568 3352
rect 383620 3340 383626 3392
rect 398926 3340 398932 3392
rect 398984 3380 398990 3392
rect 400122 3380 400128 3392
rect 398984 3352 400128 3380
rect 398984 3340 398990 3352
rect 400122 3340 400128 3352
rect 400180 3340 400186 3392
rect 407206 3340 407212 3392
rect 407264 3380 407270 3392
rect 408402 3380 408408 3392
rect 407264 3352 408408 3380
rect 407264 3340 407270 3352
rect 408402 3340 408408 3352
rect 408460 3340 408466 3392
rect 415394 3340 415400 3392
rect 415452 3380 415458 3392
rect 416682 3380 416688 3392
rect 415452 3352 416688 3380
rect 415452 3340 415458 3352
rect 416682 3340 416688 3352
rect 416740 3340 416746 3392
rect 423674 3340 423680 3392
rect 423732 3380 423738 3392
rect 424962 3380 424968 3392
rect 423732 3352 424968 3380
rect 423732 3340 423738 3352
rect 424962 3340 424968 3352
rect 425020 3340 425026 3392
rect 440326 3340 440332 3392
rect 440384 3380 440390 3392
rect 441522 3380 441528 3392
rect 440384 3352 441528 3380
rect 440384 3340 440390 3352
rect 441522 3340 441528 3352
rect 441580 3340 441586 3392
rect 448606 3340 448612 3392
rect 448664 3380 448670 3392
rect 449802 3380 449808 3392
rect 448664 3352 449808 3380
rect 448664 3340 448670 3352
rect 449802 3340 449808 3352
rect 449860 3340 449866 3392
rect 456794 3340 456800 3392
rect 456852 3380 456858 3392
rect 458082 3380 458088 3392
rect 456852 3352 458088 3380
rect 456852 3340 456858 3352
rect 458082 3340 458088 3352
rect 458140 3340 458146 3392
rect 256418 3272 256424 3324
rect 256476 3312 256482 3324
rect 288986 3312 288992 3324
rect 256476 3284 288992 3312
rect 256476 3272 256482 3284
rect 288986 3272 288992 3284
rect 289044 3272 289050 3324
rect 470566 3312 470594 3420
rect 473188 3380 473216 3488
rect 473354 3476 473360 3528
rect 473412 3516 473418 3528
rect 474182 3516 474188 3528
rect 473412 3488 474188 3516
rect 473412 3476 473418 3488
rect 474182 3476 474188 3488
rect 474240 3476 474246 3528
rect 487798 3476 487804 3528
rect 487856 3516 487862 3528
rect 556154 3516 556160 3528
rect 487856 3488 556160 3516
rect 487856 3476 487862 3488
rect 556154 3476 556160 3488
rect 556212 3476 556218 3528
rect 572714 3476 572720 3528
rect 572772 3516 572778 3528
rect 573542 3516 573548 3528
rect 572772 3488 573548 3516
rect 572772 3476 572778 3488
rect 573542 3476 573548 3488
rect 573600 3476 573606 3528
rect 583386 3448 583392 3460
rect 480226 3420 583392 3448
rect 479334 3380 479340 3392
rect 473188 3352 479340 3380
rect 479334 3340 479340 3352
rect 479392 3340 479398 3392
rect 480226 3312 480254 3420
rect 583386 3408 583392 3420
rect 583444 3408 583450 3460
rect 489914 3340 489920 3392
rect 489972 3380 489978 3392
rect 490742 3380 490748 3392
rect 489972 3352 490748 3380
rect 489972 3340 489978 3352
rect 490742 3340 490748 3352
rect 490800 3340 490806 3392
rect 470566 3284 480254 3312
rect 209746 3216 229094 3244
rect 255958 3204 255964 3256
rect 256016 3244 256022 3256
rect 274818 3244 274824 3256
rect 256016 3216 274824 3244
rect 256016 3204 256022 3216
rect 274818 3204 274824 3216
rect 274876 3204 274882 3256
rect 189902 3136 189908 3188
rect 189960 3176 189966 3188
rect 193214 3176 193220 3188
rect 189960 3148 193220 3176
rect 189960 3136 189966 3148
rect 193214 3136 193220 3148
rect 193272 3136 193278 3188
rect 203518 3136 203524 3188
rect 203576 3176 203582 3188
rect 208578 3176 208584 3188
rect 203576 3148 208584 3176
rect 203576 3136 203582 3148
rect 208578 3136 208584 3148
rect 208636 3136 208642 3188
rect 256510 3136 256516 3188
rect 256568 3176 256574 3188
rect 271230 3176 271236 3188
rect 256568 3148 271236 3176
rect 256568 3136 256574 3148
rect 271230 3136 271236 3148
rect 271288 3136 271294 3188
rect 132954 3068 132960 3120
rect 133012 3108 133018 3120
rect 135898 3108 135904 3120
rect 133012 3080 135904 3108
rect 133012 3068 133018 3080
rect 135898 3068 135904 3080
rect 135956 3068 135962 3120
rect 214466 2864 214472 2916
rect 214524 2904 214530 2916
rect 216674 2904 216680 2916
rect 214524 2876 216680 2904
rect 214524 2864 214530 2876
rect 216674 2864 216680 2876
rect 216732 2864 216738 2916
rect 207014 2796 207020 2848
rect 207072 2836 207078 2848
rect 209774 2836 209780 2848
rect 207072 2808 209780 2836
rect 207072 2796 207078 2808
rect 209774 2796 209780 2808
rect 209832 2796 209838 2848
rect 450078 2796 450084 2848
rect 450136 2836 450142 2848
rect 450906 2836 450912 2848
rect 450136 2808 450912 2836
rect 450136 2796 450142 2808
rect 450906 2796 450912 2808
rect 450964 2796 450970 2848
<< via1 >>
rect 246396 700952 246448 701004
rect 332508 700952 332560 701004
rect 246488 700884 246540 700936
rect 348792 700884 348844 700936
rect 243636 700816 243688 700868
rect 364984 700816 365036 700868
rect 240784 700748 240836 700800
rect 397460 700748 397512 700800
rect 253296 700680 253348 700732
rect 429844 700680 429896 700732
rect 218704 700612 218756 700664
rect 413652 700612 413704 700664
rect 105452 700544 105504 700596
rect 142804 700544 142856 700596
rect 249064 700544 249116 700596
rect 462320 700544 462372 700596
rect 89168 700476 89220 700528
rect 151084 700476 151136 700528
rect 233884 700476 233936 700528
rect 478512 700476 478564 700528
rect 72976 700408 73028 700460
rect 148324 700408 148376 700460
rect 243544 700408 243596 700460
rect 494796 700408 494848 700460
rect 24308 700340 24360 700392
rect 138664 700340 138716 700392
rect 240968 700340 241020 700392
rect 527180 700340 527232 700392
rect 40500 700272 40552 700324
rect 157984 700272 158036 700324
rect 202788 700272 202840 700324
rect 218152 700272 218204 700324
rect 232504 700272 232556 700324
rect 543464 700272 543516 700324
rect 253204 700204 253256 700256
rect 300124 700204 300176 700256
rect 251824 700136 251876 700188
rect 283840 700136 283892 700188
rect 238024 700068 238076 700120
rect 267648 700068 267700 700120
rect 239404 696940 239456 696992
rect 580172 696940 580224 696992
rect 3424 683136 3476 683188
rect 158076 683136 158128 683188
rect 221464 683136 221516 683188
rect 580172 683136 580224 683188
rect 3516 670692 3568 670744
rect 141424 670692 141476 670744
rect 3424 656888 3476 656940
rect 144184 656888 144236 656940
rect 234160 644512 234212 644564
rect 251272 644512 251324 644564
rect 233976 644444 234028 644496
rect 251180 644444 251232 644496
rect 234252 643084 234304 643136
rect 251180 643084 251232 643136
rect 231124 641724 231176 641776
rect 251180 641724 251232 641776
rect 239496 640296 239548 640348
rect 251180 640296 251232 640348
rect 224224 638936 224276 638988
rect 251180 638936 251232 638988
rect 228364 637576 228416 637628
rect 251180 637576 251232 637628
rect 244924 634788 244976 634840
rect 251180 634788 251232 634840
rect 225604 633428 225656 633480
rect 251272 633428 251324 633480
rect 228456 632680 228508 632732
rect 251180 632680 251232 632732
rect 3424 632068 3476 632120
rect 158168 632068 158220 632120
rect 220084 632068 220136 632120
rect 251180 632068 251232 632120
rect 232596 630640 232648 630692
rect 251180 630640 251232 630692
rect 222844 629280 222896 629332
rect 251180 629280 251232 629332
rect 231216 627920 231268 627972
rect 251180 627920 251232 627972
rect 231308 626560 231360 626612
rect 251180 626560 251232 626612
rect 245016 625132 245068 625184
rect 251180 625132 251232 625184
rect 236644 623840 236696 623892
rect 251272 623840 251324 623892
rect 228548 623772 228600 623824
rect 251180 623772 251232 623824
rect 222936 622412 222988 622464
rect 251180 622412 251232 622464
rect 242164 620984 242216 621036
rect 251180 620984 251232 621036
rect 226984 619624 227036 619676
rect 251180 619624 251232 619676
rect 3148 618264 3200 618316
rect 146944 618264 146996 618316
rect 224316 618264 224368 618316
rect 251180 618264 251232 618316
rect 221648 616836 221700 616888
rect 251180 616836 251232 616888
rect 574744 616836 574796 616888
rect 580172 616836 580224 616888
rect 239588 615476 239640 615528
rect 251180 615476 251232 615528
rect 235264 614116 235316 614168
rect 251180 614116 251232 614168
rect 246580 612824 246632 612876
rect 251272 612824 251324 612876
rect 221740 612756 221792 612808
rect 251180 612756 251232 612808
rect 238116 611328 238168 611380
rect 251180 611328 251232 611380
rect 229744 609968 229796 610020
rect 251180 609968 251232 610020
rect 229836 608608 229888 608660
rect 251180 608608 251232 608660
rect 221832 607180 221884 607232
rect 251180 607180 251232 607232
rect 3240 605820 3292 605872
rect 135904 605820 135956 605872
rect 238208 604460 238260 604512
rect 251180 604460 251232 604512
rect 227076 603100 227128 603152
rect 251180 603100 251232 603152
rect 249156 601672 249208 601724
rect 251272 601672 251324 601724
rect 235356 600312 235408 600364
rect 251180 600312 251232 600364
rect 232688 598952 232740 599004
rect 251180 598952 251232 599004
rect 247776 597524 247828 597576
rect 251180 597524 251232 597576
rect 247868 594804 247920 594856
rect 251180 594804 251232 594856
rect 223028 593376 223080 593428
rect 251180 593376 251232 593428
rect 243728 592016 243780 592068
rect 251180 592016 251232 592068
rect 111800 590724 111852 590776
rect 119620 590724 119672 590776
rect 246672 590724 246724 590776
rect 251180 590724 251232 590776
rect 111892 590656 111944 590708
rect 140044 590656 140096 590708
rect 220176 590656 220228 590708
rect 251272 590656 251324 590708
rect 111800 589364 111852 589416
rect 123484 589364 123536 589416
rect 111892 589296 111944 589348
rect 142896 589296 142948 589348
rect 241060 589296 241112 589348
rect 251180 589296 251232 589348
rect 111800 587868 111852 587920
rect 123576 587868 123628 587920
rect 229928 587868 229980 587920
rect 251180 587868 251232 587920
rect 111800 586508 111852 586560
rect 123760 586508 123812 586560
rect 112260 585760 112312 585812
rect 123668 585760 123720 585812
rect 111800 585352 111852 585404
rect 113824 585352 113876 585404
rect 245108 585148 245160 585200
rect 251180 585148 251232 585200
rect 111984 584400 112036 584452
rect 120724 584400 120776 584452
rect 111892 583856 111944 583908
rect 113916 583856 113968 583908
rect 111800 583720 111852 583772
rect 117964 583720 118016 583772
rect 232780 583720 232832 583772
rect 251180 583720 251232 583772
rect 111800 582360 111852 582412
rect 115204 582360 115256 582412
rect 230020 582360 230072 582412
rect 251180 582360 251232 582412
rect 111892 581612 111944 581664
rect 138756 581612 138808 581664
rect 111800 581000 111852 581052
rect 122104 581000 122156 581052
rect 220268 581000 220320 581052
rect 251180 581000 251232 581052
rect 111984 580252 112036 580304
rect 122196 580252 122248 580304
rect 111892 579708 111944 579760
rect 116768 579708 116820 579760
rect 249340 579708 249392 579760
rect 251272 579708 251324 579760
rect 3332 579640 3384 579692
rect 29644 579640 29696 579692
rect 111800 579640 111852 579692
rect 134524 579640 134576 579692
rect 242256 579640 242308 579692
rect 251180 579640 251232 579692
rect 111800 578280 111852 578332
rect 130384 578280 130436 578332
rect 111892 578212 111944 578264
rect 133144 578212 133196 578264
rect 227168 578212 227220 578264
rect 251180 578212 251232 578264
rect 249432 576988 249484 577040
rect 251272 576988 251324 577040
rect 111800 576852 111852 576904
rect 152556 576852 152608 576904
rect 111892 575560 111944 575612
rect 132040 575560 132092 575612
rect 111800 575492 111852 575544
rect 141516 575492 141568 575544
rect 239680 575492 239732 575544
rect 251180 575492 251232 575544
rect 111892 574336 111944 574388
rect 114008 574336 114060 574388
rect 111800 574064 111852 574116
rect 152648 574064 152700 574116
rect 231400 574064 231452 574116
rect 251180 574064 251232 574116
rect 111800 572772 111852 572824
rect 134616 572772 134668 572824
rect 111892 572704 111944 572756
rect 142988 572704 143040 572756
rect 227260 572704 227312 572756
rect 251180 572704 251232 572756
rect 111800 571412 111852 571464
rect 130476 571412 130528 571464
rect 111892 571344 111944 571396
rect 133236 571344 133288 571396
rect 220360 571344 220412 571396
rect 251180 571344 251232 571396
rect 111800 569984 111852 570036
rect 122288 569984 122340 570036
rect 111984 569916 112036 569968
rect 127624 569916 127676 569968
rect 238300 569916 238352 569968
rect 251180 569916 251232 569968
rect 111892 568624 111944 568676
rect 137284 568624 137336 568676
rect 234344 568624 234396 568676
rect 251272 568624 251324 568676
rect 111800 568556 111852 568608
rect 152740 568556 152792 568608
rect 225696 568556 225748 568608
rect 251180 568556 251232 568608
rect 111800 567196 111852 567248
rect 141608 567196 141660 567248
rect 220452 567196 220504 567248
rect 251180 567196 251232 567248
rect 111800 565904 111852 565956
rect 116584 565904 116636 565956
rect 3424 565836 3476 565888
rect 29736 565836 29788 565888
rect 111892 565836 111944 565888
rect 134708 565836 134760 565888
rect 236736 565836 236788 565888
rect 251180 565836 251232 565888
rect 111800 564476 111852 564528
rect 127716 564476 127768 564528
rect 111892 564408 111944 564460
rect 130568 564408 130620 564460
rect 234436 564408 234488 564460
rect 251180 564408 251232 564460
rect 112444 563660 112496 563712
rect 122380 563660 122432 563712
rect 111800 563048 111852 563100
rect 140136 563048 140188 563100
rect 242348 563048 242400 563100
rect 251180 563048 251232 563100
rect 111984 562300 112036 562352
rect 144276 562300 144328 562352
rect 111800 561688 111852 561740
rect 115296 561688 115348 561740
rect 243820 561688 243872 561740
rect 251180 561688 251232 561740
rect 111800 560260 111852 560312
rect 140228 560260 140280 560312
rect 236828 560260 236880 560312
rect 251180 560260 251232 560312
rect 111800 558968 111852 559020
rect 115388 558968 115440 559020
rect 111892 558900 111944 558952
rect 118056 558900 118108 558952
rect 234528 558900 234580 558952
rect 251180 558900 251232 558952
rect 111800 557608 111852 557660
rect 127808 557608 127860 557660
rect 245200 557608 245252 557660
rect 251180 557608 251232 557660
rect 111892 557540 111944 557592
rect 130660 557540 130712 557592
rect 223120 557540 223172 557592
rect 251272 557540 251324 557592
rect 112628 556792 112680 556844
rect 148416 556792 148468 556844
rect 111800 556180 111852 556232
rect 147036 556180 147088 556232
rect 246764 556180 246816 556232
rect 251180 556180 251232 556232
rect 111800 554888 111852 554940
rect 115480 554888 115532 554940
rect 111892 554752 111944 554804
rect 151176 554752 151228 554804
rect 236920 554752 236972 554804
rect 251180 554752 251232 554804
rect 111984 554004 112036 554056
rect 119344 554004 119396 554056
rect 111800 553392 111852 553444
rect 138848 553392 138900 553444
rect 232872 553392 232924 553444
rect 251180 553392 251232 553444
rect 112536 552644 112588 552696
rect 113088 552644 113140 552696
rect 111892 552100 111944 552152
rect 126244 552100 126296 552152
rect 111800 552032 111852 552084
rect 149704 552032 149756 552084
rect 221924 552032 221976 552084
rect 251180 552032 251232 552084
rect 111800 550672 111852 550724
rect 116676 550672 116728 550724
rect 111892 550604 111944 550656
rect 130752 550604 130804 550656
rect 220544 550604 220596 550656
rect 251180 550604 251232 550656
rect 111800 549312 111852 549364
rect 119436 549312 119488 549364
rect 111892 549244 111944 549296
rect 153844 549244 153896 549296
rect 247960 549244 248012 549296
rect 251180 549244 251232 549296
rect 112076 548496 112128 548548
rect 143080 548496 143132 548548
rect 111800 548088 111852 548140
rect 115572 548088 115624 548140
rect 235448 547952 235500 548004
rect 251272 547952 251324 548004
rect 111892 547884 111944 547936
rect 126520 547884 126572 547936
rect 232964 547884 233016 547936
rect 251180 547884 251232 547936
rect 111800 546456 111852 546508
rect 152832 546456 152884 546508
rect 231492 546456 231544 546508
rect 251180 546456 251232 546508
rect 111892 545164 111944 545216
rect 118148 545164 118200 545216
rect 111800 545096 111852 545148
rect 131764 545096 131816 545148
rect 227352 545096 227404 545148
rect 251180 545096 251232 545148
rect 111800 543736 111852 543788
rect 144368 543736 144420 543788
rect 227444 543736 227496 543788
rect 251180 543736 251232 543788
rect 116768 542988 116820 543040
rect 155224 542988 155276 543040
rect 111892 542444 111944 542496
rect 116860 542444 116912 542496
rect 111800 542376 111852 542428
rect 119528 542376 119580 542428
rect 113088 541628 113140 541680
rect 149796 541628 149848 541680
rect 111800 540948 111852 541000
rect 116768 540948 116820 541000
rect 249524 540948 249576 541000
rect 251180 540948 251232 541000
rect 111800 539588 111852 539640
rect 137376 539588 137428 539640
rect 235540 539588 235592 539640
rect 251180 539588 251232 539640
rect 111800 538296 111852 538348
rect 127900 538296 127952 538348
rect 111892 538228 111944 538280
rect 151268 538228 151320 538280
rect 235632 538228 235684 538280
rect 251180 538228 251232 538280
rect 111800 536868 111852 536920
rect 129004 536868 129056 536920
rect 111892 536800 111944 536852
rect 131856 536800 131908 536852
rect 235724 536800 235776 536852
rect 251180 536800 251232 536852
rect 111892 535508 111944 535560
rect 148508 535508 148560 535560
rect 111800 535440 111852 535492
rect 151360 535440 151412 535492
rect 220636 535440 220688 535492
rect 251180 535440 251232 535492
rect 113088 534692 113140 534744
rect 145564 534692 145616 534744
rect 111800 534080 111852 534132
rect 143172 534080 143224 534132
rect 235816 534080 235868 534132
rect 251180 534080 251232 534132
rect 111892 533740 111944 533792
rect 116952 533740 117004 533792
rect 113088 532720 113140 532772
rect 147128 532720 147180 532772
rect 113088 531360 113140 531412
rect 138940 531360 138992 531412
rect 112260 531292 112312 531344
rect 148600 531292 148652 531344
rect 112260 531156 112312 531208
rect 112628 531156 112680 531208
rect 112444 530000 112496 530052
rect 113088 530000 113140 530052
rect 131948 530000 132000 530052
rect 112628 529932 112680 529984
rect 153936 529932 153988 529984
rect 112444 529796 112496 529848
rect 249248 529320 249300 529372
rect 580632 529320 580684 529372
rect 247684 529252 247736 529304
rect 580172 529252 580224 529304
rect 112260 529184 112312 529236
rect 123852 529184 123904 529236
rect 132040 529184 132092 529236
rect 155316 529184 155368 529236
rect 240876 529184 240928 529236
rect 580540 529184 580592 529236
rect 112352 528572 112404 528624
rect 124864 528572 124916 528624
rect 111800 527212 111852 527264
rect 114100 527212 114152 527264
rect 2964 527144 3016 527196
rect 29828 527144 29880 527196
rect 112352 525852 112404 525904
rect 139032 525852 139084 525904
rect 113088 525784 113140 525836
rect 144460 525784 144512 525836
rect 112260 525716 112312 525768
rect 117044 525716 117096 525768
rect 112076 524424 112128 524476
rect 147220 524424 147272 524476
rect 221556 524424 221608 524476
rect 580172 524424 580224 524476
rect 111892 523064 111944 523116
rect 132040 523064 132092 523116
rect 111800 522996 111852 523048
rect 143264 522996 143316 523048
rect 111892 521704 111944 521756
rect 118240 521704 118292 521756
rect 111800 521636 111852 521688
rect 126336 521636 126388 521688
rect 112904 521160 112956 521212
rect 113180 521160 113232 521212
rect 113088 520888 113140 520940
rect 149888 520888 149940 520940
rect 111800 520344 111852 520396
rect 120816 520344 120868 520396
rect 111892 520276 111944 520328
rect 124956 520276 125008 520328
rect 111800 519596 111852 519648
rect 118332 519596 118384 519648
rect 112812 519528 112864 519580
rect 145748 519528 145800 519580
rect 112352 518168 112404 518220
rect 154028 518168 154080 518220
rect 111800 517488 111852 517540
rect 144552 517488 144604 517540
rect 111892 516196 111944 516248
rect 119712 516196 119764 516248
rect 111800 516128 111852 516180
rect 140320 516128 140372 516180
rect 113088 515380 113140 515432
rect 130844 515380 130896 515432
rect 111800 514836 111852 514888
rect 114192 514836 114244 514888
rect 3516 514768 3568 514820
rect 29920 514768 29972 514820
rect 111892 514768 111944 514820
rect 120908 514768 120960 514820
rect 111800 513408 111852 513460
rect 125048 513408 125100 513460
rect 111892 513340 111944 513392
rect 145656 513340 145708 513392
rect 112260 512592 112312 512644
rect 147312 512592 147364 512644
rect 111800 511980 111852 512032
rect 139124 511980 139176 512032
rect 111892 510688 111944 510740
rect 117136 510688 117188 510740
rect 111800 510620 111852 510672
rect 141700 510620 141752 510672
rect 234068 510620 234120 510672
rect 580172 510620 580224 510672
rect 111984 509872 112036 509924
rect 121000 509872 121052 509924
rect 111800 509260 111852 509312
rect 143356 509260 143408 509312
rect 112996 508512 113048 508564
rect 122656 508512 122708 508564
rect 111892 507900 111944 507952
rect 126612 507900 126664 507952
rect 111800 507832 111852 507884
rect 141792 507832 141844 507884
rect 111800 506472 111852 506524
rect 129096 506472 129148 506524
rect 111892 505724 111944 505776
rect 147404 505724 147456 505776
rect 111800 505112 111852 505164
rect 126428 505112 126480 505164
rect 126520 504364 126572 504416
rect 155500 504364 155552 504416
rect 111800 503888 111852 503940
rect 114284 503888 114336 503940
rect 111892 503684 111944 503736
rect 121092 503684 121144 503736
rect 111800 502392 111852 502444
rect 140412 502392 140464 502444
rect 111892 502324 111944 502376
rect 140504 502324 140556 502376
rect 111800 500964 111852 501016
rect 148692 500964 148744 501016
rect 111800 499672 111852 499724
rect 115664 499672 115716 499724
rect 111984 499536 112036 499588
rect 133328 499536 133380 499588
rect 111892 498788 111944 498840
rect 141884 498788 141936 498840
rect 111800 498176 111852 498228
rect 127992 498176 128044 498228
rect 126612 497428 126664 497480
rect 155408 497428 155460 497480
rect 233056 497428 233108 497480
rect 252192 497428 252244 497480
rect 111800 496884 111852 496936
rect 119804 496884 119856 496936
rect 111892 496816 111944 496868
rect 126796 496816 126848 496868
rect 111984 496068 112036 496120
rect 135996 496068 136048 496120
rect 111800 495728 111852 495780
rect 115756 495728 115808 495780
rect 111892 495456 111944 495508
rect 121184 495456 121236 495508
rect 225788 495456 225840 495508
rect 251180 495456 251232 495508
rect 111800 495048 111852 495100
rect 114376 495048 114428 495100
rect 111800 494028 111852 494080
rect 148784 494028 148836 494080
rect 225880 494028 225932 494080
rect 251180 494028 251232 494080
rect 111800 492668 111852 492720
rect 151452 492668 151504 492720
rect 243912 492668 243964 492720
rect 251180 492668 251232 492720
rect 111800 491376 111852 491428
rect 122472 491376 122524 491428
rect 111892 491308 111944 491360
rect 126704 491308 126756 491360
rect 225972 491308 226024 491360
rect 251180 491308 251232 491360
rect 111800 489948 111852 490000
rect 128084 489948 128136 490000
rect 111892 489880 111944 489932
rect 129188 489880 129240 489932
rect 224408 489880 224460 489932
rect 251180 489880 251232 489932
rect 111892 488588 111944 488640
rect 126520 488588 126572 488640
rect 111800 488520 111852 488572
rect 137468 488520 137520 488572
rect 241152 488520 241204 488572
rect 251180 488520 251232 488572
rect 111800 487228 111852 487280
rect 118424 487228 118476 487280
rect 111892 487160 111944 487212
rect 144644 487160 144696 487212
rect 238392 487160 238444 487212
rect 251180 487160 251232 487212
rect 111892 485868 111944 485920
rect 137560 485868 137612 485920
rect 111800 485800 111852 485852
rect 151544 485800 151596 485852
rect 246856 485800 246908 485852
rect 251180 485800 251232 485852
rect 113088 485052 113140 485104
rect 140596 485052 140648 485104
rect 111800 484372 111852 484424
rect 134800 484372 134852 484424
rect 224500 484372 224552 484424
rect 251180 484372 251232 484424
rect 111800 483080 111852 483132
rect 123944 483080 123996 483132
rect 111892 483012 111944 483064
rect 133420 483012 133472 483064
rect 224592 483012 224644 483064
rect 251180 483012 251232 483064
rect 111800 481720 111852 481772
rect 128176 481720 128228 481772
rect 111892 481652 111944 481704
rect 129280 481652 129332 481704
rect 224776 481652 224828 481704
rect 251180 481652 251232 481704
rect 126704 480904 126756 480956
rect 155592 480904 155644 480956
rect 111800 480292 111852 480344
rect 124036 480292 124088 480344
rect 111892 480224 111944 480276
rect 126612 480224 126664 480276
rect 224684 480224 224736 480276
rect 251180 480224 251232 480276
rect 239772 479476 239824 479528
rect 252376 479476 252428 479528
rect 111800 478932 111852 478984
rect 118516 478932 118568 478984
rect 111892 478864 111944 478916
rect 145840 478864 145892 478916
rect 249616 478864 249668 478916
rect 251180 478864 251232 478916
rect 111800 477640 111852 477692
rect 114468 477640 114520 477692
rect 111892 477504 111944 477556
rect 143448 477504 143500 477556
rect 223304 477504 223356 477556
rect 251180 477504 251232 477556
rect 112352 476756 112404 476808
rect 125232 476756 125284 476808
rect 111800 476076 111852 476128
rect 136088 476076 136140 476128
rect 223212 476076 223264 476128
rect 251180 476076 251232 476128
rect 111800 474784 111852 474836
rect 132132 474784 132184 474836
rect 111892 474716 111944 474768
rect 133512 474716 133564 474768
rect 227536 474716 227588 474768
rect 251180 474716 251232 474768
rect 111800 474036 111852 474088
rect 115848 474036 115900 474088
rect 111800 473424 111852 473476
rect 128268 473424 128320 473476
rect 111892 473356 111944 473408
rect 129372 473356 129424 473408
rect 242440 473356 242492 473408
rect 251180 473356 251232 473408
rect 111800 472064 111852 472116
rect 122564 472064 122616 472116
rect 111892 471996 111944 472048
rect 126704 471996 126756 472048
rect 224868 471996 224920 472048
rect 251180 471996 251232 472048
rect 111892 470636 111944 470688
rect 141976 470636 142028 470688
rect 111800 470568 111852 470620
rect 147496 470568 147548 470620
rect 230112 470568 230164 470620
rect 251180 470568 251232 470620
rect 111800 469344 111852 469396
rect 115112 469344 115164 469396
rect 245292 469276 245344 469328
rect 251180 469276 251232 469328
rect 111800 469208 111852 469260
rect 154120 469208 154172 469260
rect 227628 469208 227680 469260
rect 251272 469208 251324 469260
rect 111800 467916 111852 467968
rect 117228 467916 117280 467968
rect 111892 467848 111944 467900
rect 152924 467848 152976 467900
rect 111800 466488 111852 466540
rect 132224 466488 132276 466540
rect 111892 466420 111944 466472
rect 137652 466420 137704 466472
rect 230204 466420 230256 466472
rect 251180 466420 251232 466472
rect 111892 465128 111944 465180
rect 125140 465128 125192 465180
rect 111800 465060 111852 465112
rect 151636 465060 151688 465112
rect 249708 465060 249760 465112
rect 251640 465060 251692 465112
rect 111800 463768 111852 463820
rect 126888 463768 126940 463820
rect 111892 463700 111944 463752
rect 149980 463700 150032 463752
rect 244096 463700 244148 463752
rect 251180 463700 251232 463752
rect 111800 462408 111852 462460
rect 119896 462408 119948 462460
rect 111892 462340 111944 462392
rect 153016 462340 153068 462392
rect 244004 462340 244056 462392
rect 251180 462340 251232 462392
rect 111800 460980 111852 461032
rect 137744 460980 137796 461032
rect 111892 460912 111944 460964
rect 144736 460912 144788 460964
rect 237012 460164 237064 460216
rect 252100 460164 252152 460216
rect 111800 459552 111852 459604
rect 150072 459552 150124 459604
rect 226064 459552 226116 459604
rect 251180 459552 251232 459604
rect 111800 458260 111852 458312
rect 130936 458260 130988 458312
rect 111892 458192 111944 458244
rect 133604 458192 133656 458244
rect 248052 458192 248104 458244
rect 251180 458192 251232 458244
rect 111800 456764 111852 456816
rect 132316 456764 132368 456816
rect 238484 456764 238536 456816
rect 251180 456764 251232 456816
rect 573364 456764 573416 456816
rect 580172 456764 580224 456816
rect 111892 455472 111944 455524
rect 132408 455472 132460 455524
rect 111800 455404 111852 455456
rect 139216 455404 139268 455456
rect 239864 455404 239916 455456
rect 251180 455404 251232 455456
rect 111800 454520 111852 454572
rect 115020 454520 115072 454572
rect 111800 454044 111852 454096
rect 142068 454044 142120 454096
rect 223396 454044 223448 454096
rect 251180 454044 251232 454096
rect 111800 452684 111852 452736
rect 116400 452684 116452 452736
rect 111892 452616 111944 452668
rect 122748 452616 122800 452668
rect 111892 451324 111944 451376
rect 124128 451324 124180 451376
rect 111800 451256 111852 451308
rect 148876 451256 148928 451308
rect 241244 451256 241296 451308
rect 251180 451256 251232 451308
rect 119620 450508 119672 450560
rect 155684 450508 155736 450560
rect 111800 449964 111852 450016
rect 119252 449964 119304 450016
rect 111892 449896 111944 449948
rect 119988 449896 120040 449948
rect 226892 449896 226944 449948
rect 251180 449896 251232 449948
rect 111800 448604 111852 448656
rect 116492 448604 116544 448656
rect 111892 448536 111944 448588
rect 145932 448536 145984 448588
rect 223488 448536 223540 448588
rect 251180 448536 251232 448588
rect 111800 447108 111852 447160
rect 140688 447108 140740 447160
rect 231584 447108 231636 447160
rect 251180 447108 251232 447160
rect 251732 446428 251784 446480
rect 252284 446428 252336 446480
rect 251732 446292 251784 446344
rect 252468 446292 252520 446344
rect 226800 445748 226852 445800
rect 251180 445748 251232 445800
rect 242532 444388 242584 444440
rect 251180 444388 251232 444440
rect 231676 441600 231728 441652
rect 251180 441600 251232 441652
rect 228640 440240 228692 440292
rect 251180 440240 251232 440292
rect 230296 439492 230348 439544
rect 251732 439492 251784 439544
rect 222016 438880 222068 438932
rect 251180 438880 251232 438932
rect 246212 437452 246264 437504
rect 251180 437452 251232 437504
rect 246948 436160 247000 436212
rect 251180 436160 251232 436212
rect 231768 436092 231820 436144
rect 251272 436092 251324 436144
rect 226156 434732 226208 434784
rect 251180 434732 251232 434784
rect 238576 433304 238628 433356
rect 251180 433304 251232 433356
rect 224132 431944 224184 431996
rect 251180 431944 251232 431996
rect 228732 430584 228784 430636
rect 251180 430584 251232 430636
rect 158444 429836 158496 429888
rect 169760 429836 169812 429888
rect 245384 429156 245436 429208
rect 251180 429156 251232 429208
rect 239956 427796 240008 427848
rect 251180 427796 251232 427848
rect 245476 426504 245528 426556
rect 251272 426504 251324 426556
rect 228824 426436 228876 426488
rect 251180 426436 251232 426488
rect 222752 425076 222804 425128
rect 251180 425076 251232 425128
rect 248972 423648 249024 423700
rect 251180 423648 251232 423700
rect 3332 422288 3384 422340
rect 156604 422288 156656 422340
rect 228916 420928 228968 420980
rect 251180 420928 251232 420980
rect 226248 419500 226300 419552
rect 251180 419500 251232 419552
rect 242624 418140 242676 418192
rect 251180 418140 251232 418192
rect 244188 416780 244240 416832
rect 251180 416780 251232 416832
rect 229008 415488 229060 415540
rect 251272 415488 251324 415540
rect 224040 415420 224092 415472
rect 251180 415420 251232 415472
rect 245568 413992 245620 414044
rect 251180 413992 251232 414044
rect 219716 413924 219768 413976
rect 234252 413924 234304 413976
rect 219992 413856 220044 413908
rect 233976 413856 234028 413908
rect 220728 413788 220780 413840
rect 234160 413788 234212 413840
rect 219808 413720 219860 413772
rect 231124 413720 231176 413772
rect 248144 412632 248196 412684
rect 251180 412632 251232 412684
rect 220728 412564 220780 412616
rect 239496 412564 239548 412616
rect 219900 412088 219952 412140
rect 228364 412088 228416 412140
rect 220084 411884 220136 411936
rect 224224 411884 224276 411936
rect 223948 411272 224000 411324
rect 251180 411272 251232 411324
rect 220728 411204 220780 411256
rect 250444 411204 250496 411256
rect 219808 411136 219860 411188
rect 244924 411136 244976 411188
rect 220084 410932 220136 410984
rect 225604 410932 225656 410984
rect 3332 409844 3384 409896
rect 152464 409844 152516 409896
rect 233976 409844 234028 409896
rect 251180 409844 251232 409896
rect 220084 409776 220136 409828
rect 232596 409776 232648 409828
rect 220728 409708 220780 409760
rect 228456 409708 228508 409760
rect 219900 409640 219952 409692
rect 222844 409640 222896 409692
rect 123760 409096 123812 409148
rect 154672 409096 154724 409148
rect 234160 408484 234212 408536
rect 251180 408484 251232 408536
rect 140044 408416 140096 408468
rect 154948 408416 155000 408468
rect 220084 408416 220136 408468
rect 245016 408416 245068 408468
rect 219900 408348 219952 408400
rect 231308 408348 231360 408400
rect 220728 408280 220780 408332
rect 231216 408280 231268 408332
rect 117964 407736 118016 407788
rect 155776 407736 155828 407788
rect 231032 407124 231084 407176
rect 251180 407124 251232 407176
rect 123576 407056 123628 407108
rect 154856 407056 154908 407108
rect 220084 407056 220136 407108
rect 242164 407056 242216 407108
rect 123668 406988 123720 407040
rect 154764 406988 154816 407040
rect 220728 406988 220780 407040
rect 236644 406988 236696 407040
rect 123484 406920 123536 406972
rect 154948 406920 155000 406972
rect 142896 406852 142948 406904
rect 154580 406852 154632 406904
rect 220728 406648 220780 406700
rect 228548 406648 228600 406700
rect 219900 406376 219952 406428
rect 222936 406376 222988 406428
rect 113824 405628 113876 405680
rect 154764 405628 154816 405680
rect 220084 405628 220136 405680
rect 221648 405628 221700 405680
rect 113916 405560 113968 405612
rect 154856 405560 154908 405612
rect 155040 405560 155092 405612
rect 155316 405560 155368 405612
rect 120724 405492 120776 405544
rect 154948 405492 155000 405544
rect 123852 405424 123904 405476
rect 154580 405424 154632 405476
rect 220728 405356 220780 405408
rect 226984 405356 227036 405408
rect 219900 405288 219952 405340
rect 224316 405288 224368 405340
rect 222108 404336 222160 404388
rect 251180 404336 251232 404388
rect 115204 404268 115256 404320
rect 154672 404268 154724 404320
rect 219992 404268 220044 404320
rect 246580 404268 246632 404320
rect 122104 404200 122156 404252
rect 154948 404200 155000 404252
rect 220728 404200 220780 404252
rect 239588 404200 239640 404252
rect 122196 404132 122248 404184
rect 154856 404132 154908 404184
rect 220084 404132 220136 404184
rect 235264 404132 235316 404184
rect 138756 404064 138808 404116
rect 154764 404064 154816 404116
rect 219716 402908 219768 402960
rect 238116 402908 238168 402960
rect 130384 402840 130436 402892
rect 154764 402840 154816 402892
rect 220176 402840 220228 402892
rect 229836 402840 229888 402892
rect 133144 402772 133196 402824
rect 154856 402772 154908 402824
rect 220728 402772 220780 402824
rect 229744 402772 229796 402824
rect 134524 402704 134576 402756
rect 154672 402704 154724 402756
rect 219808 402704 219860 402756
rect 221740 402704 221792 402756
rect 122380 402636 122432 402688
rect 154948 402636 155000 402688
rect 152556 402432 152608 402484
rect 155224 402432 155276 402484
rect 231216 401616 231268 401668
rect 251180 401616 251232 401668
rect 152648 401548 152700 401600
rect 155224 401548 155276 401600
rect 220728 401548 220780 401600
rect 250536 401548 250588 401600
rect 141516 401480 141568 401532
rect 154856 401480 154908 401532
rect 220176 401480 220228 401532
rect 238208 401480 238260 401532
rect 142988 401412 143040 401464
rect 155040 401412 155092 401464
rect 114008 401344 114060 401396
rect 154948 401344 155000 401396
rect 220084 401276 220136 401328
rect 221832 401276 221884 401328
rect 122288 400868 122340 400920
rect 155132 400868 155184 400920
rect 229744 400868 229796 400920
rect 251640 400868 251692 400920
rect 251548 400800 251600 400852
rect 251916 400800 251968 400852
rect 127624 400120 127676 400172
rect 154764 400120 154816 400172
rect 220728 400120 220780 400172
rect 251548 400120 251600 400172
rect 130476 400052 130528 400104
rect 155040 400052 155092 400104
rect 220084 400052 220136 400104
rect 249156 400052 249208 400104
rect 133236 399984 133288 400036
rect 154856 399984 154908 400036
rect 220176 399984 220228 400036
rect 235356 399984 235408 400036
rect 134616 399916 134668 399968
rect 154948 399916 155000 399968
rect 219992 399916 220044 399968
rect 227076 399916 227128 399968
rect 226984 398828 227036 398880
rect 251180 398828 251232 398880
rect 152740 398760 152792 398812
rect 154580 398760 154632 398812
rect 220084 398760 220136 398812
rect 247776 398760 247828 398812
rect 141608 398692 141660 398744
rect 154672 398692 154724 398744
rect 220176 398692 220228 398744
rect 237012 398692 237064 398744
rect 144276 398624 144328 398676
rect 154856 398624 154908 398676
rect 220728 398624 220780 398676
rect 232688 398624 232740 398676
rect 149796 398556 149848 398608
rect 155040 398556 155092 398608
rect 137284 398488 137336 398540
rect 154948 398488 155000 398540
rect 127716 398080 127768 398132
rect 154764 398080 154816 398132
rect 251732 398080 251784 398132
rect 252468 398080 252520 398132
rect 3332 397468 3384 397520
rect 134524 397468 134576 397520
rect 222844 397468 222896 397520
rect 251180 397468 251232 397520
rect 116584 397400 116636 397452
rect 155040 397400 155092 397452
rect 220728 397400 220780 397452
rect 247868 397400 247920 397452
rect 122656 397332 122708 397384
rect 155132 397332 155184 397384
rect 220176 397332 220228 397384
rect 243728 397332 243780 397384
rect 130568 397264 130620 397316
rect 154856 397264 154908 397316
rect 134708 397196 134760 397248
rect 154948 397196 155000 397248
rect 220728 396856 220780 396908
rect 223028 396856 223080 396908
rect 247776 396040 247828 396092
rect 251180 396040 251232 396092
rect 112444 395972 112496 396024
rect 154764 395972 154816 396024
rect 155224 395972 155276 396024
rect 155500 395972 155552 396024
rect 220084 395972 220136 396024
rect 246672 395972 246724 396024
rect 115296 395904 115348 395956
rect 154856 395904 154908 395956
rect 220176 395904 220228 395956
rect 241060 395904 241112 395956
rect 140136 395836 140188 395888
rect 154948 395836 155000 395888
rect 220728 395836 220780 395888
rect 229928 395836 229980 395888
rect 140228 395768 140280 395820
rect 155040 395768 155092 395820
rect 148416 395700 148468 395752
rect 154672 395700 154724 395752
rect 127808 395292 127860 395344
rect 154948 395292 155000 395344
rect 221740 394680 221792 394732
rect 251180 394680 251232 394732
rect 115388 394612 115440 394664
rect 154580 394612 154632 394664
rect 220728 394612 220780 394664
rect 250628 394612 250680 394664
rect 118056 394544 118108 394596
rect 154672 394544 154724 394596
rect 219992 394544 220044 394596
rect 245108 394544 245160 394596
rect 130660 394476 130712 394528
rect 154764 394476 154816 394528
rect 220176 394476 220228 394528
rect 232780 394476 232832 394528
rect 147036 394408 147088 394460
rect 154856 394408 154908 394460
rect 129004 393932 129056 393984
rect 155132 393932 155184 393984
rect 250444 393864 250496 393916
rect 251916 393864 251968 393916
rect 221648 393320 221700 393372
rect 251180 393320 251232 393372
rect 151176 393252 151228 393304
rect 155040 393252 155092 393304
rect 220176 393252 220228 393304
rect 242256 393252 242308 393304
rect 119344 393184 119396 393236
rect 154948 393184 155000 393236
rect 220728 393184 220780 393236
rect 230020 393184 230072 393236
rect 138848 393116 138900 393168
rect 154764 393116 154816 393168
rect 143080 393048 143132 393100
rect 154856 393048 154908 393100
rect 115480 392980 115532 393032
rect 154948 392980 155000 393032
rect 220176 391960 220228 392012
rect 220452 391960 220504 392012
rect 236644 391960 236696 392012
rect 251180 391960 251232 392012
rect 220268 391892 220320 391944
rect 249432 391892 249484 391944
rect 126244 391824 126296 391876
rect 154948 391824 155000 391876
rect 220728 391824 220780 391876
rect 249340 391824 249392 391876
rect 130752 391756 130804 391808
rect 154764 391756 154816 391808
rect 220452 391756 220504 391808
rect 239680 391756 239732 391808
rect 149704 391688 149756 391740
rect 154672 391688 154724 391740
rect 116676 391620 116728 391672
rect 154948 391620 155000 391672
rect 220728 391484 220780 391536
rect 227168 391484 227220 391536
rect 219992 390532 220044 390584
rect 251180 390532 251232 390584
rect 152832 390464 152884 390516
rect 154580 390464 154632 390516
rect 220728 390464 220780 390516
rect 231400 390464 231452 390516
rect 118148 390396 118200 390448
rect 155040 390396 155092 390448
rect 119436 390328 119488 390380
rect 154948 390328 155000 390380
rect 219900 390328 219952 390380
rect 227260 390328 227312 390380
rect 145748 390260 145800 390312
rect 154856 390260 154908 390312
rect 115572 390192 115624 390244
rect 154948 390192 155000 390244
rect 119528 389784 119580 389836
rect 155224 389784 155276 389836
rect 219900 389172 219952 389224
rect 251180 389172 251232 389224
rect 116860 389104 116912 389156
rect 154856 389104 154908 389156
rect 220728 389104 220780 389156
rect 238300 389104 238352 389156
rect 130844 389036 130896 389088
rect 154764 389036 154816 389088
rect 220452 389036 220504 389088
rect 234344 389036 234396 389088
rect 131764 388968 131816 389020
rect 154672 388968 154724 389020
rect 220084 388968 220136 389020
rect 225696 388968 225748 389020
rect 144368 388900 144420 388952
rect 154948 388900 155000 388952
rect 251640 388424 251692 388476
rect 251916 388424 251968 388476
rect 249156 387812 249208 387864
rect 251456 387812 251508 387864
rect 151268 387744 151320 387796
rect 155132 387744 155184 387796
rect 220452 387744 220504 387796
rect 242348 387744 242400 387796
rect 116768 387676 116820 387728
rect 154948 387676 155000 387728
rect 220728 387676 220780 387728
rect 236736 387676 236788 387728
rect 137376 387608 137428 387660
rect 154764 387608 154816 387660
rect 220268 387608 220320 387660
rect 234436 387608 234488 387660
rect 145564 387540 145616 387592
rect 154856 387540 154908 387592
rect 112536 387472 112588 387524
rect 155040 387472 155092 387524
rect 147220 387064 147272 387116
rect 155500 387064 155552 387116
rect 151360 386316 151412 386368
rect 155040 386316 155092 386368
rect 220728 386316 220780 386368
rect 243820 386316 243872 386368
rect 131856 386248 131908 386300
rect 154672 386248 154724 386300
rect 220176 386248 220228 386300
rect 236828 386248 236880 386300
rect 148508 386180 148560 386232
rect 154856 386180 154908 386232
rect 220452 386180 220504 386232
rect 234528 386180 234580 386232
rect 127900 386112 127952 386164
rect 154948 386112 155000 386164
rect 126796 385636 126848 385688
rect 155224 385636 155276 385688
rect 112628 384956 112680 385008
rect 155132 384956 155184 385008
rect 220268 384956 220320 385008
rect 246764 384956 246816 385008
rect 116952 384888 117004 384940
rect 155040 384888 155092 384940
rect 220728 384888 220780 384940
rect 245200 384888 245252 384940
rect 143172 384820 143224 384872
rect 154948 384820 155000 384872
rect 220452 384820 220504 384872
rect 236920 384820 236972 384872
rect 147128 384752 147180 384804
rect 154856 384752 154908 384804
rect 220360 384752 220412 384804
rect 223120 384752 223172 384804
rect 148600 384684 148652 384736
rect 154672 384684 154724 384736
rect 227076 383664 227128 383716
rect 251180 383664 251232 383716
rect 220084 383596 220136 383648
rect 232872 383596 232924 383648
rect 131948 383528 132000 383580
rect 154856 383528 154908 383580
rect 138940 383460 138992 383512
rect 154948 383460 155000 383512
rect 149888 383392 149940 383444
rect 154672 383392 154724 383444
rect 124864 383324 124916 383376
rect 154948 383324 155000 383376
rect 220452 383256 220504 383308
rect 221924 383256 221976 383308
rect 234252 382236 234304 382288
rect 251180 382236 251232 382288
rect 114100 382168 114152 382220
rect 154948 382168 155000 382220
rect 220728 382168 220780 382220
rect 247960 382168 248012 382220
rect 117044 382100 117096 382152
rect 154580 382100 154632 382152
rect 220636 382100 220688 382152
rect 235448 382100 235500 382152
rect 139032 382032 139084 382084
rect 154856 382032 154908 382084
rect 220544 382032 220596 382084
rect 232964 382032 233016 382084
rect 144460 381964 144512 382016
rect 154948 381964 155000 382016
rect 112720 380808 112772 380860
rect 154948 380808 155000 380860
rect 220636 380808 220688 380860
rect 250720 380808 250772 380860
rect 118240 380740 118292 380792
rect 154764 380740 154816 380792
rect 220728 380740 220780 380792
rect 231492 380740 231544 380792
rect 126336 380672 126388 380724
rect 155040 380672 155092 380724
rect 219716 380672 219768 380724
rect 227444 380672 227496 380724
rect 132040 380604 132092 380656
rect 154856 380604 154908 380656
rect 143264 380536 143316 380588
rect 154948 380536 155000 380588
rect 220728 380468 220780 380520
rect 227352 380468 227404 380520
rect 220728 379448 220780 379500
rect 249524 379448 249576 379500
rect 120816 379380 120868 379432
rect 154856 379380 154908 379432
rect 220636 379380 220688 379432
rect 235816 379380 235868 379432
rect 124956 379312 125008 379364
rect 154948 379312 155000 379364
rect 220544 379312 220596 379364
rect 235540 379312 235592 379364
rect 147312 379244 147364 379296
rect 155040 379244 155092 379296
rect 118332 379176 118384 379228
rect 154948 379176 155000 379228
rect 139124 378768 139176 378820
rect 154672 378768 154724 378820
rect 220084 378156 220136 378208
rect 579804 378156 579856 378208
rect 112812 378088 112864 378140
rect 154948 378088 155000 378140
rect 220636 378088 220688 378140
rect 235724 378088 235776 378140
rect 119712 378020 119764 378072
rect 155040 378020 155092 378072
rect 220728 378020 220780 378072
rect 235632 378020 235684 378072
rect 120908 377952 120960 378004
rect 154764 377952 154816 378004
rect 220544 377952 220596 378004
rect 233056 377952 233108 378004
rect 140320 377884 140372 377936
rect 154856 377884 154908 377936
rect 144552 377816 144604 377868
rect 154948 377816 155000 377868
rect 114192 376660 114244 376712
rect 154948 376660 155000 376712
rect 220728 376660 220780 376712
rect 252008 376660 252060 376712
rect 121000 376592 121052 376644
rect 155040 376592 155092 376644
rect 219992 376592 220044 376644
rect 225788 376592 225840 376644
rect 125048 376524 125100 376576
rect 154856 376524 154908 376576
rect 145656 376456 145708 376508
rect 154948 376456 155000 376508
rect 143356 375980 143408 376032
rect 155132 375980 155184 376032
rect 219900 375980 219952 376032
rect 241152 375980 241204 376032
rect 219992 375844 220044 375896
rect 225880 375844 225932 375896
rect 112904 375300 112956 375352
rect 154580 375368 154632 375420
rect 154120 375300 154172 375352
rect 155040 375300 155092 375352
rect 220636 375300 220688 375352
rect 250812 375300 250864 375352
rect 117136 375232 117188 375284
rect 154948 375232 155000 375284
rect 220728 375232 220780 375284
rect 243912 375232 243964 375284
rect 141700 375164 141752 375216
rect 154856 375164 154908 375216
rect 219440 374824 219492 374876
rect 225972 374824 226024 374876
rect 118424 374620 118476 374672
rect 155592 374620 155644 374672
rect 125232 373940 125284 373992
rect 154672 373940 154724 373992
rect 220728 373940 220780 373992
rect 246856 373940 246908 373992
rect 126428 373872 126480 373924
rect 154764 373872 154816 373924
rect 220636 373872 220688 373924
rect 238392 373872 238444 373924
rect 129096 373804 129148 373856
rect 154580 373804 154632 373856
rect 220544 373804 220596 373856
rect 224408 373804 224460 373856
rect 141792 373736 141844 373788
rect 154948 373736 155000 373788
rect 147404 373668 147456 373720
rect 154856 373668 154908 373720
rect 114284 372512 114336 372564
rect 154764 372512 154816 372564
rect 219992 372512 220044 372564
rect 224776 372512 224828 372564
rect 121092 372444 121144 372496
rect 154948 372444 155000 372496
rect 140412 372376 140464 372428
rect 155132 372376 155184 372428
rect 140504 372308 140556 372360
rect 154948 372308 155000 372360
rect 220360 372308 220412 372360
rect 224500 372308 224552 372360
rect 148692 372240 148744 372292
rect 154856 372240 154908 372292
rect 220452 371968 220504 372020
rect 224592 371968 224644 372020
rect 218796 371832 218848 371884
rect 580448 371832 580500 371884
rect 3332 371220 3384 371272
rect 156696 371220 156748 371272
rect 115664 371152 115716 371204
rect 154764 371152 154816 371204
rect 220544 371152 220596 371204
rect 249616 371152 249668 371204
rect 127992 371084 128044 371136
rect 154672 371084 154724 371136
rect 220728 371084 220780 371136
rect 239772 371084 239824 371136
rect 133328 371016 133380 371068
rect 154948 371016 155000 371068
rect 220636 371016 220688 371068
rect 224684 371016 224736 371068
rect 135996 370948 136048 371000
rect 154856 370948 154908 371000
rect 141884 370880 141936 370932
rect 155132 370880 155184 370932
rect 219716 370472 219768 370524
rect 242440 370472 242492 370524
rect 220544 370132 220596 370184
rect 223304 370132 223356 370184
rect 114376 369792 114428 369844
rect 154672 369792 154724 369844
rect 115756 369724 115808 369776
rect 155132 369724 155184 369776
rect 119804 369656 119856 369708
rect 154948 369656 155000 369708
rect 121184 369588 121236 369640
rect 154856 369588 154908 369640
rect 220636 369588 220688 369640
rect 223212 369588 223264 369640
rect 148784 369520 148836 369572
rect 154764 369520 154816 369572
rect 220636 369316 220688 369368
rect 227536 369316 227588 369368
rect 219992 369112 220044 369164
rect 244096 369112 244148 369164
rect 151452 368432 151504 368484
rect 154580 368432 154632 368484
rect 220544 368432 220596 368484
rect 230112 368432 230164 368484
rect 129188 368364 129240 368416
rect 154764 368364 154816 368416
rect 220728 368364 220780 368416
rect 224868 368364 224920 368416
rect 140596 368296 140648 368348
rect 154948 368296 155000 368348
rect 122472 368228 122524 368280
rect 154856 368228 154908 368280
rect 219900 368024 219952 368076
rect 227628 368024 227680 368076
rect 150072 367820 150124 367872
rect 155316 367820 155368 367872
rect 118516 367752 118568 367804
rect 155408 367752 155460 367804
rect 219624 367752 219676 367804
rect 249708 367752 249760 367804
rect 126520 367004 126572 367056
rect 155132 367004 155184 367056
rect 220544 367004 220596 367056
rect 252192 367004 252244 367056
rect 128084 366936 128136 366988
rect 154948 366936 155000 366988
rect 220728 366936 220780 366988
rect 245292 366936 245344 366988
rect 137468 366868 137520 366920
rect 154672 366868 154724 366920
rect 220636 366868 220688 366920
rect 230204 366868 230256 366920
rect 144644 366800 144696 366852
rect 154856 366800 154908 366852
rect 124036 366324 124088 366376
rect 155224 366324 155276 366376
rect 219440 366324 219492 366376
rect 250904 366324 250956 366376
rect 151544 365644 151596 365696
rect 154948 365644 155000 365696
rect 220636 365644 220688 365696
rect 244004 365644 244056 365696
rect 133420 365576 133472 365628
rect 155132 365576 155184 365628
rect 219716 365576 219768 365628
rect 230296 365576 230348 365628
rect 134800 365508 134852 365560
rect 154856 365508 154908 365560
rect 137560 365440 137612 365492
rect 154672 365440 154724 365492
rect 112996 365372 113048 365424
rect 154764 365372 154816 365424
rect 231124 364352 231176 364404
rect 579988 364352 580040 364404
rect 123944 364284 123996 364336
rect 154764 364284 154816 364336
rect 220636 364284 220688 364336
rect 252100 364284 252152 364336
rect 126612 364216 126664 364268
rect 155040 364216 155092 364268
rect 220728 364216 220780 364268
rect 248052 364216 248104 364268
rect 128176 364148 128228 364200
rect 154856 364148 154908 364200
rect 220544 364148 220596 364200
rect 226064 364148 226116 364200
rect 129280 364080 129332 364132
rect 154948 364080 155000 364132
rect 113088 362856 113140 362908
rect 154580 362856 154632 362908
rect 114468 362788 114520 362840
rect 155040 362788 155092 362840
rect 220636 362788 220688 362840
rect 239864 362788 239916 362840
rect 143448 362720 143500 362772
rect 154856 362720 154908 362772
rect 220728 362720 220780 362772
rect 238484 362720 238536 362772
rect 145840 362652 145892 362704
rect 154948 362652 155000 362704
rect 220544 362652 220596 362704
rect 252284 362652 252336 362704
rect 122748 362176 122800 362228
rect 155408 362176 155460 362228
rect 220636 362176 220688 362228
rect 239956 362176 240008 362228
rect 220452 362108 220504 362160
rect 223396 362108 223448 362160
rect 115848 361496 115900 361548
rect 155040 361496 155092 361548
rect 220728 361496 220780 361548
rect 241244 361496 241296 361548
rect 129372 361428 129424 361480
rect 154764 361428 154816 361480
rect 132132 361360 132184 361412
rect 154856 361360 154908 361412
rect 133512 361292 133564 361344
rect 154580 361292 154632 361344
rect 136088 361224 136140 361276
rect 154948 361224 155000 361276
rect 219900 361088 219952 361140
rect 223488 361088 223540 361140
rect 220452 360884 220504 360936
rect 226892 360884 226944 360936
rect 220360 360816 220412 360868
rect 242624 360816 242676 360868
rect 122564 360136 122616 360188
rect 154580 360136 154632 360188
rect 220636 360136 220688 360188
rect 252376 360136 252428 360188
rect 126704 360068 126756 360120
rect 155040 360068 155092 360120
rect 219716 360068 219768 360120
rect 242532 360068 242584 360120
rect 128268 360000 128320 360052
rect 154948 360000 155000 360052
rect 220728 360000 220780 360052
rect 231584 360000 231636 360052
rect 141976 359932 142028 359984
rect 154856 359932 154908 359984
rect 147496 359864 147548 359916
rect 154948 359864 155000 359916
rect 219900 359456 219952 359508
rect 246212 359456 246264 359508
rect 220728 359252 220780 359304
rect 226800 359252 226852 359304
rect 152924 358708 152976 358760
rect 155592 358708 155644 358760
rect 220636 358708 220688 358760
rect 231676 358708 231728 358760
rect 117228 358640 117280 358692
rect 154948 358640 155000 358692
rect 219992 358640 220044 358692
rect 228640 358640 228692 358692
rect 137652 358572 137704 358624
rect 154764 358572 154816 358624
rect 115112 358504 115164 358556
rect 154580 358504 154632 358556
rect 220544 358028 220596 358080
rect 238576 358028 238628 358080
rect 2964 357416 3016 357468
rect 156788 357416 156840 357468
rect 151636 357348 151688 357400
rect 155040 357348 155092 357400
rect 220728 357348 220780 357400
rect 231768 357348 231820 357400
rect 126888 357280 126940 357332
rect 154764 357280 154816 357332
rect 132224 357212 132276 357264
rect 154948 357212 155000 357264
rect 220636 357212 220688 357264
rect 222016 357212 222068 357264
rect 149980 357144 150032 357196
rect 154856 357144 154908 357196
rect 125140 357076 125192 357128
rect 154948 357076 155000 357128
rect 219900 356668 219952 356720
rect 248972 356668 249024 356720
rect 153016 355988 153068 356040
rect 154580 355988 154632 356040
rect 220728 355988 220780 356040
rect 246948 355988 247000 356040
rect 137744 355920 137796 355972
rect 155040 355920 155092 355972
rect 144736 355852 144788 355904
rect 154856 355852 154908 355904
rect 119896 355784 119948 355836
rect 154948 355784 155000 355836
rect 219808 355784 219860 355836
rect 224132 355784 224184 355836
rect 220728 355716 220780 355768
rect 226156 355716 226208 355768
rect 130936 355376 130988 355428
rect 155592 355376 155644 355428
rect 119252 355308 119304 355360
rect 155132 355308 155184 355360
rect 112260 354628 112312 354680
rect 154856 354628 154908 354680
rect 220728 354628 220780 354680
rect 245384 354628 245436 354680
rect 112352 354560 112404 354612
rect 154580 354560 154632 354612
rect 116400 354492 116452 354544
rect 154948 354492 155000 354544
rect 133604 354424 133656 354476
rect 154764 354424 154816 354476
rect 220636 354356 220688 354408
rect 228732 354356 228784 354408
rect 220636 353948 220688 354000
rect 251088 353948 251140 354000
rect 115020 353200 115072 353252
rect 154764 353200 154816 353252
rect 220728 353200 220780 353252
rect 245476 353200 245528 353252
rect 132408 353132 132460 353184
rect 154948 353132 155000 353184
rect 132316 353064 132368 353116
rect 154856 353064 154908 353116
rect 139216 352996 139268 353048
rect 155040 352996 155092 353048
rect 142068 352928 142120 352980
rect 154856 352928 154908 352980
rect 220452 352724 220504 352776
rect 228824 352724 228876 352776
rect 220452 352452 220504 352504
rect 222752 352452 222804 352504
rect 258724 351908 258776 351960
rect 580172 351908 580224 351960
rect 119988 351840 120040 351892
rect 154856 351840 154908 351892
rect 220728 351840 220780 351892
rect 250996 351840 251048 351892
rect 124128 351772 124180 351824
rect 154948 351772 155000 351824
rect 145932 351704 145984 351756
rect 155040 351704 155092 351756
rect 148876 351636 148928 351688
rect 154764 351636 154816 351688
rect 219992 351296 220044 351348
rect 228916 351296 228968 351348
rect 219900 351024 219952 351076
rect 226248 351024 226300 351076
rect 116492 350480 116544 350532
rect 154580 350480 154632 350532
rect 220544 350480 220596 350532
rect 244188 350480 244240 350532
rect 140688 350412 140740 350464
rect 154948 350412 155000 350464
rect 219900 350208 219952 350260
rect 229008 350208 229060 350260
rect 220728 349800 220780 349852
rect 245568 349800 245620 349852
rect 138756 349188 138808 349240
rect 154948 349188 155000 349240
rect 126244 349120 126296 349172
rect 154856 349120 154908 349172
rect 220636 349052 220688 349104
rect 248144 349052 248196 349104
rect 220544 348984 220596 349036
rect 224040 348984 224092 349036
rect 220544 348372 220596 348424
rect 236644 348372 236696 348424
rect 220452 348032 220504 348084
rect 223948 348032 224000 348084
rect 122656 347964 122708 348016
rect 154856 347964 154908 348016
rect 119436 347896 119488 347948
rect 154948 347896 155000 347948
rect 119528 347828 119580 347880
rect 154764 347828 154816 347880
rect 116676 347760 116728 347812
rect 155040 347760 155092 347812
rect 220452 347692 220504 347744
rect 234160 347692 234212 347744
rect 220728 347624 220780 347676
rect 233976 347624 234028 347676
rect 220636 347556 220688 347608
rect 231032 347556 231084 347608
rect 118240 347012 118292 347064
rect 154948 347012 155000 347064
rect 142988 346604 143040 346656
rect 154856 346604 154908 346656
rect 136180 346536 136232 346588
rect 154948 346536 155000 346588
rect 116584 346468 116636 346520
rect 155040 346468 155092 346520
rect 113916 346400 113968 346452
rect 154580 346400 154632 346452
rect 220636 346332 220688 346384
rect 252468 346332 252520 346384
rect 220728 346264 220780 346316
rect 229744 346264 229796 346316
rect 220728 345924 220780 345976
rect 222108 345924 222160 345976
rect 122104 345652 122156 345704
rect 154856 345652 154908 345704
rect 141516 345176 141568 345228
rect 154948 345176 155000 345228
rect 113824 345108 113876 345160
rect 155040 345108 155092 345160
rect 3056 345040 3108 345092
rect 135996 345040 136048 345092
rect 140136 345040 140188 345092
rect 154948 345040 155000 345092
rect 220636 344972 220688 345024
rect 250444 344972 250496 345024
rect 220728 344904 220780 344956
rect 231216 344904 231268 344956
rect 219900 343884 219952 343936
rect 226984 343884 227036 343936
rect 131764 343816 131816 343868
rect 154580 343816 154632 343868
rect 123484 343748 123536 343800
rect 154948 343748 155000 343800
rect 120724 343680 120776 343732
rect 155040 343680 155092 343732
rect 119344 343612 119396 343664
rect 154856 343612 154908 343664
rect 220728 343544 220780 343596
rect 247776 343544 247828 343596
rect 220636 343340 220688 343392
rect 222844 343340 222896 343392
rect 115204 342864 115256 342916
rect 154580 342864 154632 342916
rect 220452 342524 220504 342576
rect 221740 342524 221792 342576
rect 144552 342388 144604 342440
rect 154856 342388 154908 342440
rect 139216 342320 139268 342372
rect 154948 342320 155000 342372
rect 115848 342252 115900 342304
rect 155040 342252 155092 342304
rect 220728 342116 220780 342168
rect 251916 342116 251968 342168
rect 219808 341912 219860 341964
rect 221648 341912 221700 341964
rect 128176 341096 128228 341148
rect 154948 341096 155000 341148
rect 124036 341028 124088 341080
rect 154764 341028 154816 341080
rect 121184 340960 121236 341012
rect 155040 340960 155092 341012
rect 117136 340892 117188 340944
rect 154856 340892 154908 340944
rect 219532 340824 219584 340876
rect 249156 340824 249208 340876
rect 219900 340484 219952 340536
rect 227076 340484 227128 340536
rect 155316 340144 155368 340196
rect 155592 340144 155644 340196
rect 147496 339736 147548 339788
rect 154948 339736 155000 339788
rect 141792 339668 141844 339720
rect 154856 339668 154908 339720
rect 137284 339600 137336 339652
rect 155040 339600 155092 339652
rect 134708 339532 134760 339584
rect 154948 339532 155000 339584
rect 133236 339464 133288 339516
rect 154764 339464 154816 339516
rect 220728 339396 220780 339448
rect 251732 339396 251784 339448
rect 220636 339328 220688 339380
rect 251640 339328 251692 339380
rect 220452 339260 220504 339312
rect 234252 339260 234304 339312
rect 117228 338716 117280 338768
rect 154580 338716 154632 338768
rect 148876 338308 148928 338360
rect 154948 338308 155000 338360
rect 144736 338240 144788 338292
rect 154856 338240 154908 338292
rect 126796 338172 126848 338224
rect 154672 338172 154724 338224
rect 125140 338104 125192 338156
rect 155040 338104 155092 338156
rect 119896 337356 119948 337408
rect 155132 337356 155184 337408
rect 112260 337016 112312 337068
rect 154580 337016 154632 337068
rect 143356 336948 143408 337000
rect 154856 336948 154908 337000
rect 139124 336880 139176 336932
rect 154764 336880 154816 336932
rect 220544 336880 220596 336932
rect 227076 336880 227128 336932
rect 133604 336812 133656 336864
rect 154948 336812 155000 336864
rect 220728 336812 220780 336864
rect 233976 336812 234028 336864
rect 151544 336744 151596 336796
rect 155040 336744 155092 336796
rect 220636 336744 220688 336796
rect 247776 336744 247828 336796
rect 220636 336064 220688 336116
rect 223948 336064 224000 336116
rect 119804 335588 119856 335640
rect 154764 335588 154816 335640
rect 145932 335520 145984 335572
rect 155040 335520 155092 335572
rect 220728 335520 220780 335572
rect 222936 335520 222988 335572
rect 133512 335452 133564 335504
rect 154856 335452 154908 335504
rect 220544 335452 220596 335504
rect 246580 335452 246632 335504
rect 128084 335384 128136 335436
rect 154672 335384 154724 335436
rect 151452 335316 151504 335368
rect 154948 335316 155000 335368
rect 155224 335316 155276 335368
rect 155684 335316 155736 335368
rect 140596 334636 140648 334688
rect 155040 334636 155092 334688
rect 115112 334568 115164 334620
rect 155500 334568 155552 334620
rect 219900 334568 219952 334620
rect 229836 334568 229888 334620
rect 132224 334092 132276 334144
rect 154948 334092 155000 334144
rect 148784 334024 148836 334076
rect 154764 334024 154816 334076
rect 219992 334024 220044 334076
rect 222844 334024 222896 334076
rect 153016 333956 153068 334008
rect 155132 333956 155184 334008
rect 220360 333956 220412 334008
rect 249616 333956 249668 334008
rect 117964 333208 118016 333260
rect 155408 333208 155460 333260
rect 219808 333072 219860 333124
rect 227720 333072 227772 333124
rect 114468 332868 114520 332920
rect 154764 332868 154816 332920
rect 145840 332800 145892 332852
rect 154580 332800 154632 332852
rect 140504 332732 140556 332784
rect 154948 332732 155000 332784
rect 129372 332664 129424 332716
rect 154856 332664 154908 332716
rect 220636 332664 220688 332716
rect 235632 332664 235684 332716
rect 220728 332596 220780 332648
rect 244924 332596 244976 332648
rect 220452 331848 220504 331900
rect 248144 331848 248196 331900
rect 219900 331576 219952 331628
rect 227536 331576 227588 331628
rect 150072 331440 150124 331492
rect 154948 331440 155000 331492
rect 219900 331440 219952 331492
rect 224132 331440 224184 331492
rect 132132 331372 132184 331424
rect 154856 331372 154908 331424
rect 129280 331304 129332 331356
rect 154948 331304 155000 331356
rect 115756 331236 115808 331288
rect 155040 331236 155092 331288
rect 220544 331236 220596 331288
rect 254952 331236 255004 331288
rect 147404 330488 147456 330540
rect 154764 330488 154816 330540
rect 144644 330012 144696 330064
rect 154948 330012 155000 330064
rect 137652 329944 137704 329996
rect 154856 329944 154908 329996
rect 219716 329944 219768 329996
rect 228916 329944 228968 329996
rect 122564 329876 122616 329928
rect 155040 329876 155092 329928
rect 220544 329876 220596 329928
rect 231676 329876 231728 329928
rect 115664 329808 115716 329860
rect 155132 329808 155184 329860
rect 220728 329808 220780 329860
rect 250444 329808 250496 329860
rect 220636 329060 220688 329112
rect 241244 329060 241296 329112
rect 219532 328992 219584 329044
rect 224868 328992 224920 329044
rect 152924 328720 152976 328772
rect 154580 328720 154632 328772
rect 149980 328652 150032 328704
rect 154948 328652 155000 328704
rect 140412 328584 140464 328636
rect 154856 328584 154908 328636
rect 132040 328516 132092 328568
rect 154580 328516 154632 328568
rect 220728 328516 220780 328568
rect 231584 328516 231636 328568
rect 112352 328448 112404 328500
rect 155040 328448 155092 328500
rect 220544 328448 220596 328500
rect 255964 328448 256016 328500
rect 220268 327904 220320 327956
rect 228824 327904 228876 327956
rect 3424 327700 3476 327752
rect 158260 327700 158312 327752
rect 227720 327700 227772 327752
rect 257344 327700 257396 327752
rect 143264 327292 143316 327344
rect 154764 327292 154816 327344
rect 121092 327224 121144 327276
rect 154948 327224 155000 327276
rect 118056 327156 118108 327208
rect 154856 327156 154908 327208
rect 220268 327156 220320 327208
rect 226064 327156 226116 327208
rect 117044 327088 117096 327140
rect 155040 327088 155092 327140
rect 220728 327088 220780 327140
rect 238300 327088 238352 327140
rect 113088 325932 113140 325984
rect 154856 325932 154908 325984
rect 137560 325864 137612 325916
rect 154948 325864 155000 325916
rect 220360 325864 220412 325916
rect 224776 325864 224828 325916
rect 131948 325796 132000 325848
rect 154580 325796 154632 325848
rect 112996 325728 113048 325780
rect 154764 325728 154816 325780
rect 220728 325728 220780 325780
rect 228732 325728 228784 325780
rect 151360 325660 151412 325712
rect 155040 325660 155092 325712
rect 220636 325660 220688 325712
rect 236920 325660 236972 325712
rect 3516 324912 3568 324964
rect 140044 324912 140096 324964
rect 219532 324912 219584 324964
rect 234344 324912 234396 324964
rect 112904 324572 112956 324624
rect 154948 324572 155000 324624
rect 220728 324572 220780 324624
rect 123944 324504 123996 324556
rect 155040 324504 155092 324556
rect 122472 324436 122524 324488
rect 154856 324436 154908 324488
rect 220268 324436 220320 324488
rect 225972 324436 226024 324488
rect 121000 324368 121052 324420
rect 154764 324368 154816 324420
rect 220360 324368 220412 324420
rect 149888 324300 149940 324352
rect 154948 324300 155000 324352
rect 219900 324300 219952 324352
rect 224684 324300 224736 324352
rect 235540 324368 235592 324420
rect 580172 324300 580224 324352
rect 3608 323552 3660 323604
rect 157892 323552 157944 323604
rect 219716 323280 219768 323332
rect 228640 323280 228692 323332
rect 112812 323212 112864 323264
rect 154948 323212 155000 323264
rect 137468 323144 137520 323196
rect 155040 323144 155092 323196
rect 130844 323076 130896 323128
rect 154948 323076 155000 323128
rect 220268 323076 220320 323128
rect 224592 323076 224644 323128
rect 114376 323008 114428 323060
rect 154856 323008 154908 323060
rect 220728 323008 220780 323060
rect 224040 323008 224092 323060
rect 220636 322940 220688 322992
rect 231492 322940 231544 322992
rect 3792 322260 3844 322312
rect 142896 322260 142948 322312
rect 3700 322192 3752 322244
rect 152556 322192 152608 322244
rect 147312 321784 147364 321836
rect 154856 321784 154908 321836
rect 126704 321716 126756 321768
rect 155040 321716 155092 321768
rect 220544 321716 220596 321768
rect 236828 321716 236880 321768
rect 116952 321648 117004 321700
rect 154948 321648 155000 321700
rect 220728 321648 220780 321700
rect 250720 321648 250772 321700
rect 115572 321580 115624 321632
rect 154764 321580 154816 321632
rect 220636 321580 220688 321632
rect 256332 321580 256384 321632
rect 228364 320900 228416 320952
rect 580908 320900 580960 320952
rect 218980 320832 219032 320884
rect 580724 320832 580776 320884
rect 220268 320560 220320 320612
rect 222752 320560 222804 320612
rect 144460 320424 144512 320476
rect 154948 320424 155000 320476
rect 143172 320356 143224 320408
rect 154856 320356 154908 320408
rect 133420 320288 133472 320340
rect 154764 320288 154816 320340
rect 133328 320220 133380 320272
rect 154948 320220 155000 320272
rect 220268 320220 220320 320272
rect 242348 320220 242400 320272
rect 112720 320152 112772 320204
rect 155040 320152 155092 320204
rect 220728 320152 220780 320204
rect 249524 320152 249576 320204
rect 220176 320016 220228 320068
rect 220268 319812 220320 319864
rect 220452 319744 220504 319796
rect 223488 319744 223540 319796
rect 229928 319676 229980 319728
rect 580356 319676 580408 319728
rect 229744 319608 229796 319660
rect 580264 319608 580316 319660
rect 226984 319540 227036 319592
rect 580540 319540 580592 319592
rect 221648 319472 221700 319524
rect 580816 319472 580868 319524
rect 118148 319404 118200 319456
rect 154672 319404 154724 319456
rect 219164 319404 219216 319456
rect 580632 319404 580684 319456
rect 148692 318996 148744 319048
rect 154856 318996 154908 319048
rect 220728 318996 220780 319048
rect 252008 318996 252060 319048
rect 130752 318928 130804 318980
rect 154764 318928 154816 318980
rect 127992 318860 128044 318912
rect 154948 318860 155000 318912
rect 220452 318860 220504 318912
rect 223396 318860 223448 318912
rect 3424 318792 3476 318844
rect 30012 318792 30064 318844
rect 114284 318792 114336 318844
rect 155040 318792 155092 318844
rect 220360 318792 220412 318844
rect 223304 318792 223356 318844
rect 254584 318792 254636 318844
rect 580448 318792 580500 318844
rect 219992 318384 220044 318436
rect 221832 318384 221884 318436
rect 122380 318044 122432 318096
rect 154580 318044 154632 318096
rect 148600 317704 148652 317756
rect 154856 317704 154908 317756
rect 145656 317636 145708 317688
rect 154948 317636 155000 317688
rect 139032 317568 139084 317620
rect 155040 317568 155092 317620
rect 122288 317500 122340 317552
rect 154764 317500 154816 317552
rect 220636 317500 220688 317552
rect 239680 317500 239732 317552
rect 119712 317432 119764 317484
rect 154672 317432 154724 317484
rect 220728 317432 220780 317484
rect 256240 317432 256292 317484
rect 220636 316480 220688 316532
rect 225880 316480 225932 316532
rect 152832 316344 152884 316396
rect 154580 316344 154632 316396
rect 115480 316276 115532 316328
rect 154856 316276 154908 316328
rect 147220 316208 147272 316260
rect 154764 316208 154816 316260
rect 130660 316140 130712 316192
rect 155040 316140 155092 316192
rect 126612 316072 126664 316124
rect 154948 316072 155000 316124
rect 220452 316072 220504 316124
rect 248052 316072 248104 316124
rect 220728 316004 220780 316056
rect 254860 316004 254912 316056
rect 127900 314848 127952 314900
rect 155040 314848 155092 314900
rect 219992 314848 220044 314900
rect 227352 314848 227404 314900
rect 125048 314780 125100 314832
rect 154856 314780 154908 314832
rect 220544 314780 220596 314832
rect 223212 314780 223264 314832
rect 123852 314712 123904 314764
rect 154764 314712 154816 314764
rect 220636 314712 220688 314764
rect 230204 314712 230256 314764
rect 122196 314644 122248 314696
rect 154948 314644 155000 314696
rect 220728 314644 220780 314696
rect 243912 314644 243964 314696
rect 111800 314576 111852 314628
rect 138756 314576 138808 314628
rect 147128 313556 147180 313608
rect 154948 313556 155000 313608
rect 134616 313488 134668 313540
rect 154580 313488 154632 313540
rect 130568 313420 130620 313472
rect 154948 313420 155000 313472
rect 220728 313420 220780 313472
rect 230112 313420 230164 313472
rect 115388 313352 115440 313404
rect 154856 313352 154908 313404
rect 220452 313352 220504 313404
rect 239588 313352 239640 313404
rect 112628 313284 112680 313336
rect 154764 313284 154816 313336
rect 220636 313284 220688 313336
rect 249432 313284 249484 313336
rect 111800 313216 111852 313268
rect 126244 313216 126296 313268
rect 111892 313148 111944 313200
rect 117964 313148 118016 313200
rect 227076 312536 227128 312588
rect 257712 312536 257764 312588
rect 220452 312400 220504 312452
rect 224500 312400 224552 312452
rect 219900 312196 219952 312248
rect 227260 312196 227312 312248
rect 123760 312128 123812 312180
rect 154948 312128 155000 312180
rect 133144 312060 133196 312112
rect 154580 312060 154632 312112
rect 127808 311992 127860 312044
rect 154764 311992 154816 312044
rect 126520 311924 126572 311976
rect 154856 311924 154908 311976
rect 220728 311924 220780 311976
rect 225788 311924 225840 311976
rect 152740 311856 152792 311908
rect 154580 311856 154632 311908
rect 220452 311856 220504 311908
rect 235448 311856 235500 311908
rect 111892 311788 111944 311840
rect 122656 311788 122708 311840
rect 229836 311788 229888 311840
rect 256700 311788 256752 311840
rect 111800 311720 111852 311772
rect 116676 311720 116728 311772
rect 154672 311176 154724 311228
rect 155408 311176 155460 311228
rect 116860 311108 116912 311160
rect 155592 311108 155644 311160
rect 114192 310768 114244 310820
rect 154856 310768 154908 310820
rect 145748 310700 145800 310752
rect 154948 310700 155000 310752
rect 138940 310632 138992 310684
rect 154856 310632 154908 310684
rect 220544 310632 220596 310684
rect 227444 310632 227496 310684
rect 119620 310564 119672 310616
rect 154764 310564 154816 310616
rect 220728 310564 220780 310616
rect 230020 310564 230072 310616
rect 151268 310496 151320 310548
rect 155040 310496 155092 310548
rect 220636 310496 220688 310548
rect 245108 310496 245160 310548
rect 111800 310428 111852 310480
rect 119528 310428 119580 310480
rect 111892 310360 111944 310412
rect 119436 310360 119488 310412
rect 233976 309748 234028 309800
rect 256792 309748 256844 309800
rect 144368 309408 144420 309460
rect 154856 309408 154908 309460
rect 220636 309408 220688 309460
rect 224408 309408 224460 309460
rect 130476 309340 130528 309392
rect 154764 309340 154816 309392
rect 127716 309272 127768 309324
rect 154948 309272 155000 309324
rect 126428 309204 126480 309256
rect 154580 309204 154632 309256
rect 220544 309204 220596 309256
rect 234252 309204 234304 309256
rect 124956 309136 125008 309188
rect 154948 309136 155000 309188
rect 220728 309136 220780 309188
rect 246764 309136 246816 309188
rect 111800 309068 111852 309120
rect 118240 309068 118292 309120
rect 247776 309068 247828 309120
rect 256700 309068 256752 309120
rect 111892 309000 111944 309052
rect 116584 309000 116636 309052
rect 149796 307980 149848 308032
rect 154948 307980 155000 308032
rect 219900 307980 219952 308032
rect 225696 307980 225748 308032
rect 141700 307912 141752 307964
rect 154764 307912 154816 307964
rect 220728 307912 220780 307964
rect 232688 307912 232740 307964
rect 123576 307844 123628 307896
rect 155040 307844 155092 307896
rect 220636 307844 220688 307896
rect 238208 307844 238260 307896
rect 117964 307776 118016 307828
rect 154856 307776 154908 307828
rect 219716 307776 219768 307828
rect 242256 307776 242308 307828
rect 111800 307708 111852 307760
rect 142988 307708 143040 307760
rect 111800 307504 111852 307556
rect 113916 307504 113968 307556
rect 148508 306620 148560 306672
rect 155040 306620 155092 306672
rect 143080 306552 143132 306604
rect 154948 306552 155000 306604
rect 130384 306484 130436 306536
rect 154856 306484 154908 306536
rect 155040 306484 155092 306536
rect 155684 306484 155736 306536
rect 220544 306484 220596 306536
rect 232872 306484 232924 306536
rect 126336 306416 126388 306468
rect 154948 306416 155000 306468
rect 155316 306416 155368 306468
rect 220728 306416 220780 306468
rect 238116 306416 238168 306468
rect 112076 306348 112128 306400
rect 154764 306348 154816 306400
rect 154856 306348 154908 306400
rect 220636 306348 220688 306400
rect 247960 306348 248012 306400
rect 111800 306280 111852 306332
rect 136180 306280 136232 306332
rect 111892 306212 111944 306264
rect 122104 306212 122156 306264
rect 136088 305600 136140 305652
rect 155500 305600 155552 305652
rect 244924 305600 244976 305652
rect 257620 305600 257672 305652
rect 154580 305532 154632 305584
rect 155684 305532 155736 305584
rect 154948 305464 155000 305516
rect 155316 305464 155368 305516
rect 220728 305328 220780 305380
rect 224316 305328 224368 305380
rect 155132 305192 155184 305244
rect 155408 305192 155460 305244
rect 127624 305124 127676 305176
rect 154856 305124 154908 305176
rect 220728 305124 220780 305176
rect 243820 305124 243872 305176
rect 124864 305056 124916 305108
rect 154764 305056 154816 305108
rect 220636 305056 220688 305108
rect 245016 305056 245068 305108
rect 3240 304988 3292 305040
rect 30104 304988 30156 305040
rect 114100 304988 114152 305040
rect 154948 304988 155000 305040
rect 220544 304988 220596 305040
rect 246672 304988 246724 305040
rect 111892 304920 111944 304972
rect 141516 304920 141568 304972
rect 111800 304852 111852 304904
rect 113824 304852 113876 304904
rect 112076 304444 112128 304496
rect 112536 304444 112588 304496
rect 119528 304240 119580 304292
rect 155132 304240 155184 304292
rect 115296 303832 115348 303884
rect 154948 303832 155000 303884
rect 140320 303764 140372 303816
rect 154580 303764 154632 303816
rect 220636 303764 220688 303816
rect 231400 303764 231452 303816
rect 116768 303696 116820 303748
rect 154856 303696 154908 303748
rect 220728 303696 220780 303748
rect 239496 303696 239548 303748
rect 152648 303628 152700 303680
rect 155500 303628 155552 303680
rect 220452 303628 220504 303680
rect 250628 303628 250680 303680
rect 111892 303560 111944 303612
rect 155316 303560 155368 303612
rect 223948 303560 224000 303612
rect 256700 303560 256752 303612
rect 111800 303492 111852 303544
rect 117228 303492 117280 303544
rect 141608 302880 141660 302932
rect 154764 302880 154816 302932
rect 114008 302472 114060 302524
rect 154948 302472 155000 302524
rect 138756 302404 138808 302456
rect 154672 302404 154724 302456
rect 129188 302336 129240 302388
rect 155132 302336 155184 302388
rect 219900 302336 219952 302388
rect 224224 302336 224276 302388
rect 126244 302268 126296 302320
rect 154856 302268 154908 302320
rect 220544 302268 220596 302320
rect 241152 302268 241204 302320
rect 220728 302200 220780 302252
rect 241060 302200 241112 302252
rect 111800 302132 111852 302184
rect 140136 302132 140188 302184
rect 111892 302064 111944 302116
rect 120724 302064 120776 302116
rect 154120 301384 154172 301436
rect 154580 301384 154632 301436
rect 140228 301044 140280 301096
rect 154580 301044 154632 301096
rect 219992 301044 220044 301096
rect 232596 301044 232648 301096
rect 137376 300976 137428 301028
rect 154856 300976 154908 301028
rect 220728 300976 220780 301028
rect 233976 300976 234028 301028
rect 120816 300908 120868 300960
rect 154764 300908 154816 300960
rect 220544 300908 220596 300960
rect 234160 300908 234212 300960
rect 119436 300840 119488 300892
rect 154672 300840 154724 300892
rect 220636 300840 220688 300892
rect 256148 300840 256200 300892
rect 111984 300772 112036 300824
rect 131764 300772 131816 300824
rect 246580 300772 246632 300824
rect 256700 300772 256752 300824
rect 111892 300704 111944 300756
rect 123484 300704 123536 300756
rect 111800 300636 111852 300688
rect 119344 300636 119396 300688
rect 142988 299684 143040 299736
rect 154672 299684 154724 299736
rect 141516 299616 141568 299668
rect 154580 299616 154632 299668
rect 131856 299548 131908 299600
rect 154764 299548 154816 299600
rect 220636 299548 220688 299600
rect 236644 299548 236696 299600
rect 113916 299480 113968 299532
rect 154856 299480 154908 299532
rect 220728 299480 220780 299532
rect 251916 299480 251968 299532
rect 222936 299412 222988 299464
rect 256700 299412 256752 299464
rect 111800 299140 111852 299192
rect 115204 299140 115256 299192
rect 111800 298800 111852 298852
rect 115848 298800 115900 298852
rect 123668 298732 123720 298784
rect 155500 298732 155552 298784
rect 148416 298324 148468 298376
rect 154948 298324 155000 298376
rect 149704 298256 149756 298308
rect 154856 298256 154908 298308
rect 219992 298256 220044 298308
rect 223120 298256 223172 298308
rect 144276 298188 144328 298240
rect 154580 298188 154632 298240
rect 220544 298188 220596 298240
rect 231308 298188 231360 298240
rect 123484 298120 123536 298172
rect 154764 298120 154816 298172
rect 220728 298120 220780 298172
rect 254768 298120 254820 298172
rect 111892 298052 111944 298104
rect 144552 298052 144604 298104
rect 111800 297916 111852 297968
rect 115112 297916 115164 297968
rect 220728 297576 220780 297628
rect 223028 297576 223080 297628
rect 147036 297372 147088 297424
rect 154672 297372 154724 297424
rect 151636 297168 151688 297220
rect 155408 297168 155460 297220
rect 138848 296828 138900 296880
rect 154580 296828 154632 296880
rect 116676 296760 116728 296812
rect 154764 296760 154816 296812
rect 220728 296760 220780 296812
rect 246580 296760 246632 296812
rect 115204 296692 115256 296744
rect 154948 296692 155000 296744
rect 220636 296692 220688 296744
rect 247868 296692 247920 296744
rect 111800 296624 111852 296676
rect 155224 296624 155276 296676
rect 220268 296624 220320 296676
rect 256700 296624 256752 296676
rect 111892 296556 111944 296608
rect 139216 296556 139268 296608
rect 145564 295604 145616 295656
rect 154580 295604 154632 295656
rect 131764 295536 131816 295588
rect 154856 295536 154908 295588
rect 129096 295468 129148 295520
rect 154764 295468 154816 295520
rect 219900 295468 219952 295520
rect 228548 295468 228600 295520
rect 129004 295400 129056 295452
rect 154672 295400 154724 295452
rect 220636 295400 220688 295452
rect 231216 295400 231268 295452
rect 113824 295332 113876 295384
rect 154948 295332 155000 295384
rect 220728 295332 220780 295384
rect 256056 295332 256108 295384
rect 111892 295264 111944 295316
rect 128176 295264 128228 295316
rect 222844 295264 222896 295316
rect 256700 295264 256752 295316
rect 111800 295196 111852 295248
rect 124036 295196 124088 295248
rect 151176 294244 151228 294296
rect 154856 294244 154908 294296
rect 140136 294176 140188 294228
rect 154672 294176 154724 294228
rect 220268 294176 220320 294228
rect 225604 294176 225656 294228
rect 122104 294108 122156 294160
rect 154580 294108 154632 294160
rect 220728 294108 220780 294160
rect 254676 294108 254728 294160
rect 120908 294040 120960 294092
rect 154764 294040 154816 294092
rect 112444 293972 112496 294024
rect 154580 293972 154632 294024
rect 219900 293972 219952 294024
rect 222936 293972 222988 294024
rect 111800 293904 111852 293956
rect 121184 293904 121236 293956
rect 111892 293836 111944 293888
rect 117136 293836 117188 293888
rect 250444 292748 250496 292800
rect 257436 292748 257488 292800
rect 120724 292680 120776 292732
rect 154580 292680 154632 292732
rect 220544 292680 220596 292732
rect 228456 292680 228508 292732
rect 119344 292612 119396 292664
rect 154672 292612 154724 292664
rect 154948 292612 155000 292664
rect 155316 292612 155368 292664
rect 220728 292612 220780 292664
rect 243728 292612 243780 292664
rect 116584 292544 116636 292596
rect 154580 292544 154632 292596
rect 220636 292544 220688 292596
rect 249340 292544 249392 292596
rect 111892 292476 111944 292528
rect 137284 292476 137336 292528
rect 249616 292476 249668 292528
rect 256700 292476 256752 292528
rect 111800 292408 111852 292460
rect 119896 292408 119948 292460
rect 144552 291796 144604 291848
rect 155132 291796 155184 291848
rect 219900 291320 219952 291372
rect 227168 291320 227220 291372
rect 220636 291252 220688 291304
rect 249156 291252 249208 291304
rect 220728 291184 220780 291236
rect 250536 291184 250588 291236
rect 111892 291116 111944 291168
rect 147496 291116 147548 291168
rect 248144 291116 248196 291168
rect 256700 291116 256752 291168
rect 111800 291048 111852 291100
rect 133236 291048 133288 291100
rect 137284 290436 137336 290488
rect 154672 290436 154724 290488
rect 220728 289960 220780 290012
rect 235356 289960 235408 290012
rect 220636 289892 220688 289944
rect 244924 289892 244976 289944
rect 220728 289824 220780 289876
rect 247776 289824 247828 289876
rect 111800 289756 111852 289808
rect 141792 289756 141844 289808
rect 255964 289756 256016 289808
rect 257804 289756 257856 289808
rect 111892 289688 111944 289740
rect 134708 289688 134760 289740
rect 220544 288532 220596 288584
rect 229836 288532 229888 288584
rect 220636 288464 220688 288516
rect 236736 288464 236788 288516
rect 220728 288396 220780 288448
rect 250444 288396 250496 288448
rect 111892 288328 111944 288380
rect 144736 288328 144788 288380
rect 235632 288328 235684 288380
rect 256700 288328 256752 288380
rect 111800 288260 111852 288312
rect 126796 288260 126848 288312
rect 220728 287376 220780 287428
rect 227076 287376 227128 287428
rect 220636 287104 220688 287156
rect 235264 287104 235316 287156
rect 219532 287036 219584 287088
rect 242164 287036 242216 287088
rect 111892 286968 111944 287020
rect 148876 286968 148928 287020
rect 111800 286900 111852 286952
rect 125140 286900 125192 286952
rect 219900 286696 219952 286748
rect 222844 286696 222896 286748
rect 219900 286084 219952 286136
rect 221740 286084 221792 286136
rect 220728 285880 220780 285932
rect 255964 285880 256016 285932
rect 220636 285744 220688 285796
rect 232780 285744 232832 285796
rect 111800 285608 111852 285660
rect 140596 285608 140648 285660
rect 111892 285540 111944 285592
rect 139124 285540 139176 285592
rect 111892 284248 111944 284300
rect 151544 284248 151596 284300
rect 111800 284180 111852 284232
rect 143356 284180 143408 284232
rect 224040 283568 224092 283620
rect 257344 283568 257396 283620
rect 111800 282820 111852 282872
rect 133604 282820 133656 282872
rect 227536 282820 227588 282872
rect 256700 282820 256752 282872
rect 133236 282140 133288 282192
rect 154948 282140 155000 282192
rect 111892 281460 111944 281512
rect 128084 281460 128136 281512
rect 111800 281392 111852 281444
rect 119804 281392 119856 281444
rect 111800 280100 111852 280152
rect 145932 280100 145984 280152
rect 254952 280100 255004 280152
rect 256700 280100 256752 280152
rect 111892 280032 111944 280084
rect 133512 280032 133564 280084
rect 111892 278672 111944 278724
rect 154120 278672 154172 278724
rect 224132 278672 224184 278724
rect 256700 278672 256752 278724
rect 111800 278604 111852 278656
rect 151452 278604 151504 278656
rect 111800 277312 111852 277364
rect 155868 277312 155920 277364
rect 111892 277244 111944 277296
rect 148784 277244 148836 277296
rect 111800 275952 111852 276004
rect 153016 275952 153068 276004
rect 231676 275952 231728 276004
rect 256700 275952 256752 276004
rect 111892 275884 111944 275936
rect 132224 275884 132276 275936
rect 111892 274592 111944 274644
rect 140504 274592 140556 274644
rect 228916 274592 228968 274644
rect 256700 274592 256752 274644
rect 111800 274524 111852 274576
rect 129372 274524 129424 274576
rect 111892 273164 111944 273216
rect 154028 273164 154080 273216
rect 111800 273028 111852 273080
rect 114468 273028 114520 273080
rect 551284 271872 551336 271924
rect 580172 271872 580224 271924
rect 111892 271804 111944 271856
rect 147404 271804 147456 271856
rect 111800 271736 111852 271788
rect 145840 271736 145892 271788
rect 111800 270444 111852 270496
rect 155776 270444 155828 270496
rect 241244 270444 241296 270496
rect 256700 270444 256752 270496
rect 111892 270376 111944 270428
rect 150072 270376 150124 270428
rect 111892 269016 111944 269068
rect 132132 269016 132184 269068
rect 111800 268948 111852 269000
rect 115756 268948 115808 269000
rect 111800 267656 111852 267708
rect 129280 267656 129332 267708
rect 111892 267588 111944 267640
rect 122564 267588 122616 267640
rect 232872 266976 232924 267028
rect 257436 266976 257488 267028
rect 3056 266364 3108 266416
rect 30196 266364 30248 266416
rect 160376 266364 160428 266416
rect 161572 266364 161624 266416
rect 111892 266296 111944 266348
rect 137652 266296 137704 266348
rect 224868 266296 224920 266348
rect 256700 266296 256752 266348
rect 111800 266228 111852 266280
rect 115664 266228 115716 266280
rect 111892 264868 111944 264920
rect 152924 264868 152976 264920
rect 231584 264868 231636 264920
rect 256700 264868 256752 264920
rect 111800 264800 111852 264852
rect 144644 264800 144696 264852
rect 111892 263508 111944 263560
rect 151636 263508 151688 263560
rect 111800 263440 111852 263492
rect 140412 263440 140464 263492
rect 161480 262896 161532 262948
rect 162400 262896 162452 262948
rect 168380 262896 168432 262948
rect 169024 262896 169076 262948
rect 169760 262896 169812 262948
rect 170680 262896 170732 262948
rect 173900 262896 173952 262948
rect 174820 262896 174872 262948
rect 176660 262896 176712 262948
rect 177304 262896 177356 262948
rect 178040 262896 178092 262948
rect 178960 262896 179012 262948
rect 186320 262896 186372 262948
rect 187240 262896 187292 262948
rect 190460 262896 190512 262948
rect 191380 262896 191432 262948
rect 111800 262148 111852 262200
rect 149980 262148 150032 262200
rect 228824 262148 228876 262200
rect 256700 262148 256752 262200
rect 194600 261264 194652 261316
rect 195520 261264 195572 261316
rect 202880 261264 202932 261316
rect 203800 261264 203852 261316
rect 112904 261060 112956 261112
rect 113088 260992 113140 261044
rect 112996 260924 113048 260976
rect 112904 260856 112956 260908
rect 111800 260788 111852 260840
rect 132040 260788 132092 260840
rect 226064 260788 226116 260840
rect 256700 260788 256752 260840
rect 111892 260720 111944 260772
rect 117044 260720 117096 260772
rect 112260 260652 112312 260704
rect 113180 260652 113232 260704
rect 215300 260380 215352 260432
rect 216220 260380 216272 260432
rect 111892 259360 111944 259412
rect 118056 259360 118108 259412
rect 111800 259292 111852 259344
rect 118148 259292 118200 259344
rect 551376 258068 551428 258120
rect 580172 258068 580224 258120
rect 111892 258000 111944 258052
rect 143264 258000 143316 258052
rect 238300 258000 238352 258052
rect 256700 258000 256752 258052
rect 111800 257932 111852 257984
rect 121092 257932 121144 257984
rect 111800 256640 111852 256692
rect 137560 256640 137612 256692
rect 234344 256640 234396 256692
rect 256700 256640 256752 256692
rect 111800 255212 111852 255264
rect 151360 255212 151412 255264
rect 3516 253920 3568 253972
rect 26884 253920 26936 253972
rect 111800 253852 111852 253904
rect 131948 253852 132000 253904
rect 236920 253852 236972 253904
rect 256700 253852 256752 253904
rect 111892 253784 111944 253836
rect 123944 253784 123996 253836
rect 111800 253716 111852 253768
rect 121000 253716 121052 253768
rect 112352 252968 112404 253020
rect 112720 252968 112772 253020
rect 111800 252492 111852 252544
rect 122472 252492 122524 252544
rect 224776 252492 224828 252544
rect 256700 252492 256752 252544
rect 111800 251132 111852 251184
rect 149888 251132 149940 251184
rect 111892 251064 111944 251116
rect 137468 251064 137520 251116
rect 111800 249704 111852 249756
rect 153936 249704 153988 249756
rect 228732 249704 228784 249756
rect 256700 249704 256752 249756
rect 111892 248344 111944 248396
rect 130844 248344 130896 248396
rect 225972 248344 226024 248396
rect 256700 248344 256752 248396
rect 111800 248276 111852 248328
rect 114376 248276 114428 248328
rect 111892 246984 111944 247036
rect 126704 246984 126756 247036
rect 111800 246916 111852 246968
rect 115572 246916 115624 246968
rect 112904 246304 112956 246356
rect 152832 246304 152884 246356
rect 111800 245556 111852 245608
rect 147312 245556 147364 245608
rect 224684 245556 224736 245608
rect 256700 245556 256752 245608
rect 111892 245488 111944 245540
rect 116952 245488 117004 245540
rect 111800 244196 111852 244248
rect 122380 244196 122432 244248
rect 235540 244196 235592 244248
rect 256700 244196 256752 244248
rect 111984 243516 112036 243568
rect 144460 243516 144512 243568
rect 111800 242836 111852 242888
rect 133420 242836 133472 242888
rect 111892 242156 111944 242208
rect 143172 242156 143224 242208
rect 111800 241408 111852 241460
rect 133328 241408 133380 241460
rect 224592 241408 224644 241460
rect 256700 241408 256752 241460
rect 112352 240728 112404 240780
rect 119712 240728 119764 240780
rect 111800 240048 111852 240100
rect 148692 240048 148744 240100
rect 231492 240048 231544 240100
rect 256700 240048 256752 240100
rect 111892 239980 111944 240032
rect 130752 239980 130804 240032
rect 111800 238688 111852 238740
rect 127992 238688 128044 238740
rect 111892 238484 111944 238536
rect 114284 238484 114336 238536
rect 227444 238008 227496 238060
rect 257804 238008 257856 238060
rect 111800 237328 111852 237380
rect 136088 237328 136140 237380
rect 228640 237328 228692 237380
rect 256700 237328 256752 237380
rect 111892 236648 111944 236700
rect 139032 236648 139084 236700
rect 111800 235900 111852 235952
rect 122288 235900 122340 235952
rect 111892 235220 111944 235272
rect 145656 235220 145708 235272
rect 111800 234540 111852 234592
rect 148600 234540 148652 234592
rect 112352 233928 112404 233980
rect 112628 233928 112680 233980
rect 111800 233860 111852 233912
rect 147220 233860 147272 233912
rect 232780 233860 232832 233912
rect 257344 233860 257396 233912
rect 236828 233180 236880 233232
rect 256700 233180 256752 233232
rect 111800 232908 111852 232960
rect 115480 232908 115532 232960
rect 112812 232500 112864 232552
rect 145748 232500 145800 232552
rect 551468 231820 551520 231872
rect 579620 231820 579672 231872
rect 111800 231752 111852 231804
rect 130660 231752 130712 231804
rect 112904 231072 112956 231124
rect 119620 231072 119672 231124
rect 111800 230392 111852 230444
rect 127900 230392 127952 230444
rect 111892 230324 111944 230376
rect 126612 230324 126664 230376
rect 111800 229032 111852 229084
rect 125048 229032 125100 229084
rect 111892 228964 111944 229016
rect 123852 228964 123904 229016
rect 250720 228964 250772 229016
rect 256700 228964 256752 229016
rect 111800 227672 111852 227724
rect 122196 227672 122248 227724
rect 222752 227672 222804 227724
rect 256700 227672 256752 227724
rect 111892 227604 111944 227656
rect 116860 227604 116912 227656
rect 111800 225972 111852 226024
rect 115388 225972 115440 226024
rect 111800 224884 111852 224936
rect 144552 224884 144604 224936
rect 249524 224884 249576 224936
rect 256700 224884 256752 224936
rect 111892 224816 111944 224868
rect 134616 224816 134668 224868
rect 112812 224408 112864 224460
rect 112996 224408 113048 224460
rect 111800 223524 111852 223576
rect 147128 223524 147180 223576
rect 242348 223524 242400 223576
rect 256700 223524 256752 223576
rect 111892 223456 111944 223508
rect 130568 223456 130620 223508
rect 111800 222096 111852 222148
rect 127808 222096 127860 222148
rect 111892 222028 111944 222080
rect 126520 222028 126572 222080
rect 111800 220736 111852 220788
rect 133144 220736 133196 220788
rect 223488 220736 223540 220788
rect 256700 220736 256752 220788
rect 111892 220668 111944 220720
rect 123760 220668 123812 220720
rect 112628 220056 112680 220108
rect 152740 220056 152792 220108
rect 223396 219376 223448 219428
rect 256700 219376 256752 219428
rect 111892 218696 111944 218748
rect 151268 218696 151320 218748
rect 551560 218016 551612 218068
rect 580172 218016 580224 218068
rect 111800 217948 111852 218000
rect 114192 217948 114244 218000
rect 223304 217948 223356 218000
rect 256700 217948 256752 218000
rect 112628 217268 112680 217320
rect 149796 217268 149848 217320
rect 111800 216588 111852 216640
rect 138940 216588 138992 216640
rect 112720 215908 112772 215960
rect 129188 215908 129240 215960
rect 111800 215228 111852 215280
rect 144368 215228 144420 215280
rect 252008 215228 252060 215280
rect 256700 215228 256752 215280
rect 111892 215160 111944 215212
rect 130476 215160 130528 215212
rect 3332 213936 3384 213988
rect 30288 213936 30340 213988
rect 111800 213868 111852 213920
rect 127716 213868 127768 213920
rect 221832 213868 221884 213920
rect 256700 213868 256752 213920
rect 111892 213800 111944 213852
rect 126428 213800 126480 213852
rect 111800 212440 111852 212492
rect 124956 212440 125008 212492
rect 111892 212372 111944 212424
rect 123576 212372 123628 212424
rect 111800 211080 111852 211132
rect 141700 211080 141752 211132
rect 239680 211080 239732 211132
rect 256700 211080 256752 211132
rect 111892 211012 111944 211064
rect 117964 211012 118016 211064
rect 111800 209720 111852 209772
rect 155684 209720 155736 209772
rect 111800 209040 111852 209092
rect 148508 209040 148560 209092
rect 112628 207748 112680 207800
rect 120908 207748 120960 207800
rect 111984 207680 112036 207732
rect 127624 207680 127676 207732
rect 112076 207612 112128 207664
rect 152648 207612 152700 207664
rect 111800 206932 111852 206984
rect 143080 206932 143132 206984
rect 254860 206932 254912 206984
rect 256700 206932 256752 206984
rect 111892 206864 111944 206916
rect 130384 206864 130436 206916
rect 111800 205572 111852 205624
rect 126336 205572 126388 205624
rect 225880 205572 225932 205624
rect 256700 205572 256752 205624
rect 111892 205504 111944 205556
rect 124864 205504 124916 205556
rect 111800 204212 111852 204264
rect 123668 204212 123720 204264
rect 111892 204008 111944 204060
rect 114100 204008 114152 204060
rect 111800 202784 111852 202836
rect 119528 202784 119580 202836
rect 248052 202784 248104 202836
rect 256700 202784 256752 202836
rect 111892 202716 111944 202768
rect 116768 202716 116820 202768
rect 112260 202104 112312 202156
rect 153844 202104 153896 202156
rect 3240 201492 3292 201544
rect 29552 201492 29604 201544
rect 230204 201424 230256 201476
rect 256700 201424 256752 201476
rect 111800 201356 111852 201408
rect 115296 201356 115348 201408
rect 112996 200744 113048 200796
rect 138848 200744 138900 200796
rect 111892 200064 111944 200116
rect 141608 200064 141660 200116
rect 111800 199996 111852 200048
rect 140320 199996 140372 200048
rect 111800 198636 111852 198688
rect 114008 198636 114060 198688
rect 227352 198636 227404 198688
rect 256700 198636 256752 198688
rect 111800 197276 111852 197328
rect 126244 197276 126296 197328
rect 243912 197276 243964 197328
rect 256700 197276 256752 197328
rect 111800 195916 111852 195968
rect 138756 195916 138808 195968
rect 111892 195848 111944 195900
rect 137376 195848 137428 195900
rect 112536 195236 112588 195288
rect 112996 195236 113048 195288
rect 111800 194488 111852 194540
rect 120816 194488 120868 194540
rect 223212 194488 223264 194540
rect 256700 194488 256752 194540
rect 111892 194420 111944 194472
rect 119436 194420 119488 194472
rect 112904 193808 112956 193860
rect 149704 193808 149756 193860
rect 111892 193128 111944 193180
rect 155592 193128 155644 193180
rect 249432 193128 249484 193180
rect 256700 193128 256752 193180
rect 111800 193060 111852 193112
rect 140228 193060 140280 193112
rect 111800 191700 111852 191752
rect 133236 191700 133288 191752
rect 111800 191156 111852 191208
rect 113916 191156 113968 191208
rect 111892 190408 111944 190460
rect 142988 190408 143040 190460
rect 239588 190408 239640 190460
rect 256700 190408 256752 190460
rect 111800 190340 111852 190392
rect 131856 190340 131908 190392
rect 111892 188980 111944 189032
rect 148416 188980 148468 189032
rect 230112 188980 230164 189032
rect 256700 188980 256752 189032
rect 111800 188912 111852 188964
rect 141516 188912 141568 188964
rect 111892 187620 111944 187672
rect 144276 187620 144328 187672
rect 111800 187552 111852 187604
rect 123484 187552 123536 187604
rect 111800 186260 111852 186312
rect 147036 186260 147088 186312
rect 227260 186260 227312 186312
rect 256700 186260 256752 186312
rect 111892 184832 111944 184884
rect 116676 184832 116728 184884
rect 224500 184832 224552 184884
rect 256700 184832 256752 184884
rect 111800 184764 111852 184816
rect 115204 184764 115256 184816
rect 112812 184152 112864 184204
rect 140136 184152 140188 184204
rect 111800 183472 111852 183524
rect 137284 183472 137336 183524
rect 111800 182112 111852 182164
rect 155500 182112 155552 182164
rect 235448 182112 235500 182164
rect 256700 182112 256752 182164
rect 111800 181772 111852 181824
rect 113824 181772 113876 181824
rect 111892 180752 111944 180804
rect 129004 180752 129056 180804
rect 225788 180752 225840 180804
rect 256700 180752 256752 180804
rect 111800 180684 111852 180736
rect 129096 180684 129148 180736
rect 111892 179324 111944 179376
rect 155408 179324 155460 179376
rect 111800 179256 111852 179308
rect 145564 179256 145616 179308
rect 552664 178032 552716 178084
rect 580172 178032 580224 178084
rect 245108 177964 245160 178016
rect 256700 177964 256752 178016
rect 111984 177284 112036 177336
rect 131764 177284 131816 177336
rect 111800 176604 111852 176656
rect 151176 176604 151228 176656
rect 230020 176604 230072 176656
rect 256700 176604 256752 176656
rect 111892 176536 111944 176588
rect 122104 176536 122156 176588
rect 111800 173816 111852 173868
rect 120724 173816 120776 173868
rect 111892 173748 111944 173800
rect 119344 173748 119396 173800
rect 111800 172456 111852 172508
rect 155224 172456 155276 172508
rect 246764 172456 246816 172508
rect 256700 172456 256752 172508
rect 111892 171028 111944 171080
rect 155316 171028 155368 171080
rect 234252 171028 234304 171080
rect 256700 171028 256752 171080
rect 111800 170960 111852 171012
rect 116584 170960 116636 171012
rect 224408 168308 224460 168360
rect 256700 168308 256752 168360
rect 242256 166948 242308 167000
rect 256700 166948 256752 167000
rect 225696 164160 225748 164212
rect 256700 164160 256752 164212
rect 238208 162800 238260 162852
rect 256700 162800 256752 162852
rect 3424 160760 3476 160812
rect 134616 160760 134668 160812
rect 3332 160692 3384 160744
rect 156880 160692 156932 160744
rect 232688 160012 232740 160064
rect 256700 160012 256752 160064
rect 3608 159332 3660 159384
rect 158352 159332 158404 159384
rect 3516 157972 3568 158024
rect 155224 157972 155276 158024
rect 241152 157972 241204 158024
rect 257528 157972 257580 158024
rect 247960 155864 248012 155916
rect 256700 155864 256752 155916
rect 238116 154504 238168 154556
rect 256700 154504 256752 154556
rect 550088 151784 550140 151836
rect 579988 151784 580040 151836
rect 246672 151716 246724 151768
rect 256700 151716 256752 151768
rect 245016 150356 245068 150408
rect 256700 150356 256752 150408
rect 3424 149064 3476 149116
rect 156972 149064 157024 149116
rect 224316 147568 224368 147620
rect 256700 147568 256752 147620
rect 243820 146208 243872 146260
rect 256700 146208 256752 146260
rect 250628 143488 250680 143540
rect 256700 143488 256752 143540
rect 231400 142060 231452 142112
rect 256700 142060 256752 142112
rect 194600 140700 194652 140752
rect 195520 140700 195572 140752
rect 186320 140632 186372 140684
rect 187240 140632 187292 140684
rect 178040 140428 178092 140480
rect 178960 140428 179012 140480
rect 236736 140020 236788 140072
rect 257436 140020 257488 140072
rect 215300 139884 215352 139936
rect 216220 139884 216272 139936
rect 173900 139408 173952 139460
rect 174820 139408 174872 139460
rect 239496 139340 239548 139392
rect 256700 139340 256752 139392
rect 551652 137980 551704 138032
rect 580172 137980 580224 138032
rect 168380 137300 168432 137352
rect 169024 137300 169076 137352
rect 169760 137300 169812 137352
rect 170680 137300 170732 137352
rect 176660 137300 176712 137352
rect 177304 137300 177356 137352
rect 190460 137300 190512 137352
rect 191380 137300 191432 137352
rect 202880 137300 202932 137352
rect 203800 137300 203852 137352
rect 3424 136620 3476 136672
rect 134708 136620 134760 136672
rect 224224 135192 224276 135244
rect 256700 135192 256752 135244
rect 161388 133900 161440 133952
rect 161664 133900 161716 133952
rect 30104 133832 30156 133884
rect 151268 133832 151320 133884
rect 241060 133832 241112 133884
rect 256700 133832 256752 133884
rect 29920 133764 29972 133816
rect 151176 133764 151228 133816
rect 29552 133696 29604 133748
rect 151360 133696 151412 133748
rect 30288 133628 30340 133680
rect 154028 133628 154080 133680
rect 30196 133560 30248 133612
rect 154120 133560 154172 133612
rect 29736 133492 29788 133544
rect 153844 133492 153896 133544
rect 30012 133424 30064 133476
rect 154212 133424 154264 133476
rect 26884 133356 26936 133408
rect 151452 133356 151504 133408
rect 29828 133288 29880 133340
rect 157156 133288 157208 133340
rect 29644 133220 29696 133272
rect 157064 133220 157116 133272
rect 6920 133152 6972 133204
rect 153936 133152 153988 133204
rect 136548 130364 136600 130416
rect 154948 130364 155000 130416
rect 234160 129684 234212 129736
rect 256700 129684 256752 129736
rect 136548 127576 136600 127628
rect 154948 127576 155000 127628
rect 232596 126896 232648 126948
rect 256700 126896 256752 126948
rect 136548 125536 136600 125588
rect 154948 125604 155000 125656
rect 233976 125536 234028 125588
rect 256700 125536 256752 125588
rect 136180 124108 136232 124160
rect 154488 124108 154540 124160
rect 135260 121388 135312 121440
rect 154948 121456 155000 121508
rect 236644 121388 236696 121440
rect 256700 121388 256752 121440
rect 149060 120096 149112 120148
rect 154580 120096 154632 120148
rect 251916 120028 251968 120080
rect 256700 120028 256752 120080
rect 220452 119824 220504 119876
rect 224224 119824 224276 119876
rect 135444 118600 135496 118652
rect 149060 118600 149112 118652
rect 149060 117308 149112 117360
rect 154580 117308 154632 117360
rect 231308 117240 231360 117292
rect 256700 117240 256752 117292
rect 136548 115880 136600 115932
rect 149060 115880 149112 115932
rect 223120 115880 223172 115932
rect 256700 115880 256752 115932
rect 136548 113092 136600 113144
rect 155408 113092 155460 113144
rect 254768 112888 254820 112940
rect 256700 112888 256752 112940
rect 550180 111800 550232 111852
rect 580172 111800 580224 111852
rect 247868 111732 247920 111784
rect 256700 111732 256752 111784
rect 3424 110440 3476 110492
rect 22744 110440 22796 110492
rect 136548 110372 136600 110424
rect 154764 110372 154816 110424
rect 223028 108944 223080 108996
rect 256700 108944 256752 108996
rect 136548 107584 136600 107636
rect 154948 107584 155000 107636
rect 246580 107584 246632 107636
rect 256700 107584 256752 107636
rect 136732 104864 136784 104916
rect 154580 104864 154632 104916
rect 136548 104796 136600 104848
rect 154856 104796 154908 104848
rect 220360 104796 220412 104848
rect 256700 104796 256752 104848
rect 136180 103436 136232 103488
rect 155500 103436 155552 103488
rect 231216 103436 231268 103488
rect 256700 103436 256752 103488
rect 139400 102144 139452 102196
rect 154580 102144 154632 102196
rect 138848 100716 138900 100768
rect 154948 100716 155000 100768
rect 136180 100648 136232 100700
rect 155316 100648 155368 100700
rect 228548 100648 228600 100700
rect 256700 100648 256752 100700
rect 147036 99356 147088 99408
rect 154948 99356 155000 99408
rect 3424 96636 3476 96688
rect 24124 96636 24176 96688
rect 225604 96568 225656 96620
rect 256700 96568 256752 96620
rect 136548 96228 136600 96280
rect 139400 96228 139452 96280
rect 142160 95208 142212 95260
rect 154948 95208 155000 95260
rect 222936 95140 222988 95192
rect 256700 95140 256752 95192
rect 137284 94460 137336 94512
rect 154856 94460 154908 94512
rect 140136 92488 140188 92540
rect 154580 92488 154632 92540
rect 136088 92420 136140 92472
rect 138848 92420 138900 92472
rect 254676 92420 254728 92472
rect 256700 92420 256752 92472
rect 138756 91060 138808 91112
rect 154948 91060 155000 91112
rect 224224 90992 224276 91044
rect 256700 90992 256752 91044
rect 141608 89700 141660 89752
rect 154948 89700 155000 89752
rect 136548 89632 136600 89684
rect 147036 89632 147088 89684
rect 249340 88272 249392 88324
rect 256700 88272 256752 88324
rect 135812 87320 135864 87372
rect 142160 87320 142212 87372
rect 144276 86980 144328 87032
rect 154948 86980 155000 87032
rect 243728 86912 243780 86964
rect 256700 86912 256752 86964
rect 135260 86844 135312 86896
rect 137284 86844 137336 86896
rect 137376 85552 137428 85604
rect 154948 85552 155000 85604
rect 151636 84192 151688 84244
rect 154948 84192 155000 84244
rect 228456 84124 228508 84176
rect 256700 84124 256752 84176
rect 227168 82764 227220 82816
rect 256700 82764 256752 82816
rect 136548 82220 136600 82272
rect 140136 82220 140188 82272
rect 138848 81404 138900 81456
rect 154948 81404 155000 81456
rect 140228 80044 140280 80096
rect 154764 80044 154816 80096
rect 249156 79976 249208 80028
rect 256700 79976 256752 80028
rect 136088 79704 136140 79756
rect 138756 79704 138808 79756
rect 250536 78616 250588 78668
rect 256700 78616 256752 78668
rect 147036 77256 147088 77308
rect 154948 77256 155000 77308
rect 220268 77188 220320 77240
rect 224868 77188 224920 77240
rect 235356 77188 235408 77240
rect 256700 77188 256752 77240
rect 136548 77052 136600 77104
rect 141608 77052 141660 77104
rect 141516 75896 141568 75948
rect 154948 75896 155000 75948
rect 137284 74536 137336 74588
rect 154948 74536 155000 74588
rect 244924 74468 244976 74520
rect 256700 74468 256752 74520
rect 136548 73720 136600 73772
rect 144276 73720 144328 73772
rect 224868 73108 224920 73160
rect 256700 73108 256752 73160
rect 135720 72428 135772 72480
rect 151636 72428 151688 72480
rect 151544 71748 151596 71800
rect 154580 71748 154632 71800
rect 135352 71612 135404 71664
rect 137376 71612 137428 71664
rect 247776 70320 247828 70372
rect 256700 70320 256752 70372
rect 143080 69028 143132 69080
rect 154580 69028 154632 69080
rect 229836 68960 229888 69012
rect 256700 68960 256752 69012
rect 137376 68280 137428 68332
rect 154948 68280 155000 68332
rect 138756 66240 138808 66292
rect 154948 66240 155000 66292
rect 136088 66172 136140 66224
rect 138848 66172 138900 66224
rect 140136 64880 140188 64932
rect 154580 64880 154632 64932
rect 250444 64404 250496 64456
rect 256700 64404 256752 64456
rect 136548 64132 136600 64184
rect 140228 64132 140280 64184
rect 138848 62092 138900 62144
rect 154580 62092 154632 62144
rect 135628 62024 135680 62076
rect 147036 62024 147088 62076
rect 235264 62024 235316 62076
rect 256700 62024 256752 62076
rect 144276 60732 144328 60784
rect 154948 60732 155000 60784
rect 227076 60664 227128 60716
rect 256700 60664 256752 60716
rect 147036 59372 147088 59424
rect 154948 59372 155000 59424
rect 551744 59372 551796 59424
rect 580080 59372 580132 59424
rect 136548 58964 136600 59016
rect 141516 58964 141568 59016
rect 222844 57876 222896 57928
rect 256700 57876 256752 57928
rect 141516 56584 141568 56636
rect 154948 56584 155000 56636
rect 221740 56516 221792 56568
rect 256700 56516 256752 56568
rect 135260 56380 135312 56432
rect 137284 56380 137336 56432
rect 142988 55224 143040 55276
rect 154948 55224 155000 55276
rect 242164 54476 242216 54528
rect 256700 54476 256752 54528
rect 136548 53728 136600 53780
rect 151544 53728 151596 53780
rect 142804 52776 142856 52828
rect 158444 52640 158496 52692
rect 175602 52640 175654 52692
rect 175878 52640 175930 52692
rect 157064 52572 157116 52624
rect 157156 52504 157208 52556
rect 177258 52640 177310 52692
rect 148416 52436 148468 52488
rect 154948 52436 155000 52488
rect 159916 52368 159968 52420
rect 176982 52368 177034 52420
rect 136640 51960 136692 52012
rect 156604 52028 156656 52080
rect 159824 52028 159876 52080
rect 154212 51892 154264 51944
rect 159916 51960 159968 52012
rect 161434 51892 161486 51944
rect 161802 51892 161854 51944
rect 161894 51892 161946 51944
rect 162998 51892 163050 51944
rect 161066 51824 161118 51876
rect 154120 51756 154172 51808
rect 153200 51688 153252 51740
rect 160698 51756 160750 51808
rect 161618 51824 161670 51876
rect 159364 51620 159416 51672
rect 151452 51552 151504 51604
rect 151084 51484 151136 51536
rect 159272 51484 159324 51536
rect 135996 51416 136048 51468
rect 135904 51348 135956 51400
rect 159456 51348 159508 51400
rect 134708 51280 134760 51332
rect 160192 51280 160244 51332
rect 160928 51620 160980 51672
rect 161112 51620 161164 51672
rect 161296 51484 161348 51536
rect 161756 51688 161808 51740
rect 162998 51756 163050 51808
rect 161848 51620 161900 51672
rect 161940 51552 161992 51604
rect 163734 51892 163786 51944
rect 164010 51892 164062 51944
rect 164194 51892 164246 51944
rect 164378 51892 164430 51944
rect 164562 51892 164614 51944
rect 163366 51824 163418 51876
rect 163550 51756 163602 51808
rect 163412 51688 163464 51740
rect 164286 51824 164338 51876
rect 164148 51620 164200 51672
rect 164516 51756 164568 51808
rect 164424 51688 164476 51740
rect 164930 51892 164982 51944
rect 165022 51892 165074 51944
rect 165114 51892 165166 51944
rect 164838 51824 164890 51876
rect 164608 51620 164660 51672
rect 164240 51552 164292 51604
rect 161756 51484 161808 51536
rect 163596 51484 163648 51536
rect 163964 51484 164016 51536
rect 164976 51756 165028 51808
rect 165068 51688 165120 51740
rect 165482 51892 165534 51944
rect 165666 51892 165718 51944
rect 165758 51892 165810 51944
rect 165942 51892 165994 51944
rect 166034 51892 166086 51944
rect 166218 51892 166270 51944
rect 166310 51892 166362 51944
rect 167138 51892 167190 51944
rect 167322 51892 167374 51944
rect 167414 51892 167466 51944
rect 167874 51892 167926 51944
rect 168058 51892 168110 51944
rect 168150 51892 168202 51944
rect 169162 51892 169214 51944
rect 169346 51892 169398 51944
rect 169622 51892 169674 51944
rect 165528 51756 165580 51808
rect 166402 51824 166454 51876
rect 166586 51824 166638 51876
rect 167046 51824 167098 51876
rect 165896 51688 165948 51740
rect 165988 51688 166040 51740
rect 166172 51688 166224 51740
rect 166264 51688 166316 51740
rect 166494 51756 166546 51808
rect 165712 51620 165764 51672
rect 166356 51620 166408 51672
rect 165068 51484 165120 51536
rect 166080 51552 166132 51604
rect 165620 51416 165672 51468
rect 166448 51416 166500 51468
rect 167230 51824 167282 51876
rect 167000 51688 167052 51740
rect 167184 51688 167236 51740
rect 167506 51824 167558 51876
rect 167414 51756 167466 51808
rect 167092 51620 167144 51672
rect 167368 51620 167420 51672
rect 167460 51620 167512 51672
rect 168012 51688 168064 51740
rect 168242 51824 168294 51876
rect 168886 51824 168938 51876
rect 168104 51620 168156 51672
rect 168702 51756 168754 51808
rect 168840 51688 168892 51740
rect 168748 51620 168800 51672
rect 167828 51552 167880 51604
rect 168196 51552 168248 51604
rect 168380 51552 168432 51604
rect 169898 51824 169950 51876
rect 169300 51620 169352 51672
rect 169576 51620 169628 51672
rect 170128 51620 170180 51672
rect 170726 51892 170778 51944
rect 172014 51892 172066 51944
rect 174682 51892 174734 51944
rect 170358 51824 170410 51876
rect 170910 51824 170962 51876
rect 171002 51824 171054 51876
rect 172290 51824 172342 51876
rect 170588 51688 170640 51740
rect 170496 51552 170548 51604
rect 166908 51484 166960 51536
rect 170128 51484 170180 51536
rect 170312 51484 170364 51536
rect 170864 51620 170916 51672
rect 171968 51620 172020 51672
rect 172152 51620 172204 51672
rect 172934 51756 172986 51808
rect 173026 51756 173078 51808
rect 173302 51824 173354 51876
rect 173394 51756 173446 51808
rect 173578 51756 173630 51808
rect 172980 51620 173032 51672
rect 173072 51620 173124 51672
rect 173164 51620 173216 51672
rect 173348 51620 173400 51672
rect 173624 51620 173676 51672
rect 175694 51892 175746 51944
rect 176522 51892 176574 51944
rect 176062 51824 176114 51876
rect 175740 51688 175792 51740
rect 170680 51484 170732 51536
rect 169760 51348 169812 51400
rect 135352 50940 135404 50992
rect 137376 50940 137428 50992
rect 159824 51212 159876 51264
rect 166908 51212 166960 51264
rect 175648 51552 175700 51604
rect 175740 51552 175792 51604
rect 170956 51484 171008 51536
rect 171876 51416 171928 51468
rect 175648 51416 175700 51468
rect 176016 51552 176068 51604
rect 176614 51756 176666 51808
rect 176568 51620 176620 51672
rect 176798 51892 176850 51944
rect 176384 51552 176436 51604
rect 178362 51892 178414 51944
rect 216680 52776 216732 52828
rect 216036 52708 216088 52760
rect 255872 52504 255924 52556
rect 253388 52436 253440 52488
rect 200258 52368 200310 52420
rect 182778 52028 182830 52080
rect 184342 52028 184394 52080
rect 188114 52028 188166 52080
rect 179006 51892 179058 51944
rect 179098 51892 179150 51944
rect 179374 51892 179426 51944
rect 178822 51824 178874 51876
rect 177074 51756 177126 51808
rect 177120 51552 177172 51604
rect 176108 51484 176160 51536
rect 178500 51552 178552 51604
rect 179282 51824 179334 51876
rect 179466 51824 179518 51876
rect 179558 51824 179610 51876
rect 179052 51688 179104 51740
rect 178960 51416 179012 51468
rect 173440 51348 173492 51400
rect 175740 51348 175792 51400
rect 179604 51688 179656 51740
rect 179420 51620 179472 51672
rect 179512 51552 179564 51604
rect 180110 51892 180162 51944
rect 180202 51892 180254 51944
rect 180478 51892 180530 51944
rect 181122 51892 181174 51944
rect 181214 51892 181266 51944
rect 180018 51824 180070 51876
rect 180570 51824 180622 51876
rect 180432 51756 180484 51808
rect 180662 51756 180714 51808
rect 180846 51756 180898 51808
rect 180524 51688 180576 51740
rect 180616 51620 180668 51672
rect 180340 51484 180392 51536
rect 181582 51824 181634 51876
rect 181260 51756 181312 51808
rect 181168 51620 181220 51672
rect 181858 51756 181910 51808
rect 181628 51688 181680 51740
rect 181168 51484 181220 51536
rect 181444 51484 181496 51536
rect 181720 51484 181772 51536
rect 180800 51416 180852 51468
rect 173716 51280 173768 51332
rect 180064 51348 180116 51400
rect 181076 51348 181128 51400
rect 182226 51892 182278 51944
rect 182318 51892 182370 51944
rect 182502 51892 182554 51944
rect 182594 51892 182646 51944
rect 182686 51892 182738 51944
rect 182870 51892 182922 51944
rect 182134 51824 182186 51876
rect 182364 51756 182416 51808
rect 182548 51688 182600 51740
rect 182272 51620 182324 51672
rect 182732 51620 182784 51672
rect 182640 51552 182692 51604
rect 182916 51552 182968 51604
rect 183146 51892 183198 51944
rect 183238 51892 183290 51944
rect 183330 51892 183382 51944
rect 183698 51892 183750 51944
rect 183882 51892 183934 51944
rect 183974 51892 184026 51944
rect 184066 51892 184118 51944
rect 184250 51892 184302 51944
rect 183284 51756 183336 51808
rect 183192 51688 183244 51740
rect 182088 51484 182140 51536
rect 183008 51484 183060 51536
rect 182732 51348 182784 51400
rect 183652 51756 183704 51808
rect 184388 51824 184440 51876
rect 184204 51756 184256 51808
rect 184020 51688 184072 51740
rect 184112 51688 184164 51740
rect 184388 51688 184440 51740
rect 183928 51620 183980 51672
rect 184296 51620 184348 51672
rect 184894 51892 184946 51944
rect 185170 51892 185222 51944
rect 185262 51892 185314 51944
rect 185354 51892 185406 51944
rect 185446 51892 185498 51944
rect 185078 51756 185130 51808
rect 185216 51688 185268 51740
rect 185308 51688 185360 51740
rect 185400 51688 185452 51740
rect 185032 51620 185084 51672
rect 185124 51620 185176 51672
rect 185584 51620 185636 51672
rect 184848 51484 184900 51536
rect 185584 51484 185636 51536
rect 185906 51892 185958 51944
rect 185814 51824 185866 51876
rect 185768 51416 185820 51468
rect 186274 51892 186326 51944
rect 186550 51892 186602 51944
rect 186090 51824 186142 51876
rect 186366 51824 186418 51876
rect 186826 51824 186878 51876
rect 187470 51892 187522 51944
rect 187838 51892 187890 51944
rect 189494 52164 189546 52216
rect 190414 52028 190466 52080
rect 192254 52028 192306 52080
rect 186228 51620 186280 51672
rect 186504 51620 186556 51672
rect 187286 51824 187338 51876
rect 187378 51824 187430 51876
rect 186964 51620 187016 51672
rect 187148 51620 187200 51672
rect 186320 51552 186372 51604
rect 187424 51620 187476 51672
rect 187516 51620 187568 51672
rect 186044 51484 186096 51536
rect 186596 51484 186648 51536
rect 186780 51484 186832 51536
rect 187700 51484 187752 51536
rect 188206 51824 188258 51876
rect 188298 51824 188350 51876
rect 188482 51824 188534 51876
rect 187976 51484 188028 51536
rect 188344 51620 188396 51672
rect 178960 51280 179012 51332
rect 180892 51280 180944 51332
rect 185860 51348 185912 51400
rect 187976 51348 188028 51400
rect 188666 51756 188718 51808
rect 175096 51212 175148 51264
rect 188436 51280 188488 51332
rect 189218 51892 189270 51944
rect 188942 51824 188994 51876
rect 189172 51484 189224 51536
rect 189264 51484 189316 51536
rect 190138 51892 190190 51944
rect 190230 51892 190282 51944
rect 189586 51824 189638 51876
rect 189770 51824 189822 51876
rect 190184 51756 190236 51808
rect 189448 51620 189500 51672
rect 189724 51620 189776 51672
rect 191334 51892 191386 51944
rect 190782 51824 190834 51876
rect 190874 51824 190926 51876
rect 191242 51824 191294 51876
rect 190368 51484 190420 51536
rect 190552 51484 190604 51536
rect 188896 51416 188948 51468
rect 191104 51484 191156 51536
rect 190828 51416 190880 51468
rect 191610 51892 191662 51944
rect 192070 51892 192122 51944
rect 191702 51824 191754 51876
rect 191794 51756 191846 51808
rect 191886 51756 191938 51808
rect 191978 51756 192030 51808
rect 191748 51552 191800 51604
rect 191840 51552 191892 51604
rect 192116 51688 192168 51740
rect 192024 51552 192076 51604
rect 191656 51484 191708 51536
rect 191380 51416 191432 51468
rect 191932 51416 191984 51468
rect 192622 51892 192674 51944
rect 193174 51824 193226 51876
rect 192576 51756 192628 51808
rect 192944 51484 192996 51536
rect 193450 51824 193502 51876
rect 216036 52368 216088 52420
rect 216220 52300 216272 52352
rect 214426 52164 214478 52216
rect 216312 52164 216364 52216
rect 194002 51892 194054 51944
rect 194094 51892 194146 51944
rect 194186 51892 194238 51944
rect 194278 51892 194330 51944
rect 191564 51348 191616 51400
rect 194370 51824 194422 51876
rect 194462 51824 194514 51876
rect 194048 51688 194100 51740
rect 194140 51688 194192 51740
rect 194324 51552 194376 51604
rect 194416 51552 194468 51604
rect 194738 51892 194790 51944
rect 194922 51892 194974 51944
rect 194784 51756 194836 51808
rect 195198 51892 195250 51944
rect 195290 51892 195342 51944
rect 195382 51892 195434 51944
rect 195566 51892 195618 51944
rect 196026 51892 196078 51944
rect 196210 51892 196262 51944
rect 196486 51892 196538 51944
rect 196854 51892 196906 51944
rect 197222 51892 197274 51944
rect 197314 51892 197366 51944
rect 197682 51892 197734 51944
rect 198050 51892 198102 51944
rect 195060 51620 195112 51672
rect 195658 51824 195710 51876
rect 195336 51688 195388 51740
rect 195428 51620 195480 51672
rect 195612 51620 195664 51672
rect 195244 51552 195296 51604
rect 195520 51552 195572 51604
rect 194600 51484 194652 51536
rect 195980 51484 196032 51536
rect 196532 51620 196584 51672
rect 197406 51824 197458 51876
rect 197498 51824 197550 51876
rect 197268 51688 197320 51740
rect 197360 51688 197412 51740
rect 196716 51552 196768 51604
rect 197176 51552 197228 51604
rect 197544 51552 197596 51604
rect 196808 51484 196860 51536
rect 196900 51484 196952 51536
rect 197866 51824 197918 51876
rect 197728 51552 197780 51604
rect 197958 51756 198010 51808
rect 198004 51620 198056 51672
rect 197820 51484 197872 51536
rect 199062 51892 199114 51944
rect 198786 51824 198838 51876
rect 198510 51756 198562 51808
rect 198464 51620 198516 51672
rect 198740 51620 198792 51672
rect 198280 51552 198332 51604
rect 198648 51552 198700 51604
rect 199338 51824 199390 51876
rect 199522 51824 199574 51876
rect 199798 51824 199850 51876
rect 199982 51824 200034 51876
rect 200074 51824 200126 51876
rect 199200 51620 199252 51672
rect 199660 51620 199712 51672
rect 199844 51620 199896 51672
rect 199936 51620 199988 51672
rect 199384 51552 199436 51604
rect 199016 51484 199068 51536
rect 200718 51824 200770 51876
rect 201086 51824 201138 51876
rect 200212 51620 200264 51672
rect 201730 51892 201782 51944
rect 202190 51892 202242 51944
rect 203018 51892 203070 51944
rect 202006 51824 202058 51876
rect 201638 51756 201690 51808
rect 201776 51756 201828 51808
rect 201684 51620 201736 51672
rect 201868 51620 201920 51672
rect 202650 51824 202702 51876
rect 202926 51824 202978 51876
rect 203386 51824 203438 51876
rect 203570 51824 203622 51876
rect 203662 51824 203714 51876
rect 203754 51824 203806 51876
rect 204030 51824 204082 51876
rect 202236 51620 202288 51672
rect 201040 51552 201092 51604
rect 200948 51484 201000 51536
rect 196716 51416 196768 51468
rect 198556 51416 198608 51468
rect 203064 51620 203116 51672
rect 203432 51620 203484 51672
rect 203524 51620 203576 51672
rect 203616 51552 203668 51604
rect 202604 51484 202656 51536
rect 203248 51484 203300 51536
rect 203892 51620 203944 51672
rect 204398 51892 204450 51944
rect 204260 51620 204312 51672
rect 204076 51552 204128 51604
rect 204582 51892 204634 51944
rect 204674 51892 204726 51944
rect 204766 51892 204818 51944
rect 204858 51892 204910 51944
rect 204950 51892 205002 51944
rect 205042 51892 205094 51944
rect 205318 51892 205370 51944
rect 205502 51892 205554 51944
rect 205594 51892 205646 51944
rect 205686 51892 205738 51944
rect 205778 51892 205830 51944
rect 206238 51892 206290 51944
rect 206606 51892 206658 51944
rect 206698 51892 206750 51944
rect 208630 52028 208682 52080
rect 216128 52096 216180 52148
rect 258724 52096 258776 52148
rect 204628 51688 204680 51740
rect 204720 51688 204772 51740
rect 204444 51484 204496 51536
rect 204950 51756 205002 51808
rect 205272 51756 205324 51808
rect 205456 51756 205508 51808
rect 205870 51824 205922 51876
rect 205732 51756 205784 51808
rect 205640 51688 205692 51740
rect 205364 51620 205416 51672
rect 205962 51756 206014 51808
rect 206422 51824 206474 51876
rect 206606 51756 206658 51808
rect 206790 51824 206842 51876
rect 206974 51892 207026 51944
rect 206744 51688 206796 51740
rect 205640 51552 205692 51604
rect 205916 51552 205968 51604
rect 206192 51552 206244 51604
rect 206376 51552 206428 51604
rect 206284 51484 206336 51536
rect 206928 51756 206980 51808
rect 206928 51620 206980 51672
rect 207158 51892 207210 51944
rect 207894 51892 207946 51944
rect 208262 51892 208314 51944
rect 208354 51892 208406 51944
rect 208446 51892 208498 51944
rect 209090 51892 209142 51944
rect 209458 51892 209510 51944
rect 207020 51552 207072 51604
rect 207434 51824 207486 51876
rect 207710 51824 207762 51876
rect 207250 51756 207302 51808
rect 207204 51552 207256 51604
rect 207756 51620 207808 51672
rect 207664 51552 207716 51604
rect 208216 51688 208268 51740
rect 208308 51688 208360 51740
rect 208538 51824 208590 51876
rect 208906 51824 208958 51876
rect 208400 51620 208452 51672
rect 207388 51484 207440 51536
rect 207480 51484 207532 51536
rect 208676 51688 208728 51740
rect 208952 51620 209004 51672
rect 209044 51620 209096 51672
rect 208676 51552 208728 51604
rect 210010 51892 210062 51944
rect 209918 51824 209970 51876
rect 209504 51620 209556 51672
rect 209596 51552 209648 51604
rect 209688 51484 209740 51536
rect 210654 51892 210706 51944
rect 210838 51824 210890 51876
rect 210608 51756 210660 51808
rect 210792 51620 210844 51672
rect 210056 51552 210108 51604
rect 211390 51892 211442 51944
rect 211482 51756 211534 51808
rect 211252 51552 211304 51604
rect 211436 51552 211488 51604
rect 212770 51892 212822 51944
rect 212862 51892 212914 51944
rect 212954 51892 213006 51944
rect 213230 51892 213282 51944
rect 213414 51892 213466 51944
rect 213690 51892 213742 51944
rect 213782 51892 213834 51944
rect 213966 51892 214018 51944
rect 214886 51892 214938 51944
rect 215070 51892 215122 51944
rect 215162 51892 215214 51944
rect 215254 51892 215306 51944
rect 215438 51892 215490 51944
rect 215714 51892 215766 51944
rect 215806 51892 215858 51944
rect 215944 51892 215996 51944
rect 211758 51824 211810 51876
rect 212034 51824 212086 51876
rect 212586 51824 212638 51876
rect 211712 51620 211764 51672
rect 212540 51688 212592 51740
rect 212816 51756 212868 51808
rect 213046 51824 213098 51876
rect 212908 51688 212960 51740
rect 213276 51688 213328 51740
rect 213506 51824 213558 51876
rect 212172 51552 212224 51604
rect 212724 51552 212776 51604
rect 213000 51552 213052 51604
rect 210332 51484 210384 51536
rect 210976 51484 211028 51536
rect 211620 51484 211672 51536
rect 212448 51484 212500 51536
rect 213690 51756 213742 51808
rect 213552 51552 213604 51604
rect 213644 51552 213696 51604
rect 214058 51824 214110 51876
rect 214150 51824 214202 51876
rect 213920 51688 213972 51740
rect 214012 51688 214064 51740
rect 215116 51756 215168 51808
rect 215208 51756 215260 51808
rect 214840 51688 214892 51740
rect 214104 51620 214156 51672
rect 214932 51552 214984 51604
rect 215760 51756 215812 51808
rect 215852 51756 215904 51808
rect 234712 51824 234764 51876
rect 253572 51756 253624 51808
rect 216588 51688 216640 51740
rect 238760 51688 238812 51740
rect 216128 51620 216180 51672
rect 253480 51620 253532 51672
rect 216404 51552 216456 51604
rect 258816 51552 258868 51604
rect 242900 51484 242952 51536
rect 216220 51416 216272 51468
rect 256332 51416 256384 51468
rect 194508 51348 194560 51400
rect 194784 51348 194836 51400
rect 201592 51348 201644 51400
rect 202052 51348 202104 51400
rect 256240 51348 256292 51400
rect 256148 51280 256200 51332
rect 159456 51144 159508 51196
rect 176384 51144 176436 51196
rect 178776 51144 178828 51196
rect 179144 51144 179196 51196
rect 238024 51212 238076 51264
rect 171876 51076 171928 51128
rect 175004 51076 175056 51128
rect 253204 51144 253256 51196
rect 180248 51076 180300 51128
rect 180800 51076 180852 51128
rect 188896 51076 188948 51128
rect 220820 51076 220872 51128
rect 160192 51008 160244 51060
rect 162860 51008 162912 51060
rect 173440 51008 173492 51060
rect 174912 51008 174964 51060
rect 246488 51008 246540 51060
rect 255964 51008 256016 51060
rect 256700 51008 256752 51060
rect 173716 50940 173768 50992
rect 175280 50940 175332 50992
rect 246396 50940 246448 50992
rect 156696 50804 156748 50856
rect 159824 50804 159876 50856
rect 159272 50736 159324 50788
rect 170956 50872 171008 50924
rect 172244 50872 172296 50924
rect 231124 50872 231176 50924
rect 171784 50804 171836 50856
rect 220176 50804 220228 50856
rect 175556 50736 175608 50788
rect 148324 50668 148376 50720
rect 175924 50668 175976 50720
rect 179236 50736 179288 50788
rect 220084 50736 220136 50788
rect 218060 50668 218112 50720
rect 151360 50600 151412 50652
rect 179052 50600 179104 50652
rect 179788 50600 179840 50652
rect 180524 50600 180576 50652
rect 188712 50600 188764 50652
rect 188896 50600 188948 50652
rect 189172 50600 189224 50652
rect 190368 50600 190420 50652
rect 201592 50600 201644 50652
rect 204628 50600 204680 50652
rect 253204 50600 253256 50652
rect 159824 50532 159876 50584
rect 178040 50532 178092 50584
rect 178408 50532 178460 50584
rect 179512 50532 179564 50584
rect 134524 50464 134576 50516
rect 177948 50464 178000 50516
rect 196440 50532 196492 50584
rect 202052 50532 202104 50584
rect 205640 50532 205692 50584
rect 206100 50532 206152 50584
rect 206284 50532 206336 50584
rect 208032 50532 208084 50584
rect 200488 50464 200540 50516
rect 214932 50532 214984 50584
rect 258724 50532 258776 50584
rect 253296 50464 253348 50516
rect 154028 50396 154080 50448
rect 177764 50396 177816 50448
rect 179512 50396 179564 50448
rect 179880 50396 179932 50448
rect 183836 50396 183888 50448
rect 184940 50396 184992 50448
rect 188712 50396 188764 50448
rect 197544 50396 197596 50448
rect 160376 50328 160428 50380
rect 160560 50328 160612 50380
rect 172336 50328 172388 50380
rect 179236 50328 179288 50380
rect 190644 50328 190696 50380
rect 207112 50328 207164 50380
rect 207296 50328 207348 50380
rect 207480 50328 207532 50380
rect 144184 50260 144236 50312
rect 176568 50260 176620 50312
rect 188344 50260 188396 50312
rect 141424 50192 141476 50244
rect 176016 50192 176068 50244
rect 188068 50192 188120 50244
rect 188804 50192 188856 50244
rect 159456 50124 159508 50176
rect 161848 50124 161900 50176
rect 171232 50124 171284 50176
rect 171876 50124 171928 50176
rect 174268 50124 174320 50176
rect 178868 50124 178920 50176
rect 184940 50124 184992 50176
rect 185584 50124 185636 50176
rect 190184 50124 190236 50176
rect 190368 50124 190420 50176
rect 193404 50124 193456 50176
rect 193956 50124 194008 50176
rect 138664 50056 138716 50108
rect 176292 50056 176344 50108
rect 204260 50260 204312 50312
rect 210608 50328 210660 50380
rect 210700 50328 210752 50380
rect 210884 50328 210936 50380
rect 211804 50328 211856 50380
rect 211988 50328 212040 50380
rect 213460 50396 213512 50448
rect 214196 50396 214248 50448
rect 256608 50396 256660 50448
rect 210332 50260 210384 50312
rect 214932 50260 214984 50312
rect 204996 50192 205048 50244
rect 206192 50192 206244 50244
rect 207480 50192 207532 50244
rect 207848 50192 207900 50244
rect 208032 50192 208084 50244
rect 208308 50192 208360 50244
rect 208492 50192 208544 50244
rect 209412 50192 209464 50244
rect 211988 50192 212040 50244
rect 252560 50328 252612 50380
rect 580080 50328 580132 50380
rect 580816 50328 580868 50380
rect 204812 50124 204864 50176
rect 205088 50124 205140 50176
rect 205180 50124 205232 50176
rect 205640 50124 205692 50176
rect 206100 50124 206152 50176
rect 206376 50124 206428 50176
rect 208400 50124 208452 50176
rect 208584 50124 208636 50176
rect 223580 50056 223632 50108
rect 158076 49988 158128 50040
rect 161480 49988 161532 50040
rect 175648 49988 175700 50040
rect 178132 49988 178184 50040
rect 205364 49988 205416 50040
rect 205916 49988 205968 50040
rect 207204 49988 207256 50040
rect 207388 49988 207440 50040
rect 208400 49988 208452 50040
rect 209136 49988 209188 50040
rect 212724 49988 212776 50040
rect 213092 49988 213144 50040
rect 158536 49920 158588 49972
rect 168472 49920 168524 49972
rect 207112 49920 207164 49972
rect 211988 49920 212040 49972
rect 158168 49852 158220 49904
rect 176752 49852 176804 49904
rect 181996 49852 182048 49904
rect 182180 49852 182232 49904
rect 204076 49852 204128 49904
rect 211252 49852 211304 49904
rect 181812 49784 181864 49836
rect 184664 49784 184716 49836
rect 201040 49784 201092 49836
rect 216588 49920 216640 49972
rect 212908 49852 212960 49904
rect 213368 49852 213420 49904
rect 212632 49784 212684 49836
rect 220176 49784 220228 49836
rect 182180 49716 182232 49768
rect 184020 49716 184072 49768
rect 204444 49716 204496 49768
rect 207848 49716 207900 49768
rect 212540 49716 212592 49768
rect 212724 49716 212776 49768
rect 212908 49716 212960 49768
rect 256056 49716 256108 49768
rect 158628 49648 158680 49700
rect 161940 49648 161992 49700
rect 187700 49648 187752 49700
rect 188068 49648 188120 49700
rect 203892 49648 203944 49700
rect 208032 49648 208084 49700
rect 158168 49580 158220 49632
rect 159456 49580 159508 49632
rect 160836 49580 160888 49632
rect 161020 49580 161072 49632
rect 175372 49580 175424 49632
rect 234620 49580 234672 49632
rect 160192 49512 160244 49564
rect 161112 49512 161164 49564
rect 173164 49512 173216 49564
rect 177028 49512 177080 49564
rect 157800 49444 157852 49496
rect 167000 49444 167052 49496
rect 172152 49444 172204 49496
rect 228364 49512 228416 49564
rect 209688 49444 209740 49496
rect 157984 49376 158036 49428
rect 160100 49376 160152 49428
rect 160560 49308 160612 49360
rect 161388 49308 161440 49360
rect 178500 49376 178552 49428
rect 186780 49376 186832 49428
rect 187700 49376 187752 49428
rect 193680 49376 193732 49428
rect 212908 49376 212960 49428
rect 172520 49308 172572 49360
rect 176936 49308 176988 49360
rect 211988 49308 212040 49360
rect 218244 49308 218296 49360
rect 220176 49444 220228 49496
rect 260104 49376 260156 49428
rect 259000 49308 259052 49360
rect 158352 49172 158404 49224
rect 172704 49240 172756 49292
rect 177948 49240 178000 49292
rect 186780 49240 186832 49292
rect 186964 49240 187016 49292
rect 203708 49240 203760 49292
rect 206652 49240 206704 49292
rect 208308 49240 208360 49292
rect 258632 49240 258684 49292
rect 167460 49172 167512 49224
rect 168472 49172 168524 49224
rect 171968 49172 172020 49224
rect 173808 49172 173860 49224
rect 208216 49172 208268 49224
rect 258908 49172 258960 49224
rect 157708 49104 157760 49156
rect 165804 49104 165856 49156
rect 179604 49104 179656 49156
rect 179880 49104 179932 49156
rect 186964 49104 187016 49156
rect 187148 49104 187200 49156
rect 157616 49036 157668 49088
rect 165528 49036 165580 49088
rect 172796 49036 172848 49088
rect 177856 49036 177908 49088
rect 179788 49036 179840 49088
rect 188068 49036 188120 49088
rect 161388 48968 161440 49020
rect 176200 48968 176252 49020
rect 179604 48968 179656 49020
rect 187332 48968 187384 49020
rect 173256 48900 173308 48952
rect 177948 48900 178000 48952
rect 179420 48900 179472 48952
rect 179788 48900 179840 48952
rect 182364 48900 182416 48952
rect 184572 48900 184624 48952
rect 161572 48832 161624 48884
rect 162124 48832 162176 48884
rect 177120 48832 177172 48884
rect 183928 48832 183980 48884
rect 186228 48832 186280 48884
rect 187332 48832 187384 48884
rect 197544 48900 197596 48952
rect 198096 48900 198148 48952
rect 209596 49036 209648 49088
rect 259184 49104 259236 49156
rect 211988 48968 212040 49020
rect 209136 48900 209188 48952
rect 209780 48900 209832 48952
rect 210240 48900 210292 48952
rect 210608 48900 210660 48952
rect 210884 48832 210936 48884
rect 156880 48424 156932 48476
rect 179328 48764 179380 48816
rect 196256 48764 196308 48816
rect 196532 48764 196584 48816
rect 210056 48764 210108 48816
rect 210424 48764 210476 48816
rect 211528 48764 211580 48816
rect 211988 48764 212040 48816
rect 161756 48696 161808 48748
rect 162032 48696 162084 48748
rect 163228 48696 163280 48748
rect 163596 48696 163648 48748
rect 163688 48696 163740 48748
rect 169024 48696 169076 48748
rect 169484 48696 169536 48748
rect 177304 48696 177356 48748
rect 183376 48696 183428 48748
rect 200028 48696 200080 48748
rect 204444 48696 204496 48748
rect 205732 48696 205784 48748
rect 259276 49036 259328 49088
rect 159640 48628 159692 48680
rect 162768 48628 162820 48680
rect 163136 48628 163188 48680
rect 161480 48560 161532 48612
rect 165252 48560 165304 48612
rect 159732 48492 159784 48544
rect 163044 48492 163096 48544
rect 158444 48424 158496 48476
rect 161204 48424 161256 48476
rect 163596 48424 163648 48476
rect 164516 48424 164568 48476
rect 164792 48424 164844 48476
rect 165252 48424 165304 48476
rect 155224 48356 155276 48408
rect 178684 48628 178736 48680
rect 179052 48628 179104 48680
rect 183744 48628 183796 48680
rect 186688 48628 186740 48680
rect 188620 48628 188672 48680
rect 197360 48628 197412 48680
rect 198004 48628 198056 48680
rect 199200 48628 199252 48680
rect 203984 48628 204036 48680
rect 206284 48628 206336 48680
rect 259368 48968 259420 49020
rect 214012 48900 214064 48952
rect 216128 48900 216180 48952
rect 215300 48832 215352 48884
rect 215760 48832 215812 48884
rect 214104 48764 214156 48816
rect 214288 48764 214340 48816
rect 214380 48764 214432 48816
rect 214932 48764 214984 48816
rect 215576 48764 215628 48816
rect 216036 48764 216088 48816
rect 214012 48696 214064 48748
rect 214748 48696 214800 48748
rect 215668 48628 215720 48680
rect 215944 48628 215996 48680
rect 172060 48492 172112 48544
rect 254584 48560 254636 48612
rect 177672 48492 177724 48544
rect 179788 48492 179840 48544
rect 184204 48492 184256 48544
rect 185032 48492 185084 48544
rect 173624 48424 173676 48476
rect 208308 48492 208360 48544
rect 210148 48492 210200 48544
rect 210976 48492 211028 48544
rect 212540 48492 212592 48544
rect 213184 48492 213236 48544
rect 214196 48492 214248 48544
rect 214472 48492 214524 48544
rect 196072 48424 196124 48476
rect 199844 48424 199896 48476
rect 200120 48424 200172 48476
rect 203892 48424 203944 48476
rect 208124 48424 208176 48476
rect 215944 48424 215996 48476
rect 179144 48356 179196 48408
rect 179972 48356 180024 48408
rect 180524 48356 180576 48408
rect 184020 48356 184072 48408
rect 198280 48356 198332 48408
rect 202512 48356 202564 48408
rect 203156 48356 203208 48408
rect 204628 48356 204680 48408
rect 210884 48356 210936 48408
rect 216680 48356 216732 48408
rect 164424 48288 164476 48340
rect 164976 48288 165028 48340
rect 179236 48288 179288 48340
rect 179512 48288 179564 48340
rect 196532 48288 196584 48340
rect 196992 48288 197044 48340
rect 202052 48288 202104 48340
rect 203708 48288 203760 48340
rect 213184 48288 213236 48340
rect 213552 48288 213604 48340
rect 214380 48288 214432 48340
rect 216312 48288 216364 48340
rect 156972 48084 157024 48136
rect 178408 48220 178460 48272
rect 162124 48152 162176 48204
rect 162492 48152 162544 48204
rect 162860 48152 162912 48204
rect 164240 48152 164292 48204
rect 164792 48152 164844 48204
rect 165620 48152 165672 48204
rect 175188 48152 175240 48204
rect 251824 48220 251876 48272
rect 161664 48084 161716 48136
rect 162400 48084 162452 48136
rect 165068 48084 165120 48136
rect 165344 48084 165396 48136
rect 174728 48084 174780 48136
rect 243636 48152 243688 48204
rect 201500 48084 201552 48136
rect 253664 48084 253716 48136
rect 156788 48016 156840 48068
rect 178224 48016 178276 48068
rect 180800 48016 180852 48068
rect 183836 48016 183888 48068
rect 190644 48016 190696 48068
rect 190828 48016 190880 48068
rect 190920 48016 190972 48068
rect 191380 48016 191432 48068
rect 196164 48016 196216 48068
rect 196440 48016 196492 48068
rect 205640 48016 205692 48068
rect 259092 48016 259144 48068
rect 146944 47948 146996 48000
rect 176844 47948 176896 48000
rect 179604 47948 179656 48000
rect 180616 47948 180668 48000
rect 189908 47948 189960 48000
rect 244280 47948 244332 48000
rect 164700 47880 164752 47932
rect 165436 47880 165488 47932
rect 169116 47880 169168 47932
rect 169760 47880 169812 47932
rect 179696 47880 179748 47932
rect 180064 47880 180116 47932
rect 190368 47880 190420 47932
rect 248420 47880 248472 47932
rect 190460 47812 190512 47864
rect 251180 47812 251232 47864
rect 159364 47744 159416 47796
rect 169668 47744 169720 47796
rect 195704 47744 195756 47796
rect 256424 47744 256476 47796
rect 134524 47676 134576 47728
rect 160836 47676 160888 47728
rect 191932 47676 191984 47728
rect 255964 47676 256016 47728
rect 134616 47608 134668 47660
rect 168288 47608 168340 47660
rect 192024 47608 192076 47660
rect 256516 47608 256568 47660
rect 133144 47540 133196 47592
rect 166724 47540 166776 47592
rect 167276 47540 167328 47592
rect 167644 47540 167696 47592
rect 173256 47540 173308 47592
rect 182640 47540 182692 47592
rect 191564 47540 191616 47592
rect 255320 47540 255372 47592
rect 152464 47472 152516 47524
rect 177764 47472 177816 47524
rect 193220 47472 193272 47524
rect 193864 47472 193916 47524
rect 203064 47472 203116 47524
rect 253756 47472 253808 47524
rect 136548 47404 136600 47456
rect 143080 47404 143132 47456
rect 159548 47404 159600 47456
rect 160284 47404 160336 47456
rect 163228 47404 163280 47456
rect 164148 47404 164200 47456
rect 167460 47404 167512 47456
rect 167736 47404 167788 47456
rect 176660 47404 176712 47456
rect 181812 47404 181864 47456
rect 189356 47404 189408 47456
rect 190368 47404 190420 47456
rect 193680 47404 193732 47456
rect 194600 47404 194652 47456
rect 194784 47404 194836 47456
rect 195520 47404 195572 47456
rect 196164 47404 196216 47456
rect 197084 47404 197136 47456
rect 205824 47404 205876 47456
rect 224224 47404 224276 47456
rect 175464 47336 175516 47388
rect 218152 47336 218204 47388
rect 167000 47268 167052 47320
rect 167828 47268 167880 47320
rect 178868 47268 178920 47320
rect 184388 47268 184440 47320
rect 189448 47268 189500 47320
rect 190184 47268 190236 47320
rect 177764 47200 177816 47252
rect 181536 47200 181588 47252
rect 177488 47132 177540 47184
rect 180892 47132 180944 47184
rect 181260 47132 181312 47184
rect 181444 47132 181496 47184
rect 184388 47132 184440 47184
rect 184848 47132 184900 47184
rect 178684 47064 178736 47116
rect 183284 47064 183336 47116
rect 198832 47064 198884 47116
rect 199200 47064 199252 47116
rect 178776 46996 178828 47048
rect 181904 46996 181956 47048
rect 159456 46928 159508 46980
rect 163412 46928 163464 46980
rect 168564 46928 168616 46980
rect 169208 46928 169260 46980
rect 177580 46928 177632 46980
rect 180340 46928 180392 46980
rect 183560 46928 183612 46980
rect 184940 46928 184992 46980
rect 185860 46928 185912 46980
rect 186044 46928 186096 46980
rect 186964 46928 187016 46980
rect 190092 46928 190144 46980
rect 204628 46928 204680 46980
rect 205180 46928 205232 46980
rect 172980 46860 173032 46912
rect 247684 46860 247736 46912
rect 167368 46792 167420 46844
rect 168104 46792 168156 46844
rect 173532 46792 173584 46844
rect 240876 46792 240928 46844
rect 151268 46724 151320 46776
rect 178592 46724 178644 46776
rect 204352 46724 204404 46776
rect 204628 46724 204680 46776
rect 153844 46656 153896 46708
rect 177212 46656 177264 46708
rect 188436 46656 188488 46708
rect 151176 46588 151228 46640
rect 177396 46588 177448 46640
rect 189540 46588 189592 46640
rect 161848 46520 161900 46572
rect 162216 46520 162268 46572
rect 191012 46520 191064 46572
rect 138664 46452 138716 46504
rect 159916 46452 159968 46504
rect 185216 46452 185268 46504
rect 185860 46452 185912 46504
rect 153200 46384 153252 46436
rect 182916 46384 182968 46436
rect 186780 46384 186832 46436
rect 191012 46384 191064 46436
rect 134708 46316 134760 46368
rect 168380 46316 168432 46368
rect 171324 46316 171376 46368
rect 171508 46316 171560 46368
rect 175280 46316 175332 46368
rect 182364 46316 182416 46368
rect 185216 46316 185268 46368
rect 185768 46316 185820 46368
rect 190460 46316 190512 46368
rect 191196 46316 191248 46368
rect 143540 46248 143592 46300
rect 182088 46248 182140 46300
rect 182916 46248 182968 46300
rect 183468 46248 183520 46300
rect 186596 46248 186648 46300
rect 188528 46248 188580 46300
rect 190736 46248 190788 46300
rect 191288 46248 191340 46300
rect 135996 46180 136048 46232
rect 180248 46180 180300 46232
rect 185308 46180 185360 46232
rect 185768 46180 185820 46232
rect 188068 46180 188120 46232
rect 188712 46180 188764 46232
rect 192484 46180 192536 46232
rect 192760 46180 192812 46232
rect 201500 46656 201552 46708
rect 201776 46656 201828 46708
rect 201408 46588 201460 46640
rect 201868 46588 201920 46640
rect 211068 46520 211120 46572
rect 211712 46520 211764 46572
rect 204444 46452 204496 46504
rect 205272 46452 205324 46504
rect 211344 46452 211396 46504
rect 211804 46452 211856 46504
rect 201592 46384 201644 46436
rect 202328 46384 202380 46436
rect 204352 46384 204404 46436
rect 204996 46384 205048 46436
rect 211160 46384 211212 46436
rect 211712 46384 211764 46436
rect 212632 46384 212684 46436
rect 212816 46384 212868 46436
rect 227720 46316 227772 46368
rect 237380 46248 237432 46300
rect 259460 46180 259512 46232
rect 161940 46112 161992 46164
rect 162584 46112 162636 46164
rect 166356 46112 166408 46164
rect 166908 46112 166960 46164
rect 169760 46112 169812 46164
rect 170036 46112 170088 46164
rect 171508 46112 171560 46164
rect 171692 46112 171744 46164
rect 177488 46112 177540 46164
rect 177764 46112 177816 46164
rect 197360 46112 197412 46164
rect 198372 46112 198424 46164
rect 201684 46112 201736 46164
rect 202052 46112 202104 46164
rect 203064 46112 203116 46164
rect 203432 46112 203484 46164
rect 204444 46112 204496 46164
rect 204720 46112 204772 46164
rect 205732 46112 205784 46164
rect 206468 46112 206520 46164
rect 207112 46112 207164 46164
rect 207940 46112 207992 46164
rect 210424 46112 210476 46164
rect 210700 46112 210752 46164
rect 211804 46112 211856 46164
rect 212080 46112 212132 46164
rect 212448 46112 212500 46164
rect 212816 46112 212868 46164
rect 170128 46044 170180 46096
rect 170956 46044 171008 46096
rect 185308 46044 185360 46096
rect 185952 46044 186004 46096
rect 189264 46044 189316 46096
rect 190000 46044 190052 46096
rect 193312 46044 193364 46096
rect 193956 46044 194008 46096
rect 199108 46044 199160 46096
rect 199568 46044 199620 46096
rect 200212 46044 200264 46096
rect 201316 46044 201368 46096
rect 201500 46044 201552 46096
rect 202236 46044 202288 46096
rect 202880 46044 202932 46096
rect 203524 46044 203576 46096
rect 204260 46044 204312 46096
rect 204812 46044 204864 46096
rect 205824 46044 205876 46096
rect 206560 46044 206612 46096
rect 168932 45976 168984 46028
rect 169576 45976 169628 46028
rect 170036 45976 170088 46028
rect 170680 45976 170732 46028
rect 171140 45976 171192 46028
rect 171692 45976 171744 46028
rect 198832 45976 198884 46028
rect 199476 45976 199528 46028
rect 200304 45976 200356 46028
rect 200672 45976 200724 46028
rect 200764 45976 200816 46028
rect 201132 45976 201184 46028
rect 201684 45976 201736 46028
rect 202420 45976 202472 46028
rect 204720 45976 204772 46028
rect 205088 45976 205140 46028
rect 193312 45908 193364 45960
rect 194140 45908 194192 45960
rect 207296 45908 207348 45960
rect 207756 45908 207808 45960
rect 167736 45840 167788 45892
rect 168196 45840 168248 45892
rect 198740 45840 198792 45892
rect 199476 45840 199528 45892
rect 200304 45840 200356 45892
rect 201224 45840 201276 45892
rect 211344 45772 211396 45824
rect 212172 45772 212224 45824
rect 198740 45704 198792 45756
rect 199660 45704 199712 45756
rect 135628 45500 135680 45552
rect 138756 45500 138808 45552
rect 158720 45432 158772 45484
rect 160008 45432 160060 45484
rect 185584 45228 185636 45280
rect 189724 45228 189776 45280
rect 162952 45160 163004 45212
rect 164056 45160 164108 45212
rect 168380 45024 168432 45076
rect 177120 45024 177172 45076
rect 155960 44956 156012 45008
rect 183100 45024 183152 45076
rect 143632 44888 143684 44940
rect 181996 44956 182048 45008
rect 188436 44956 188488 45008
rect 226340 44956 226392 45008
rect 178040 44888 178092 44940
rect 184664 44888 184716 44940
rect 190276 44888 190328 44940
rect 249800 44888 249852 44940
rect 139400 44820 139452 44872
rect 181628 44820 181680 44872
rect 190920 44820 190972 44872
rect 253940 44820 253992 44872
rect 203156 44412 203208 44464
rect 203616 44412 203668 44464
rect 171140 44140 171192 44192
rect 180524 44140 180576 44192
rect 203708 44140 203760 44192
rect 203984 44140 204036 44192
rect 187608 44072 187660 44124
rect 191104 44072 191156 44124
rect 208768 44004 208820 44056
rect 209228 44004 209280 44056
rect 174820 43868 174872 43920
rect 182824 43868 182876 43920
rect 208768 43868 208820 43920
rect 209320 43868 209372 43920
rect 174636 43800 174688 43852
rect 157340 43528 157392 43580
rect 183192 43732 183244 43784
rect 184112 43664 184164 43716
rect 190368 43664 190420 43716
rect 190184 43596 190236 43648
rect 189908 43528 189960 43580
rect 236000 43596 236052 43648
rect 136548 43460 136600 43512
rect 140136 43460 140188 43512
rect 151820 43460 151872 43512
rect 174820 43460 174872 43512
rect 176752 43460 176804 43512
rect 184572 43460 184624 43512
rect 191380 43460 191432 43512
rect 240140 43528 240192 43580
rect 136640 43392 136692 43444
rect 180892 43392 180944 43444
rect 242992 43460 243044 43512
rect 258080 43392 258132 43444
rect 197084 43324 197136 43376
rect 197544 43324 197596 43376
rect 201408 43324 201460 43376
rect 201776 43324 201828 43376
rect 211068 43324 211120 43376
rect 211528 43324 211580 43376
rect 160928 43256 160980 43308
rect 161296 43256 161348 43308
rect 192024 42984 192076 43036
rect 192300 42984 192352 43036
rect 213000 42984 213052 43036
rect 213828 42984 213880 43036
rect 163320 42848 163372 42900
rect 163964 42848 164016 42900
rect 192300 42848 192352 42900
rect 192668 42848 192720 42900
rect 186044 42780 186096 42832
rect 189908 42780 189960 42832
rect 165988 42576 166040 42628
rect 166264 42576 166316 42628
rect 165896 42440 165948 42492
rect 166816 42440 166868 42492
rect 170496 42032 170548 42084
rect 580908 42032 580960 42084
rect 170588 41964 170640 42016
rect 580724 41964 580776 42016
rect 171692 41896 171744 41948
rect 580448 41896 580500 41948
rect 173808 41828 173860 41880
rect 580540 41828 580592 41880
rect 166264 41624 166316 41676
rect 166632 41624 166684 41676
rect 172520 41420 172572 41472
rect 173348 41420 173400 41472
rect 170312 41352 170364 41404
rect 580172 41352 580224 41404
rect 136088 41284 136140 41336
rect 138848 41284 138900 41336
rect 171600 41284 171652 41336
rect 580356 41284 580408 41336
rect 171508 41216 171560 41268
rect 580264 41216 580316 41268
rect 172152 41148 172204 41200
rect 580816 41148 580868 41200
rect 170404 41080 170456 41132
rect 550180 41080 550232 41132
rect 171692 41012 171744 41064
rect 551468 41012 551520 41064
rect 193956 40808 194008 40860
rect 287060 40808 287112 40860
rect 198188 40740 198240 40792
rect 350540 40740 350592 40792
rect 200948 40672 201000 40724
rect 382280 40672 382332 40724
rect 170036 39992 170088 40044
rect 580080 39992 580132 40044
rect 170220 39924 170272 39976
rect 551744 39924 551796 39976
rect 170128 39856 170180 39908
rect 551652 39856 551704 39908
rect 171232 39788 171284 39840
rect 551560 39788 551612 39840
rect 171324 39720 171376 39772
rect 551284 39720 551336 39772
rect 171416 39652 171468 39704
rect 551376 39652 551428 39704
rect 198096 39516 198148 39568
rect 347780 39516 347832 39568
rect 199476 39448 199528 39500
rect 357440 39448 357492 39500
rect 203708 39380 203760 39432
rect 365720 39380 365772 39432
rect 199384 39312 199436 39364
rect 361580 39312 361632 39364
rect 172520 38564 172572 38616
rect 574744 38564 574796 38616
rect 172612 38496 172664 38548
rect 573364 38496 573416 38548
rect 196808 38292 196860 38344
rect 332600 38292 332652 38344
rect 202144 38224 202196 38276
rect 400220 38224 400272 38276
rect 209228 38156 209280 38208
rect 462964 38156 463016 38208
rect 207664 38088 207716 38140
rect 474740 38088 474792 38140
rect 136548 38020 136600 38072
rect 144276 38020 144328 38072
rect 210608 38020 210660 38072
rect 505100 38020 505152 38072
rect 210516 37952 210568 38004
rect 507860 37952 507912 38004
rect 140780 37884 140832 37936
rect 181352 37884 181404 37936
rect 213368 37884 213420 37936
rect 539600 37884 539652 37936
rect 200856 37068 200908 37120
rect 385040 37068 385092 37120
rect 211988 37000 212040 37052
rect 450544 37000 450596 37052
rect 211896 36932 211948 36984
rect 479524 36932 479576 36984
rect 213276 36864 213328 36916
rect 543740 36864 543792 36916
rect 213184 36796 213236 36848
rect 547880 36796 547932 36848
rect 216036 36728 216088 36780
rect 554780 36728 554832 36780
rect 154580 36660 154632 36712
rect 182456 36660 182508 36712
rect 214748 36660 214800 36712
rect 557540 36660 557592 36712
rect 169944 36592 169996 36644
rect 580356 36592 580408 36644
rect 169760 36524 169812 36576
rect 580264 36524 580316 36576
rect 136548 35844 136600 35896
rect 147036 35844 147088 35896
rect 193864 35436 193916 35488
rect 298100 35436 298152 35488
rect 199292 35368 199344 35420
rect 364340 35368 364392 35420
rect 209044 35300 209096 35352
rect 489920 35300 489972 35352
rect 209136 35232 209188 35284
rect 494060 35232 494112 35284
rect 138020 35164 138072 35216
rect 181720 35164 181772 35216
rect 214656 35164 214708 35216
rect 561680 35164 561732 35216
rect 199568 33872 199620 33924
rect 324320 33872 324372 33924
rect 196716 33804 196768 33856
rect 324412 33804 324464 33856
rect 169760 33736 169812 33788
rect 184480 33736 184532 33788
rect 214564 33736 214616 33788
rect 564440 33736 564492 33788
rect 136548 32988 136600 33040
rect 141516 32988 141568 33040
rect 205272 32512 205324 32564
rect 372620 32512 372672 32564
rect 210424 32444 210476 32496
rect 512000 32444 512052 32496
rect 188252 32376 188304 32428
rect 213184 32376 213236 32428
rect 215852 32376 215904 32428
rect 576860 32376 576912 32428
rect 195428 31288 195480 31340
rect 311900 31288 311952 31340
rect 196624 31220 196676 31272
rect 331220 31220 331272 31272
rect 207940 31152 207992 31204
rect 425060 31152 425112 31204
rect 214472 31084 214524 31136
rect 487804 31084 487856 31136
rect 211804 31016 211856 31068
rect 529940 31016 529992 31068
rect 195336 29928 195388 29980
rect 313280 29928 313332 29980
rect 198004 29860 198056 29912
rect 340880 29860 340932 29912
rect 202052 29792 202104 29844
rect 394700 29792 394752 29844
rect 213092 29724 213144 29776
rect 538220 29724 538272 29776
rect 215760 29656 215812 29708
rect 572720 29656 572772 29708
rect 179420 29588 179472 29640
rect 579620 29588 579672 29640
rect 135444 29044 135496 29096
rect 142988 29044 143040 29096
rect 192484 28568 192536 28620
rect 281540 28568 281592 28620
rect 195244 28500 195296 28552
rect 307760 28500 307812 28552
rect 195152 28432 195204 28484
rect 309140 28432 309192 28484
rect 199200 28364 199252 28416
rect 358820 28364 358872 28416
rect 200764 28296 200816 28348
rect 386420 28296 386472 28348
rect 136548 28228 136600 28280
rect 148416 28228 148468 28280
rect 214380 28228 214432 28280
rect 558920 28228 558972 28280
rect 193772 27208 193824 27260
rect 292672 27208 292724 27260
rect 197912 27140 197964 27192
rect 345020 27140 345072 27192
rect 200672 27072 200724 27124
rect 378140 27072 378192 27124
rect 203340 27004 203392 27056
rect 415400 27004 415452 27056
rect 151912 26936 151964 26988
rect 183008 26936 183060 26988
rect 214288 26936 214340 26988
rect 560300 26936 560352 26988
rect 135260 26868 135312 26920
rect 181536 26868 181588 26920
rect 215668 26868 215720 26920
rect 572812 26868 572864 26920
rect 3424 25712 3476 25764
rect 179880 25712 179932 25764
rect 196532 25712 196584 25764
rect 333980 25712 334032 25764
rect 3516 25644 3568 25696
rect 179788 25644 179840 25696
rect 185400 25644 185452 25696
rect 186780 25644 186832 25696
rect 199108 25644 199160 25696
rect 368480 25644 368532 25696
rect 3792 25576 3844 25628
rect 179696 25576 179748 25628
rect 200580 25576 200632 25628
rect 383660 25576 383712 25628
rect 3700 25508 3752 25560
rect 179236 25508 179288 25560
rect 213000 25508 213052 25560
rect 545120 25508 545172 25560
rect 3608 25440 3660 25492
rect 179144 25440 179196 25492
rect 24124 25372 24176 25424
rect 179972 25372 180024 25424
rect 89720 24760 89772 24812
rect 157800 24760 157852 24812
rect 95240 24692 95292 24744
rect 168288 24692 168340 24744
rect 81440 24624 81492 24676
rect 166908 24624 166960 24676
rect 71780 24556 71832 24608
rect 157616 24556 157668 24608
rect 64880 24488 64932 24540
rect 165252 24488 165304 24540
rect 60740 24420 60792 24472
rect 164976 24420 165028 24472
rect 195060 24420 195112 24472
rect 316040 24420 316092 24472
rect 57980 24352 58032 24404
rect 163596 24352 163648 24404
rect 199016 24352 199068 24404
rect 362960 24352 363012 24404
rect 46940 24284 46992 24336
rect 158628 24284 158680 24336
rect 200488 24284 200540 24336
rect 382372 24284 382424 24336
rect 45560 24216 45612 24268
rect 159640 24216 159692 24268
rect 208952 24216 209004 24268
rect 488540 24216 488592 24268
rect 38660 24148 38712 24200
rect 159732 24148 159784 24200
rect 214104 24148 214156 24200
rect 556252 24148 556304 24200
rect 35900 24080 35952 24132
rect 162584 24080 162636 24132
rect 214196 24080 214248 24132
rect 563060 24080 563112 24132
rect 107660 24012 107712 24064
rect 158536 24012 158588 24064
rect 120080 23944 120132 23996
rect 169024 23944 169076 23996
rect 110420 23876 110472 23928
rect 157708 23876 157760 23928
rect 193680 23332 193732 23384
rect 299480 23332 299532 23384
rect 196440 23264 196492 23316
rect 325700 23264 325752 23316
rect 197820 23196 197872 23248
rect 349160 23196 349212 23248
rect 201868 23128 201920 23180
rect 396080 23128 396132 23180
rect 201960 23060 202012 23112
rect 398840 23060 398892 23112
rect 204812 22992 204864 23044
rect 440332 22992 440384 23044
rect 85580 22924 85632 22976
rect 166264 22924 166316 22976
rect 210240 22924 210292 22976
rect 503720 22924 503772 22976
rect 31760 22856 31812 22908
rect 162124 22856 162176 22908
rect 210332 22856 210384 22908
rect 506480 22856 506532 22908
rect 13820 22788 13872 22840
rect 160560 22788 160612 22840
rect 211712 22788 211764 22840
rect 517520 22788 517572 22840
rect 9680 22720 9732 22772
rect 160652 22720 160704 22772
rect 179420 22720 179472 22772
rect 184388 22720 184440 22772
rect 185308 22720 185360 22772
rect 193680 22720 193732 22772
rect 214012 22720 214064 22772
rect 564532 22720 564584 22772
rect 121460 21700 121512 21752
rect 169116 21700 169168 21752
rect 78680 21632 78732 21684
rect 166172 21632 166224 21684
rect 190828 21632 190880 21684
rect 260840 21632 260892 21684
rect 53840 21564 53892 21616
rect 162860 21564 162912 21616
rect 258632 21564 258684 21616
rect 471980 21564 472032 21616
rect 49700 21496 49752 21548
rect 163412 21496 163464 21548
rect 204720 21496 204772 21548
rect 441620 21496 441672 21548
rect 15200 21428 15252 21480
rect 158444 21428 158496 21480
rect 211620 21428 211672 21480
rect 520280 21428 520332 21480
rect 4160 21360 4212 21412
rect 159548 21360 159600 21412
rect 212908 21360 212960 21412
rect 540980 21360 541032 21412
rect 3424 20612 3476 20664
rect 177580 20612 177632 20664
rect 190644 20544 190696 20596
rect 262220 20544 262272 20596
rect 169852 20476 169904 20528
rect 269764 20476 269816 20528
rect 253756 20408 253808 20460
rect 411260 20408 411312 20460
rect 200396 20340 200448 20392
rect 379520 20340 379572 20392
rect 259368 20272 259420 20324
rect 454040 20272 454092 20324
rect 122840 20204 122892 20256
rect 168932 20204 168984 20256
rect 203524 20204 203576 20256
rect 404360 20204 404412 20256
rect 102140 20136 102192 20188
rect 167644 20136 167696 20188
rect 205180 20136 205232 20188
rect 415492 20136 415544 20188
rect 82820 20068 82872 20120
rect 166080 20068 166132 20120
rect 203248 20068 203300 20120
rect 422300 20068 422352 20120
rect 67640 20000 67692 20052
rect 164884 20000 164936 20052
rect 204628 20000 204680 20052
rect 429200 20000 429252 20052
rect 34520 19932 34572 19984
rect 162032 19932 162084 19984
rect 186688 19932 186740 19984
rect 203524 19932 203576 19984
rect 206284 19932 206336 19984
rect 456800 19932 456852 19984
rect 192208 19184 192260 19236
rect 273260 19184 273312 19236
rect 192392 19116 192444 19168
rect 276020 19116 276072 19168
rect 192300 19048 192352 19100
rect 280160 19048 280212 19100
rect 193588 18980 193640 19032
rect 291200 18980 291252 19032
rect 193496 18912 193548 18964
rect 293960 18912 294012 18964
rect 194968 18844 195020 18896
rect 305000 18844 305052 18896
rect 69020 18776 69072 18828
rect 164700 18776 164752 18828
rect 196348 18776 196400 18828
rect 329840 18776 329892 18828
rect 69112 18708 69164 18760
rect 164792 18708 164844 18760
rect 206652 18708 206704 18760
rect 418160 18708 418212 18760
rect 11060 18640 11112 18692
rect 160376 18640 160428 18692
rect 215944 18640 215996 18692
rect 436100 18640 436152 18692
rect 6920 18572 6972 18624
rect 160468 18572 160520 18624
rect 260196 18572 260248 18624
rect 536840 18572 536892 18624
rect 255872 17892 255924 17944
rect 397460 17892 397512 17944
rect 210148 17824 210200 17876
rect 468484 17824 468536 17876
rect 207388 17756 207440 17808
rect 466460 17756 466512 17808
rect 207572 17688 207624 17740
rect 470600 17688 470652 17740
rect 207480 17620 207532 17672
rect 473360 17620 473412 17672
rect 211436 17552 211488 17604
rect 521660 17552 521712 17604
rect 126980 17484 127032 17536
rect 180248 17484 180300 17536
rect 211528 17484 211580 17536
rect 524420 17484 524472 17536
rect 125600 17416 125652 17468
rect 179604 17416 179656 17468
rect 211344 17416 211396 17468
rect 528560 17416 528612 17468
rect 60832 17348 60884 17400
rect 164608 17348 164660 17400
rect 212724 17348 212776 17400
rect 535460 17348 535512 17400
rect 51080 17280 51132 17332
rect 163320 17280 163372 17332
rect 212632 17280 212684 17332
rect 539692 17280 539744 17332
rect 33140 17212 33192 17264
rect 161940 17212 161992 17264
rect 212816 17212 212868 17264
rect 546500 17212 546552 17264
rect 194876 17144 194928 17196
rect 316132 17144 316184 17196
rect 202972 16328 203024 16380
rect 414296 16328 414348 16380
rect 203064 16260 203116 16312
rect 417424 16260 417476 16312
rect 116400 16192 116452 16244
rect 168840 16192 168892 16244
rect 203156 16192 203208 16244
rect 420920 16192 420972 16244
rect 104072 16124 104124 16176
rect 167368 16124 167420 16176
rect 204536 16124 204588 16176
rect 432052 16124 432104 16176
rect 102232 16056 102284 16108
rect 167460 16056 167512 16108
rect 204444 16056 204496 16108
rect 435088 16056 435140 16108
rect 98184 15988 98236 16040
rect 167552 15988 167604 16040
rect 204352 15988 204404 16040
rect 439136 15988 439188 16040
rect 28448 15920 28500 15972
rect 161848 15920 161900 15972
rect 208860 15920 208912 15972
rect 490012 15920 490064 15972
rect 2872 15852 2924 15904
rect 158720 15852 158772 15904
rect 189264 15852 189316 15904
rect 203984 15852 204036 15904
rect 210056 15852 210108 15904
rect 507216 15852 507268 15904
rect 202420 15104 202472 15156
rect 339500 15104 339552 15156
rect 196164 15036 196216 15088
rect 336280 15036 336332 15088
rect 197636 14968 197688 15020
rect 342904 14968 342956 15020
rect 197728 14900 197780 14952
rect 346952 14900 347004 14952
rect 259276 14832 259328 14884
rect 447416 14832 447468 14884
rect 206192 14764 206244 14816
rect 453304 14764 453356 14816
rect 206100 14696 206152 14748
rect 456892 14696 456944 14748
rect 114008 14628 114060 14680
rect 168748 14628 168800 14680
rect 207204 14628 207256 14680
rect 469864 14628 469916 14680
rect 87512 14560 87564 14612
rect 165896 14560 165948 14612
rect 207296 14560 207348 14612
rect 473452 14560 473504 14612
rect 80888 14492 80940 14544
rect 165988 14492 166040 14544
rect 207112 14492 207164 14544
rect 476488 14492 476540 14544
rect 13544 14424 13596 14476
rect 160284 14424 160336 14476
rect 212540 14424 212592 14476
rect 542728 14424 542780 14476
rect 197176 14356 197228 14408
rect 332692 14356 332744 14408
rect 196256 14288 196308 14340
rect 328736 14288 328788 14340
rect 114744 13268 114796 13320
rect 168656 13268 168708 13320
rect 192116 13268 192168 13320
rect 272432 13268 272484 13320
rect 63224 13200 63276 13252
rect 164516 13200 164568 13252
rect 259184 13200 259236 13252
rect 465172 13200 465224 13252
rect 30104 13132 30156 13184
rect 161664 13132 161716 13184
rect 209964 13132 210016 13184
rect 500592 13132 500644 13184
rect 26240 13064 26292 13116
rect 161756 13064 161808 13116
rect 215576 13064 215628 13116
rect 578608 13064 578660 13116
rect 185216 12384 185268 12436
rect 192024 12384 192076 12436
rect 253664 12384 253716 12436
rect 394240 12384 394292 12436
rect 203800 12316 203852 12368
rect 376024 12316 376076 12368
rect 200304 12248 200356 12300
rect 389456 12248 389508 12300
rect 205916 12180 205968 12232
rect 448612 12180 448664 12232
rect 206008 12112 206060 12164
rect 451648 12112 451700 12164
rect 205732 12044 205784 12096
rect 455696 12044 455748 12096
rect 128912 11976 128964 12028
rect 178960 11976 179012 12028
rect 205824 11976 205876 12028
rect 459192 11976 459244 12028
rect 99840 11908 99892 11960
rect 167276 11908 167328 11960
rect 207020 11908 207072 11960
rect 465816 11908 465868 11960
rect 77392 11840 77444 11892
rect 165804 11840 165856 11892
rect 208768 11840 208820 11892
rect 493048 11840 493100 11892
rect 53288 11772 53340 11824
rect 163228 11772 163280 11824
rect 166080 11772 166132 11824
rect 179052 11772 179104 11824
rect 211252 11772 211304 11824
rect 523776 11772 523828 11824
rect 8760 11704 8812 11756
rect 161020 11704 161072 11756
rect 176660 11704 176712 11756
rect 177856 11704 177908 11756
rect 211160 11704 211212 11756
rect 527824 11704 527876 11756
rect 143540 11636 143592 11688
rect 144736 11636 144788 11688
rect 192116 11636 192168 11688
rect 276112 11636 276164 11688
rect 182364 11432 182416 11484
rect 184204 11432 184256 11484
rect 192760 10548 192812 10600
rect 279056 10548 279108 10600
rect 118792 10480 118844 10532
rect 168564 10480 168616 10532
rect 194508 10480 194560 10532
rect 297272 10480 297324 10532
rect 100760 10412 100812 10464
rect 167184 10412 167236 10464
rect 201776 10412 201828 10464
rect 398932 10412 398984 10464
rect 97448 10344 97500 10396
rect 167828 10344 167880 10396
rect 187148 10344 187200 10396
rect 194600 10344 194652 10396
rect 208676 10344 208728 10396
rect 486424 10344 486476 10396
rect 86408 10276 86460 10328
rect 166448 10276 166500 10328
rect 186596 10276 186648 10328
rect 206192 10276 206244 10328
rect 215484 10276 215536 10328
rect 575112 10276 575164 10328
rect 197544 9596 197596 9648
rect 344560 9596 344612 9648
rect 253480 9528 253532 9580
rect 413100 9528 413152 9580
rect 198924 9460 198976 9512
rect 361120 9460 361172 9512
rect 188160 9392 188212 9444
rect 220452 9392 220504 9444
rect 253572 9392 253624 9444
rect 430856 9392 430908 9444
rect 189172 9324 189224 9376
rect 241704 9324 241756 9376
rect 253204 9324 253256 9376
rect 434444 9324 434496 9376
rect 200120 9256 200172 9308
rect 388260 9256 388312 9308
rect 200212 9188 200264 9240
rect 391848 9188 391900 9240
rect 202880 9120 202932 9172
rect 420184 9120 420236 9172
rect 119896 9052 119948 9104
rect 169208 9052 169260 9104
rect 206744 9052 206796 9104
rect 460388 9052 460440 9104
rect 71504 8984 71556 9036
rect 161480 8984 161532 9036
rect 208584 8984 208636 9036
rect 482836 8984 482888 9036
rect 45468 8916 45520 8968
rect 163136 8916 163188 8968
rect 208492 8916 208544 8968
rect 485228 8916 485280 8968
rect 253296 8848 253348 8900
rect 381176 8848 381228 8900
rect 194784 7964 194836 8016
rect 315028 7964 315080 8016
rect 197452 7896 197504 7948
rect 350448 7896 350500 7948
rect 84476 7828 84528 7880
rect 166356 7828 166408 7880
rect 197360 7828 197412 7880
rect 352840 7828 352892 7880
rect 64328 7760 64380 7812
rect 164424 7760 164476 7812
rect 198832 7760 198884 7812
rect 367008 7760 367060 7812
rect 59636 7692 59688 7744
rect 165436 7692 165488 7744
rect 201684 7692 201736 7744
rect 406016 7692 406068 7744
rect 48964 7624 49016 7676
rect 163044 7624 163096 7676
rect 209872 7624 209924 7676
rect 510068 7624 510120 7676
rect 27712 7556 27764 7608
rect 161572 7556 161624 7608
rect 215392 7556 215444 7608
rect 571524 7556 571576 7608
rect 3424 6808 3476 6860
rect 135996 6808 136048 6860
rect 187792 6808 187844 6860
rect 216864 6808 216916 6860
rect 269764 6808 269816 6860
rect 580172 6808 580224 6860
rect 187884 6740 187936 6792
rect 222752 6740 222804 6792
rect 256240 6740 256292 6792
rect 328000 6740 328052 6792
rect 191840 6672 191892 6724
rect 270040 6672 270092 6724
rect 187976 6604 188028 6656
rect 226432 6604 226484 6656
rect 256608 6604 256660 6656
rect 342168 6604 342220 6656
rect 193312 6536 193364 6588
rect 299664 6536 299716 6588
rect 194692 6468 194744 6520
rect 311440 6468 311492 6520
rect 188068 6400 188120 6452
rect 229836 6400 229888 6452
rect 256332 6400 256384 6452
rect 377680 6400 377732 6452
rect 162492 6332 162544 6384
rect 182916 6332 182968 6384
rect 201592 6332 201644 6384
rect 403624 6332 403676 6384
rect 105728 6264 105780 6316
rect 167736 6264 167788 6316
rect 204260 6264 204312 6316
rect 437940 6264 437992 6316
rect 66720 6196 66772 6248
rect 165068 6196 165120 6248
rect 209780 6196 209832 6248
rect 502984 6196 503036 6248
rect 52552 6128 52604 6180
rect 162952 6128 163004 6180
rect 213920 6128 213972 6180
rect 553768 6128 553820 6180
rect 256148 6060 256200 6112
rect 306748 6060 306800 6112
rect 253388 5992 253440 6044
rect 290188 5992 290240 6044
rect 185124 5516 185176 5568
rect 188528 5516 188580 5568
rect 195612 5108 195664 5160
rect 307944 5108 307996 5160
rect 195980 5040 196032 5092
rect 323308 5040 323360 5092
rect 18236 4972 18288 5024
rect 160928 4972 160980 5024
rect 198740 4972 198792 5024
rect 368204 4972 368256 5024
rect 44272 4904 44324 4956
rect 163596 4904 163648 4956
rect 201500 4904 201552 4956
rect 402520 4904 402572 4956
rect 31300 4836 31352 4888
rect 162308 4836 162360 4888
rect 208400 4836 208452 4888
rect 492312 4904 492364 4956
rect 160100 4768 160152 4820
rect 182732 4768 182784 4820
rect 215300 4768 215352 4820
rect 576308 4768 576360 4820
rect 276020 4156 276072 4208
rect 276756 4156 276808 4208
rect 284300 4156 284352 4208
rect 285036 4156 285088 4208
rect 124680 4088 124732 4140
rect 159364 4088 159416 4140
rect 168472 4088 168524 4140
rect 173164 4088 173216 4140
rect 189724 4088 189776 4140
rect 190828 4088 190880 4140
rect 193220 4088 193272 4140
rect 296076 4088 296128 4140
rect 92756 4020 92808 4072
rect 134800 4020 134852 4072
rect 190000 4020 190052 4072
rect 201500 4020 201552 4072
rect 259092 4020 259144 4072
rect 440240 4020 440292 4072
rect 89168 3952 89220 4004
rect 133144 3952 133196 4004
rect 191196 3952 191248 4004
rect 205088 3952 205140 4004
rect 258816 3952 258868 4004
rect 448520 3952 448572 4004
rect 462964 3952 463016 4004
rect 487620 3952 487672 4004
rect 57244 3884 57296 3936
rect 133236 3884 133288 3936
rect 134156 3884 134208 3936
rect 177396 3884 177448 3936
rect 186412 3884 186464 3936
rect 200304 3884 200356 3936
rect 213184 3884 213236 3936
rect 225144 3884 225196 3936
rect 260104 3884 260156 3936
rect 461584 3884 461636 3936
rect 468484 3884 468536 3936
rect 511264 3884 511316 3936
rect 25320 3816 25372 3868
rect 137284 3816 137336 3868
rect 150624 3816 150676 3868
rect 173256 3816 173308 3868
rect 186320 3816 186372 3868
rect 210976 3816 211028 3868
rect 258908 3816 258960 3868
rect 480536 3816 480588 3868
rect 43076 3748 43128 3800
rect 159456 3748 159508 3800
rect 186504 3748 186556 3800
rect 207388 3748 207440 3800
rect 207848 3748 207900 3800
rect 433248 3748 433300 3800
rect 479524 3748 479576 3800
rect 526628 3748 526680 3800
rect 11152 3680 11204 3732
rect 134524 3680 134576 3732
rect 136456 3680 136508 3732
rect 177488 3680 177540 3732
rect 188620 3680 188672 3732
rect 203892 3680 203944 3732
rect 203984 3680 204036 3732
rect 246396 3680 246448 3732
rect 259000 3680 259052 3732
rect 484032 3680 484084 3732
rect 6460 3612 6512 3664
rect 138664 3612 138716 3664
rect 142436 3612 142488 3664
rect 178776 3612 178828 3664
rect 188804 3612 188856 3664
rect 219256 3612 219308 3664
rect 224224 3612 224276 3664
rect 450084 3612 450136 3664
rect 450544 3612 450596 3664
rect 523040 3612 523092 3664
rect 24216 3544 24268 3596
rect 158168 3544 158220 3596
rect 164884 3544 164936 3596
rect 174544 3544 174596 3596
rect 184940 3544 184992 3596
rect 185860 3544 185912 3596
rect 189080 3544 189132 3596
rect 234620 3544 234672 3596
rect 258724 3544 258776 3596
rect 501788 3544 501840 3596
rect 514760 3544 514812 3596
rect 515588 3544 515640 3596
rect 531320 3544 531372 3596
rect 532148 3544 532200 3596
rect 539600 3544 539652 3596
rect 540428 3544 540480 3596
rect 17040 3476 17092 3528
rect 18604 3476 18656 3528
rect 19432 3476 19484 3528
rect 158076 3476 158128 3528
rect 161296 3476 161348 3528
rect 572 3408 624 3460
rect 157984 3408 158036 3460
rect 158904 3408 158956 3460
rect 60740 3340 60792 3392
rect 61660 3340 61712 3392
rect 77300 3340 77352 3392
rect 78220 3340 78272 3392
rect 102140 3340 102192 3392
rect 103336 3340 103388 3392
rect 106924 3340 106976 3392
rect 134616 3340 134668 3392
rect 117596 3272 117648 3324
rect 134708 3272 134760 3324
rect 168380 3408 168432 3460
rect 169576 3408 169628 3460
rect 173164 3476 173216 3528
rect 174636 3476 174688 3528
rect 189816 3476 189868 3528
rect 174268 3408 174320 3460
rect 178868 3408 178920 3460
rect 191472 3408 191524 3460
rect 211804 3476 211856 3528
rect 213368 3476 213420 3528
rect 217324 3476 217376 3528
rect 177304 3340 177356 3392
rect 188436 3340 188488 3392
rect 178684 3272 178736 3324
rect 184848 3272 184900 3324
rect 189724 3272 189776 3324
rect 191104 3340 191156 3392
rect 202696 3340 202748 3392
rect 199108 3272 199160 3324
rect 190092 3204 190144 3256
rect 197912 3204 197964 3256
rect 215668 3408 215720 3460
rect 226340 3408 226392 3460
rect 227536 3408 227588 3460
rect 210424 3340 210476 3392
rect 212172 3340 212224 3392
rect 251180 3408 251232 3460
rect 252376 3408 252428 3460
rect 256056 3408 256108 3460
rect 257068 3340 257120 3392
rect 271144 3408 271196 3460
rect 292580 3340 292632 3392
rect 299480 3340 299532 3392
rect 300768 3340 300820 3392
rect 307760 3340 307812 3392
rect 309048 3340 309100 3392
rect 316040 3340 316092 3392
rect 317328 3340 317380 3392
rect 324412 3340 324464 3392
rect 325608 3340 325660 3392
rect 332600 3340 332652 3392
rect 333888 3340 333940 3392
rect 357440 3340 357492 3392
rect 358728 3340 358780 3392
rect 374000 3340 374052 3392
rect 375288 3340 375340 3392
rect 382280 3340 382332 3392
rect 383568 3340 383620 3392
rect 398932 3340 398984 3392
rect 400128 3340 400180 3392
rect 407212 3340 407264 3392
rect 408408 3340 408460 3392
rect 415400 3340 415452 3392
rect 416688 3340 416740 3392
rect 423680 3340 423732 3392
rect 424968 3340 425020 3392
rect 440332 3340 440384 3392
rect 441528 3340 441580 3392
rect 448612 3340 448664 3392
rect 449808 3340 449860 3392
rect 456800 3340 456852 3392
rect 458088 3340 458140 3392
rect 256424 3272 256476 3324
rect 288992 3272 289044 3324
rect 473360 3476 473412 3528
rect 474188 3476 474240 3528
rect 487804 3476 487856 3528
rect 556160 3476 556212 3528
rect 572720 3476 572772 3528
rect 573548 3476 573600 3528
rect 479340 3340 479392 3392
rect 583392 3408 583444 3460
rect 489920 3340 489972 3392
rect 490748 3340 490800 3392
rect 255964 3204 256016 3256
rect 274824 3204 274876 3256
rect 189908 3136 189960 3188
rect 193220 3136 193272 3188
rect 203524 3136 203576 3188
rect 208584 3136 208636 3188
rect 256516 3136 256568 3188
rect 271236 3136 271288 3188
rect 132960 3068 133012 3120
rect 135904 3068 135956 3120
rect 214472 2864 214524 2916
rect 216680 2864 216732 2916
rect 207020 2796 207072 2848
rect 209780 2796 209832 2848
rect 450084 2796 450136 2848
rect 450912 2796 450964 2848
<< metal2 >>
rect 6932 703582 7972 703610
rect 3422 684312 3478 684321
rect 3422 684247 3478 684256
rect 3436 683194 3464 684247
rect 3424 683188 3476 683194
rect 3424 683130 3476 683136
rect 3514 671256 3570 671265
rect 3514 671191 3570 671200
rect 3528 670750 3556 671191
rect 3516 670744 3568 670750
rect 3516 670686 3568 670692
rect 3422 658200 3478 658209
rect 3422 658135 3478 658144
rect 3436 656946 3464 658135
rect 3424 656940 3476 656946
rect 3424 656882 3476 656888
rect 3424 632120 3476 632126
rect 3422 632088 3424 632097
rect 3476 632088 3478 632097
rect 3422 632023 3478 632032
rect 3146 619168 3202 619177
rect 3146 619103 3202 619112
rect 3160 618322 3188 619103
rect 3148 618316 3200 618322
rect 3148 618258 3200 618264
rect 3238 606112 3294 606121
rect 3238 606047 3294 606056
rect 3252 605878 3280 606047
rect 3240 605872 3292 605878
rect 3240 605814 3292 605820
rect 3330 580000 3386 580009
rect 3330 579935 3386 579944
rect 3344 579698 3372 579935
rect 3332 579692 3384 579698
rect 3332 579634 3384 579640
rect 3422 566944 3478 566953
rect 3422 566879 3478 566888
rect 3436 565894 3464 566879
rect 3424 565888 3476 565894
rect 3424 565830 3476 565836
rect 3422 553888 3478 553897
rect 3422 553823 3478 553832
rect 2962 527912 3018 527921
rect 2962 527847 3018 527856
rect 2976 527202 3004 527847
rect 2964 527196 3016 527202
rect 2964 527138 3016 527144
rect 3330 423600 3386 423609
rect 3330 423535 3386 423544
rect 3344 422346 3372 423535
rect 3332 422340 3384 422346
rect 3332 422282 3384 422288
rect 3330 410544 3386 410553
rect 3330 410479 3386 410488
rect 3344 409902 3372 410479
rect 3332 409896 3384 409902
rect 3332 409838 3384 409844
rect 3332 397520 3384 397526
rect 3330 397488 3332 397497
rect 3384 397488 3386 397497
rect 3330 397423 3386 397432
rect 3330 371376 3386 371385
rect 3330 371311 3386 371320
rect 3344 371278 3372 371311
rect 3332 371272 3384 371278
rect 3332 371214 3384 371220
rect 2962 358456 3018 358465
rect 2962 358391 3018 358400
rect 2976 357474 3004 358391
rect 2964 357468 3016 357474
rect 2964 357410 3016 357416
rect 3054 345400 3110 345409
rect 3054 345335 3110 345344
rect 3068 345098 3096 345335
rect 3056 345092 3108 345098
rect 3056 345034 3108 345040
rect 3436 327758 3464 553823
rect 3514 514856 3570 514865
rect 3514 514791 3516 514800
rect 3568 514791 3570 514800
rect 3516 514762 3568 514768
rect 3514 501800 3570 501809
rect 3514 501735 3570 501744
rect 3424 327752 3476 327758
rect 3424 327694 3476 327700
rect 3528 324970 3556 501735
rect 3606 475688 3662 475697
rect 3606 475623 3662 475632
rect 3516 324964 3568 324970
rect 3516 324906 3568 324912
rect 3620 323610 3648 475623
rect 3698 462632 3754 462641
rect 3698 462567 3754 462576
rect 3608 323604 3660 323610
rect 3608 323546 3660 323552
rect 3712 322250 3740 462567
rect 3790 449576 3846 449585
rect 3790 449511 3846 449520
rect 3804 322318 3832 449511
rect 3792 322312 3844 322318
rect 3792 322254 3844 322260
rect 3700 322244 3752 322250
rect 3700 322186 3752 322192
rect 3422 319288 3478 319297
rect 3422 319223 3478 319232
rect 3436 318850 3464 319223
rect 3424 318844 3476 318850
rect 3424 318786 3476 318792
rect 3238 306232 3294 306241
rect 3238 306167 3294 306176
rect 3252 305046 3280 306167
rect 3240 305040 3292 305046
rect 3240 304982 3292 304988
rect 3422 293176 3478 293185
rect 3422 293111 3478 293120
rect 3054 267200 3110 267209
rect 3054 267135 3110 267144
rect 3068 266422 3096 267135
rect 3056 266416 3108 266422
rect 3056 266358 3108 266364
rect 3330 214976 3386 214985
rect 3330 214911 3386 214920
rect 3344 213994 3372 214911
rect 3332 213988 3384 213994
rect 3332 213930 3384 213936
rect 3238 201920 3294 201929
rect 3238 201855 3294 201864
rect 3252 201550 3280 201855
rect 3240 201544 3292 201550
rect 3240 201486 3292 201492
rect 3330 162888 3386 162897
rect 3330 162823 3386 162832
rect 3344 160750 3372 162823
rect 3436 160818 3464 293111
rect 3514 254144 3570 254153
rect 3514 254079 3570 254088
rect 3528 253978 3556 254079
rect 3516 253972 3568 253978
rect 3516 253914 3568 253920
rect 3514 241088 3570 241097
rect 3514 241023 3570 241032
rect 3424 160812 3476 160818
rect 3424 160754 3476 160760
rect 3332 160744 3384 160750
rect 3332 160686 3384 160692
rect 3528 158030 3556 241023
rect 3606 188864 3662 188873
rect 3606 188799 3662 188808
rect 3620 159390 3648 188799
rect 3608 159384 3660 159390
rect 3608 159326 3660 159332
rect 3516 158024 3568 158030
rect 3516 157966 3568 157972
rect 3422 149832 3478 149841
rect 3422 149767 3478 149776
rect 3436 149122 3464 149767
rect 3424 149116 3476 149122
rect 3424 149058 3476 149064
rect 3422 136776 3478 136785
rect 3422 136711 3478 136720
rect 3436 136678 3464 136711
rect 3424 136672 3476 136678
rect 3424 136614 3476 136620
rect 6932 133210 6960 703582
rect 7944 703474 7972 703582
rect 8086 703520 8198 704960
rect 24278 703520 24390 704960
rect 40470 703520 40582 704960
rect 56754 703520 56866 704960
rect 72946 703520 73058 704960
rect 89138 703520 89250 704960
rect 105422 703520 105534 704960
rect 121614 703520 121726 704960
rect 136652 703582 137692 703610
rect 8128 703474 8156 703520
rect 7944 703446 8156 703474
rect 24320 700398 24348 703520
rect 24308 700392 24360 700398
rect 24308 700334 24360 700340
rect 40512 700330 40540 703520
rect 72988 700466 73016 703520
rect 89180 700534 89208 703520
rect 105464 700602 105492 703520
rect 105452 700596 105504 700602
rect 105452 700538 105504 700544
rect 89168 700528 89220 700534
rect 89168 700470 89220 700476
rect 72976 700460 73028 700466
rect 72976 700402 73028 700408
rect 40500 700324 40552 700330
rect 40500 700266 40552 700272
rect 135904 605872 135956 605878
rect 135904 605814 135956 605820
rect 111890 591696 111946 591705
rect 111890 591631 111946 591640
rect 111798 591016 111854 591025
rect 111798 590951 111854 590960
rect 111812 590782 111840 590951
rect 111800 590776 111852 590782
rect 111800 590718 111852 590724
rect 111904 590714 111932 591631
rect 119620 590776 119672 590782
rect 119620 590718 119672 590724
rect 111892 590708 111944 590714
rect 111892 590650 111944 590656
rect 111890 590336 111946 590345
rect 111890 590271 111946 590280
rect 111798 589656 111854 589665
rect 111798 589591 111854 589600
rect 111812 589422 111840 589591
rect 111800 589416 111852 589422
rect 111800 589358 111852 589364
rect 111904 589354 111932 590271
rect 111892 589348 111944 589354
rect 111892 589290 111944 589296
rect 111798 588976 111854 588985
rect 111798 588911 111854 588920
rect 111812 587926 111840 588911
rect 112258 588296 112314 588305
rect 112258 588231 112314 588240
rect 111800 587920 111852 587926
rect 111800 587862 111852 587868
rect 111798 587616 111854 587625
rect 111798 587551 111854 587560
rect 111812 586566 111840 587551
rect 111800 586560 111852 586566
rect 111800 586502 111852 586508
rect 111798 586256 111854 586265
rect 111798 586191 111854 586200
rect 111812 585410 111840 586191
rect 112272 585818 112300 588231
rect 112718 586936 112774 586945
rect 112718 586871 112774 586880
rect 112260 585812 112312 585818
rect 112260 585754 112312 585760
rect 111982 585576 112038 585585
rect 111982 585511 112038 585520
rect 111800 585404 111852 585410
rect 111800 585346 111852 585352
rect 111890 584896 111946 584905
rect 111890 584831 111946 584840
rect 111798 584216 111854 584225
rect 111798 584151 111854 584160
rect 111812 583778 111840 584151
rect 111904 583914 111932 584831
rect 111996 584458 112024 585511
rect 111984 584452 112036 584458
rect 111984 584394 112036 584400
rect 111892 583908 111944 583914
rect 111892 583850 111944 583856
rect 111800 583772 111852 583778
rect 111800 583714 111852 583720
rect 111798 583536 111854 583545
rect 111798 583471 111854 583480
rect 111812 582418 111840 583471
rect 111890 582856 111946 582865
rect 111890 582791 111946 582800
rect 111800 582412 111852 582418
rect 111800 582354 111852 582360
rect 111798 582176 111854 582185
rect 111798 582111 111854 582120
rect 111812 581058 111840 582111
rect 111904 581670 111932 582791
rect 111892 581664 111944 581670
rect 111892 581606 111944 581612
rect 111982 581496 112038 581505
rect 111982 581431 112038 581440
rect 111800 581052 111852 581058
rect 111800 580994 111852 581000
rect 111890 580816 111946 580825
rect 111890 580751 111946 580760
rect 111798 580136 111854 580145
rect 111798 580071 111854 580080
rect 111812 579698 111840 580071
rect 111904 579766 111932 580751
rect 111996 580310 112024 581431
rect 111984 580304 112036 580310
rect 111984 580246 112036 580252
rect 111892 579760 111944 579766
rect 111892 579702 111944 579708
rect 29644 579692 29696 579698
rect 29644 579634 29696 579640
rect 111800 579692 111852 579698
rect 111800 579634 111852 579640
rect 26884 253972 26936 253978
rect 26884 253914 26936 253920
rect 26896 133414 26924 253914
rect 29552 201544 29604 201550
rect 29552 201486 29604 201492
rect 29564 133754 29592 201486
rect 29552 133748 29604 133754
rect 29552 133690 29604 133696
rect 26884 133408 26936 133414
rect 26884 133350 26936 133356
rect 29656 133278 29684 579634
rect 111890 579456 111946 579465
rect 111890 579391 111946 579400
rect 111798 578776 111854 578785
rect 111798 578711 111854 578720
rect 111812 578338 111840 578711
rect 111800 578332 111852 578338
rect 111800 578274 111852 578280
rect 111904 578270 111932 579391
rect 111892 578264 111944 578270
rect 111892 578206 111944 578212
rect 111798 578096 111854 578105
rect 111798 578031 111854 578040
rect 111812 576910 111840 578031
rect 112442 577416 112498 577425
rect 112442 577351 112498 577360
rect 111800 576904 111852 576910
rect 111800 576846 111852 576852
rect 111890 576736 111946 576745
rect 111890 576671 111946 576680
rect 111798 576056 111854 576065
rect 111798 575991 111854 576000
rect 111812 575550 111840 575991
rect 111904 575618 111932 576671
rect 111892 575612 111944 575618
rect 111892 575554 111944 575560
rect 111800 575544 111852 575550
rect 111800 575486 111852 575492
rect 111890 575376 111946 575385
rect 111890 575311 111946 575320
rect 111798 574696 111854 574705
rect 111798 574631 111854 574640
rect 111812 574122 111840 574631
rect 111904 574394 111932 575311
rect 111892 574388 111944 574394
rect 111892 574330 111944 574336
rect 111800 574116 111852 574122
rect 111800 574058 111852 574064
rect 111890 574016 111946 574025
rect 111890 573951 111946 573960
rect 111798 573336 111854 573345
rect 111798 573271 111854 573280
rect 111812 572830 111840 573271
rect 111800 572824 111852 572830
rect 111800 572766 111852 572772
rect 111904 572762 111932 573951
rect 111892 572756 111944 572762
rect 111892 572698 111944 572704
rect 111890 572656 111946 572665
rect 111890 572591 111946 572600
rect 111798 571976 111854 571985
rect 111798 571911 111854 571920
rect 111812 571470 111840 571911
rect 111800 571464 111852 571470
rect 111800 571406 111852 571412
rect 111904 571402 111932 572591
rect 111892 571396 111944 571402
rect 111892 571338 111944 571344
rect 111982 571296 112038 571305
rect 111982 571231 112038 571240
rect 111798 570616 111854 570625
rect 111798 570551 111854 570560
rect 111812 570042 111840 570551
rect 111800 570036 111852 570042
rect 111800 569978 111852 569984
rect 111996 569974 112024 571231
rect 111984 569968 112036 569974
rect 111890 569936 111946 569945
rect 111984 569910 112036 569916
rect 111890 569871 111946 569880
rect 111798 569256 111854 569265
rect 111798 569191 111854 569200
rect 111812 568614 111840 569191
rect 111904 568682 111932 569871
rect 111892 568676 111944 568682
rect 111892 568618 111944 568624
rect 111800 568608 111852 568614
rect 111800 568550 111852 568556
rect 111982 568576 112038 568585
rect 111982 568511 112038 568520
rect 111800 567248 111852 567254
rect 111798 567216 111800 567225
rect 111852 567216 111854 567225
rect 111798 567151 111854 567160
rect 111890 566536 111946 566545
rect 111890 566471 111946 566480
rect 111800 565956 111852 565962
rect 111800 565898 111852 565904
rect 29736 565888 29788 565894
rect 111812 565865 111840 565898
rect 111904 565894 111932 566471
rect 111892 565888 111944 565894
rect 29736 565830 29788 565836
rect 111798 565856 111854 565865
rect 29748 133550 29776 565830
rect 111892 565830 111944 565836
rect 111798 565791 111854 565800
rect 111890 565176 111946 565185
rect 111890 565111 111946 565120
rect 111800 564528 111852 564534
rect 111798 564496 111800 564505
rect 111852 564496 111854 564505
rect 111904 564466 111932 565111
rect 111798 564431 111854 564440
rect 111892 564460 111944 564466
rect 111892 564402 111944 564408
rect 111798 563136 111854 563145
rect 111798 563071 111800 563080
rect 111852 563071 111854 563080
rect 111800 563042 111852 563048
rect 111996 562358 112024 568511
rect 112350 567896 112406 567905
rect 112350 567831 112406 567840
rect 111984 562352 112036 562358
rect 111984 562294 112036 562300
rect 112364 562306 112392 567831
rect 112456 563718 112484 577351
rect 112444 563712 112496 563718
rect 112444 563654 112496 563660
rect 112626 562456 112682 562465
rect 112626 562391 112682 562400
rect 112364 562278 112576 562306
rect 111798 561776 111854 561785
rect 111798 561711 111800 561720
rect 111852 561711 111854 561720
rect 111800 561682 111852 561688
rect 112442 561096 112498 561105
rect 112442 561031 112498 561040
rect 111798 560416 111854 560425
rect 111798 560351 111854 560360
rect 111812 560318 111840 560351
rect 111800 560312 111852 560318
rect 111800 560254 111852 560260
rect 111890 559736 111946 559745
rect 111890 559671 111946 559680
rect 111798 559056 111854 559065
rect 111798 558991 111800 559000
rect 111852 558991 111854 559000
rect 111800 558962 111852 558968
rect 111904 558958 111932 559671
rect 111892 558952 111944 558958
rect 111892 558894 111944 558900
rect 111890 558376 111946 558385
rect 111890 558311 111946 558320
rect 111798 557696 111854 557705
rect 111798 557631 111800 557640
rect 111852 557631 111854 557640
rect 111800 557602 111852 557608
rect 111904 557598 111932 558311
rect 111892 557592 111944 557598
rect 111892 557534 111944 557540
rect 111798 557016 111854 557025
rect 111798 556951 111854 556960
rect 111812 556238 111840 556951
rect 111982 556336 112038 556345
rect 111982 556271 112038 556280
rect 111800 556232 111852 556238
rect 111800 556174 111852 556180
rect 111890 555656 111946 555665
rect 111890 555591 111946 555600
rect 111798 554976 111854 554985
rect 111798 554911 111800 554920
rect 111852 554911 111854 554920
rect 111800 554882 111852 554888
rect 111904 554810 111932 555591
rect 111892 554804 111944 554810
rect 111892 554746 111944 554752
rect 111996 554062 112024 556271
rect 112074 554296 112130 554305
rect 112074 554231 112130 554240
rect 111984 554056 112036 554062
rect 111984 553998 112036 554004
rect 111798 553616 111854 553625
rect 111798 553551 111854 553560
rect 111812 553450 111840 553551
rect 111800 553444 111852 553450
rect 111800 553386 111852 553392
rect 111890 552936 111946 552945
rect 111890 552871 111946 552880
rect 111798 552256 111854 552265
rect 111798 552191 111854 552200
rect 111812 552090 111840 552191
rect 111904 552158 111932 552871
rect 111892 552152 111944 552158
rect 111892 552094 111944 552100
rect 111800 552084 111852 552090
rect 111800 552026 111852 552032
rect 111890 551576 111946 551585
rect 111890 551511 111946 551520
rect 111798 550896 111854 550905
rect 111798 550831 111854 550840
rect 111812 550730 111840 550831
rect 111800 550724 111852 550730
rect 111800 550666 111852 550672
rect 111904 550662 111932 551511
rect 111892 550656 111944 550662
rect 111892 550598 111944 550604
rect 111890 550216 111946 550225
rect 111890 550151 111946 550160
rect 111798 549536 111854 549545
rect 111798 549471 111854 549480
rect 111812 549370 111840 549471
rect 111800 549364 111852 549370
rect 111800 549306 111852 549312
rect 111904 549302 111932 550151
rect 111892 549296 111944 549302
rect 111892 549238 111944 549244
rect 111890 548856 111946 548865
rect 111890 548791 111946 548800
rect 111798 548176 111854 548185
rect 111798 548111 111800 548120
rect 111852 548111 111854 548120
rect 111800 548082 111852 548088
rect 111904 547942 111932 548791
rect 112088 548554 112116 554231
rect 112076 548548 112128 548554
rect 112076 548490 112128 548496
rect 111892 547936 111944 547942
rect 111892 547878 111944 547884
rect 111798 546816 111854 546825
rect 111798 546751 111854 546760
rect 111812 546514 111840 546751
rect 111800 546508 111852 546514
rect 111800 546450 111852 546456
rect 111890 546136 111946 546145
rect 111890 546071 111946 546080
rect 111798 545456 111854 545465
rect 111798 545391 111854 545400
rect 111812 545154 111840 545391
rect 111904 545222 111932 546071
rect 111892 545216 111944 545222
rect 111892 545158 111944 545164
rect 111800 545148 111852 545154
rect 111800 545090 111852 545096
rect 111798 544096 111854 544105
rect 111798 544031 111854 544040
rect 111812 543794 111840 544031
rect 111800 543788 111852 543794
rect 111800 543730 111852 543736
rect 111890 543416 111946 543425
rect 111890 543351 111946 543360
rect 111798 542736 111854 542745
rect 111798 542671 111854 542680
rect 111812 542434 111840 542671
rect 111904 542502 111932 543351
rect 111892 542496 111944 542502
rect 111892 542438 111944 542444
rect 111800 542428 111852 542434
rect 111800 542370 111852 542376
rect 111798 542056 111854 542065
rect 111798 541991 111854 542000
rect 111812 541006 111840 541991
rect 111800 541000 111852 541006
rect 111800 540942 111852 540948
rect 112350 540696 112406 540705
rect 112350 540631 112406 540640
rect 111798 540016 111854 540025
rect 111798 539951 111854 539960
rect 111812 539646 111840 539951
rect 111800 539640 111852 539646
rect 111800 539582 111852 539588
rect 111890 539336 111946 539345
rect 111890 539271 111946 539280
rect 111798 538656 111854 538665
rect 111798 538591 111854 538600
rect 111812 538354 111840 538591
rect 111800 538348 111852 538354
rect 111800 538290 111852 538296
rect 111904 538286 111932 539271
rect 111892 538280 111944 538286
rect 111892 538222 111944 538228
rect 111890 537976 111946 537985
rect 111890 537911 111946 537920
rect 111798 537296 111854 537305
rect 111798 537231 111854 537240
rect 111812 536926 111840 537231
rect 111800 536920 111852 536926
rect 111800 536862 111852 536868
rect 111904 536858 111932 537911
rect 111892 536852 111944 536858
rect 111892 536794 111944 536800
rect 111890 536616 111946 536625
rect 111890 536551 111946 536560
rect 111798 535936 111854 535945
rect 111798 535871 111854 535880
rect 111812 535498 111840 535871
rect 111904 535566 111932 536551
rect 111892 535560 111944 535566
rect 111892 535502 111944 535508
rect 111800 535492 111852 535498
rect 111800 535434 111852 535440
rect 111798 535256 111854 535265
rect 111798 535191 111854 535200
rect 111812 534138 111840 535191
rect 111890 534576 111946 534585
rect 111890 534511 111946 534520
rect 111800 534132 111852 534138
rect 111800 534074 111852 534080
rect 111904 533798 111932 534511
rect 111892 533792 111944 533798
rect 111892 533734 111944 533740
rect 112258 532536 112314 532545
rect 112258 532471 112314 532480
rect 112272 531350 112300 532471
rect 112260 531344 112312 531350
rect 112260 531286 112312 531292
rect 112260 531208 112312 531214
rect 112260 531150 112312 531156
rect 112272 529242 112300 531150
rect 112364 529938 112392 540631
rect 112456 530058 112484 561031
rect 112548 552702 112576 562278
rect 112640 556850 112668 562391
rect 112628 556844 112680 556850
rect 112628 556786 112680 556792
rect 112536 552696 112588 552702
rect 112536 552638 112588 552644
rect 112732 534074 112760 586871
rect 113824 585404 113876 585410
rect 113824 585346 113876 585352
rect 112994 563816 113050 563825
rect 112994 563751 113050 563760
rect 112810 547496 112866 547505
rect 112810 547431 112866 547440
rect 112640 534046 112760 534074
rect 112640 531214 112668 534046
rect 112718 533896 112774 533905
rect 112718 533831 112774 533840
rect 112628 531208 112680 531214
rect 112628 531150 112680 531156
rect 112626 530496 112682 530505
rect 112626 530431 112682 530440
rect 112444 530052 112496 530058
rect 112444 529994 112496 530000
rect 112640 529990 112668 530431
rect 112628 529984 112680 529990
rect 112364 529910 112576 529938
rect 112628 529926 112680 529932
rect 112444 529848 112496 529854
rect 112350 529816 112406 529825
rect 112444 529790 112496 529796
rect 112350 529751 112406 529760
rect 112260 529236 112312 529242
rect 112260 529178 112312 529184
rect 112364 528630 112392 529751
rect 112352 528624 112404 528630
rect 112352 528566 112404 528572
rect 111798 528456 111854 528465
rect 111798 528391 111854 528400
rect 111812 527270 111840 528391
rect 112258 527776 112314 527785
rect 112258 527711 112314 527720
rect 111800 527264 111852 527270
rect 111800 527206 111852 527212
rect 29828 527196 29880 527202
rect 29828 527138 29880 527144
rect 29736 133544 29788 133550
rect 29736 133486 29788 133492
rect 29840 133346 29868 527138
rect 112272 525774 112300 527711
rect 112350 527096 112406 527105
rect 112350 527031 112406 527040
rect 112364 525910 112392 527031
rect 112352 525904 112404 525910
rect 112352 525846 112404 525852
rect 112260 525768 112312 525774
rect 112074 525736 112130 525745
rect 112260 525710 112312 525716
rect 112074 525671 112130 525680
rect 112088 524482 112116 525671
rect 112076 524476 112128 524482
rect 112076 524418 112128 524424
rect 111890 524376 111946 524385
rect 111890 524311 111946 524320
rect 111798 523696 111854 523705
rect 111798 523631 111854 523640
rect 111812 523054 111840 523631
rect 111904 523122 111932 524311
rect 111892 523116 111944 523122
rect 111892 523058 111944 523064
rect 111800 523048 111852 523054
rect 111800 522990 111852 522996
rect 111890 523016 111946 523025
rect 111890 522951 111946 522960
rect 111798 522336 111854 522345
rect 111798 522271 111854 522280
rect 111812 521694 111840 522271
rect 111904 521762 111932 522951
rect 111892 521756 111944 521762
rect 111892 521698 111944 521704
rect 111800 521688 111852 521694
rect 111800 521630 111852 521636
rect 111890 521656 111946 521665
rect 111890 521591 111946 521600
rect 111798 520976 111854 520985
rect 111798 520911 111854 520920
rect 111812 520402 111840 520911
rect 111800 520396 111852 520402
rect 111800 520338 111852 520344
rect 111904 520334 111932 521591
rect 111892 520328 111944 520334
rect 111798 520296 111854 520305
rect 111892 520270 111944 520276
rect 111798 520231 111854 520240
rect 111812 519654 111840 520231
rect 111800 519648 111852 519654
rect 111800 519590 111852 519596
rect 112350 519616 112406 519625
rect 112350 519551 112406 519560
rect 112258 518936 112314 518945
rect 112258 518871 112314 518880
rect 111798 517576 111854 517585
rect 111798 517511 111800 517520
rect 111852 517511 111854 517520
rect 111800 517482 111852 517488
rect 111890 516896 111946 516905
rect 111890 516831 111946 516840
rect 111904 516254 111932 516831
rect 111892 516248 111944 516254
rect 111798 516216 111854 516225
rect 111892 516190 111944 516196
rect 111798 516151 111800 516160
rect 111852 516151 111854 516160
rect 111800 516122 111852 516128
rect 111890 515536 111946 515545
rect 111890 515471 111946 515480
rect 111800 514888 111852 514894
rect 111798 514856 111800 514865
rect 111852 514856 111854 514865
rect 29920 514820 29972 514826
rect 111904 514826 111932 515471
rect 111798 514791 111854 514800
rect 111892 514820 111944 514826
rect 29920 514762 29972 514768
rect 111892 514762 111944 514768
rect 29932 133822 29960 514762
rect 111890 514176 111946 514185
rect 111890 514111 111946 514120
rect 111798 513496 111854 513505
rect 111798 513431 111800 513440
rect 111852 513431 111854 513440
rect 111800 513402 111852 513408
rect 111904 513398 111932 514111
rect 111892 513392 111944 513398
rect 111892 513334 111944 513340
rect 111982 512816 112038 512825
rect 111982 512751 112038 512760
rect 111798 512136 111854 512145
rect 111798 512071 111854 512080
rect 111812 512038 111840 512071
rect 111800 512032 111852 512038
rect 111800 511974 111852 511980
rect 111890 511456 111946 511465
rect 111890 511391 111946 511400
rect 111798 510776 111854 510785
rect 111904 510746 111932 511391
rect 111798 510711 111854 510720
rect 111892 510740 111944 510746
rect 111812 510678 111840 510711
rect 111892 510682 111944 510688
rect 111800 510672 111852 510678
rect 111800 510614 111852 510620
rect 111996 509930 112024 512751
rect 112272 512650 112300 518871
rect 112364 518226 112392 519551
rect 112352 518220 112404 518226
rect 112352 518162 112404 518168
rect 112260 512644 112312 512650
rect 112260 512586 112312 512592
rect 111984 509924 112036 509930
rect 111984 509866 112036 509872
rect 111798 509416 111854 509425
rect 111798 509351 111854 509360
rect 111812 509318 111840 509351
rect 111800 509312 111852 509318
rect 111800 509254 111852 509260
rect 111890 508736 111946 508745
rect 111890 508671 111946 508680
rect 111798 508056 111854 508065
rect 111798 507991 111854 508000
rect 111812 507890 111840 507991
rect 111904 507958 111932 508671
rect 111892 507952 111944 507958
rect 111892 507894 111944 507900
rect 111800 507884 111852 507890
rect 111800 507826 111852 507832
rect 111798 507376 111854 507385
rect 111798 507311 111854 507320
rect 111812 506530 111840 507311
rect 111890 506696 111946 506705
rect 111890 506631 111946 506640
rect 111800 506524 111852 506530
rect 111800 506466 111852 506472
rect 111798 506016 111854 506025
rect 111798 505951 111854 505960
rect 111812 505170 111840 505951
rect 111904 505782 111932 506631
rect 111892 505776 111944 505782
rect 111892 505718 111944 505724
rect 112350 505336 112406 505345
rect 112350 505271 112406 505280
rect 111800 505164 111852 505170
rect 111800 505106 111852 505112
rect 111890 504656 111946 504665
rect 111890 504591 111946 504600
rect 111798 503976 111854 503985
rect 111798 503911 111800 503920
rect 111852 503911 111854 503920
rect 111800 503882 111852 503888
rect 111904 503742 111932 504591
rect 111892 503736 111944 503742
rect 111892 503678 111944 503684
rect 111890 503296 111946 503305
rect 111890 503231 111946 503240
rect 111798 502616 111854 502625
rect 111798 502551 111854 502560
rect 111812 502450 111840 502551
rect 111800 502444 111852 502450
rect 111800 502386 111852 502392
rect 111904 502382 111932 503231
rect 111892 502376 111944 502382
rect 111892 502318 111944 502324
rect 111798 501936 111854 501945
rect 111798 501871 111854 501880
rect 111812 501022 111840 501871
rect 111890 501256 111946 501265
rect 111890 501191 111946 501200
rect 111800 501016 111852 501022
rect 111800 500958 111852 500964
rect 111798 499896 111854 499905
rect 111798 499831 111854 499840
rect 111812 499730 111840 499831
rect 111800 499724 111852 499730
rect 111800 499666 111852 499672
rect 111904 498846 111932 501191
rect 111982 500576 112038 500585
rect 111982 500511 112038 500520
rect 111996 499594 112024 500511
rect 111984 499588 112036 499594
rect 111984 499530 112036 499536
rect 111982 499216 112038 499225
rect 111982 499151 112038 499160
rect 111892 498840 111944 498846
rect 111892 498782 111944 498788
rect 111798 498536 111854 498545
rect 111798 498471 111854 498480
rect 111812 498234 111840 498471
rect 111800 498228 111852 498234
rect 111800 498170 111852 498176
rect 111890 497856 111946 497865
rect 111890 497791 111946 497800
rect 111798 497176 111854 497185
rect 111798 497111 111854 497120
rect 111812 496942 111840 497111
rect 111800 496936 111852 496942
rect 111800 496878 111852 496884
rect 111904 496874 111932 497791
rect 111892 496868 111944 496874
rect 111892 496810 111944 496816
rect 111890 496496 111946 496505
rect 111890 496431 111946 496440
rect 111798 495816 111854 495825
rect 111798 495751 111800 495760
rect 111852 495751 111854 495760
rect 111800 495722 111852 495728
rect 111904 495514 111932 496431
rect 111996 496126 112024 499151
rect 111984 496120 112036 496126
rect 111984 496062 112036 496068
rect 111892 495508 111944 495514
rect 111892 495450 111944 495456
rect 111798 495136 111854 495145
rect 111798 495071 111800 495080
rect 111852 495071 111854 495080
rect 111800 495042 111852 495048
rect 111798 494456 111854 494465
rect 111798 494391 111854 494400
rect 111812 494086 111840 494391
rect 111800 494080 111852 494086
rect 111800 494022 111852 494028
rect 111798 493776 111854 493785
rect 111798 493711 111854 493720
rect 111812 492726 111840 493711
rect 111800 492720 111852 492726
rect 111800 492662 111852 492668
rect 111890 492416 111946 492425
rect 111890 492351 111946 492360
rect 111798 491736 111854 491745
rect 111798 491671 111854 491680
rect 111812 491434 111840 491671
rect 111800 491428 111852 491434
rect 111800 491370 111852 491376
rect 111904 491366 111932 492351
rect 111892 491360 111944 491366
rect 111892 491302 111944 491308
rect 111890 491056 111946 491065
rect 111890 490991 111946 491000
rect 111798 490376 111854 490385
rect 111798 490311 111854 490320
rect 111812 490006 111840 490311
rect 111800 490000 111852 490006
rect 111800 489942 111852 489948
rect 111904 489938 111932 490991
rect 111892 489932 111944 489938
rect 111892 489874 111944 489880
rect 111890 489696 111946 489705
rect 111890 489631 111946 489640
rect 111798 489016 111854 489025
rect 111798 488951 111854 488960
rect 111812 488578 111840 488951
rect 111904 488646 111932 489631
rect 111892 488640 111944 488646
rect 111892 488582 111944 488588
rect 111800 488572 111852 488578
rect 111800 488514 111852 488520
rect 111890 488336 111946 488345
rect 111890 488271 111946 488280
rect 111798 487656 111854 487665
rect 111798 487591 111854 487600
rect 111812 487286 111840 487591
rect 111800 487280 111852 487286
rect 111800 487222 111852 487228
rect 111904 487218 111932 488271
rect 111892 487212 111944 487218
rect 111892 487154 111944 487160
rect 111890 486976 111946 486985
rect 111890 486911 111946 486920
rect 111798 486296 111854 486305
rect 111798 486231 111854 486240
rect 111812 485858 111840 486231
rect 111904 485926 111932 486911
rect 111892 485920 111944 485926
rect 111892 485862 111944 485868
rect 111800 485852 111852 485858
rect 111800 485794 111852 485800
rect 111798 484936 111854 484945
rect 111798 484871 111854 484880
rect 111812 484430 111840 484871
rect 111800 484424 111852 484430
rect 111800 484366 111852 484372
rect 111890 484256 111946 484265
rect 111890 484191 111946 484200
rect 111798 483576 111854 483585
rect 111798 483511 111854 483520
rect 111812 483138 111840 483511
rect 111800 483132 111852 483138
rect 111800 483074 111852 483080
rect 111904 483070 111932 484191
rect 111892 483064 111944 483070
rect 111892 483006 111944 483012
rect 111890 482896 111946 482905
rect 111890 482831 111946 482840
rect 111798 482216 111854 482225
rect 111798 482151 111854 482160
rect 111812 481778 111840 482151
rect 111800 481772 111852 481778
rect 111800 481714 111852 481720
rect 111904 481710 111932 482831
rect 111892 481704 111944 481710
rect 111892 481646 111944 481652
rect 111890 481536 111946 481545
rect 111890 481471 111946 481480
rect 111798 480856 111854 480865
rect 111798 480791 111854 480800
rect 111812 480350 111840 480791
rect 111800 480344 111852 480350
rect 111800 480286 111852 480292
rect 111904 480282 111932 481471
rect 111892 480276 111944 480282
rect 111892 480218 111944 480224
rect 111890 480176 111946 480185
rect 111890 480111 111946 480120
rect 111798 479496 111854 479505
rect 111798 479431 111854 479440
rect 111812 478990 111840 479431
rect 111800 478984 111852 478990
rect 111800 478926 111852 478932
rect 111904 478922 111932 480111
rect 111892 478916 111944 478922
rect 111892 478858 111944 478864
rect 111890 478816 111946 478825
rect 111890 478751 111946 478760
rect 111798 478136 111854 478145
rect 111798 478071 111854 478080
rect 111812 477698 111840 478071
rect 111800 477692 111852 477698
rect 111800 477634 111852 477640
rect 111904 477562 111932 478751
rect 111892 477556 111944 477562
rect 111892 477498 111944 477504
rect 112364 476814 112392 505271
rect 112352 476808 112404 476814
rect 111798 476776 111854 476785
rect 112352 476750 112404 476756
rect 111798 476711 111854 476720
rect 111812 476134 111840 476711
rect 111800 476128 111852 476134
rect 111800 476070 111852 476076
rect 111890 476096 111946 476105
rect 111890 476031 111946 476040
rect 111798 475416 111854 475425
rect 111798 475351 111854 475360
rect 111812 474842 111840 475351
rect 111800 474836 111852 474842
rect 111800 474778 111852 474784
rect 111904 474774 111932 476031
rect 111892 474768 111944 474774
rect 111798 474736 111854 474745
rect 111892 474710 111944 474716
rect 111798 474671 111854 474680
rect 111812 474094 111840 474671
rect 111800 474088 111852 474094
rect 111800 474030 111852 474036
rect 111890 474056 111946 474065
rect 111890 473991 111946 474000
rect 111800 473476 111852 473482
rect 111800 473418 111852 473424
rect 111812 473385 111840 473418
rect 111904 473414 111932 473991
rect 111892 473408 111944 473414
rect 111798 473376 111854 473385
rect 111892 473350 111944 473356
rect 111798 473311 111854 473320
rect 111890 472696 111946 472705
rect 111890 472631 111946 472640
rect 111800 472116 111852 472122
rect 111800 472058 111852 472064
rect 111812 472025 111840 472058
rect 111904 472054 111932 472631
rect 111892 472048 111944 472054
rect 111798 472016 111854 472025
rect 111892 471990 111944 471996
rect 111798 471951 111854 471960
rect 111890 471336 111946 471345
rect 111890 471271 111946 471280
rect 111904 470694 111932 471271
rect 111892 470688 111944 470694
rect 111798 470656 111854 470665
rect 111892 470630 111944 470636
rect 111798 470591 111800 470600
rect 111852 470591 111854 470600
rect 111800 470562 111852 470568
rect 111798 469976 111854 469985
rect 111798 469911 111854 469920
rect 111812 469402 111840 469911
rect 111800 469396 111852 469402
rect 111800 469338 111852 469344
rect 111798 469296 111854 469305
rect 111798 469231 111800 469240
rect 111852 469231 111854 469240
rect 111800 469202 111852 469208
rect 111890 468616 111946 468625
rect 111890 468551 111946 468560
rect 111800 467968 111852 467974
rect 111798 467936 111800 467945
rect 111852 467936 111854 467945
rect 111904 467906 111932 468551
rect 111798 467871 111854 467880
rect 111892 467900 111944 467906
rect 111892 467842 111944 467848
rect 111890 467256 111946 467265
rect 111890 467191 111946 467200
rect 111798 466576 111854 466585
rect 111798 466511 111800 466520
rect 111852 466511 111854 466520
rect 111800 466482 111852 466488
rect 111904 466478 111932 467191
rect 111892 466472 111944 466478
rect 111892 466414 111944 466420
rect 111890 465896 111946 465905
rect 111890 465831 111946 465840
rect 111798 465216 111854 465225
rect 111904 465186 111932 465831
rect 111798 465151 111854 465160
rect 111892 465180 111944 465186
rect 111812 465118 111840 465151
rect 111892 465122 111944 465128
rect 111800 465112 111852 465118
rect 111800 465054 111852 465060
rect 111890 464536 111946 464545
rect 111890 464471 111946 464480
rect 111798 463856 111854 463865
rect 111798 463791 111800 463800
rect 111852 463791 111854 463800
rect 111800 463762 111852 463768
rect 111904 463758 111932 464471
rect 111892 463752 111944 463758
rect 111892 463694 111944 463700
rect 111890 463176 111946 463185
rect 111890 463111 111946 463120
rect 111798 462496 111854 462505
rect 111798 462431 111800 462440
rect 111852 462431 111854 462440
rect 111800 462402 111852 462408
rect 111904 462398 111932 463111
rect 111892 462392 111944 462398
rect 111892 462334 111944 462340
rect 111890 461816 111946 461825
rect 111890 461751 111946 461760
rect 111798 461136 111854 461145
rect 111798 461071 111854 461080
rect 111812 461038 111840 461071
rect 111800 461032 111852 461038
rect 111800 460974 111852 460980
rect 111904 460970 111932 461751
rect 111892 460964 111944 460970
rect 111892 460906 111944 460912
rect 111798 460456 111854 460465
rect 111798 460391 111854 460400
rect 111812 459610 111840 460391
rect 112350 459776 112406 459785
rect 112350 459711 112406 459720
rect 111800 459604 111852 459610
rect 111800 459546 111852 459552
rect 111890 459096 111946 459105
rect 111890 459031 111946 459040
rect 111798 458416 111854 458425
rect 111798 458351 111854 458360
rect 111812 458318 111840 458351
rect 111800 458312 111852 458318
rect 111800 458254 111852 458260
rect 111904 458250 111932 459031
rect 111892 458244 111944 458250
rect 111892 458186 111944 458192
rect 112258 457736 112314 457745
rect 112258 457671 112314 457680
rect 111798 457056 111854 457065
rect 111798 456991 111854 457000
rect 111812 456822 111840 456991
rect 111800 456816 111852 456822
rect 111800 456758 111852 456764
rect 111890 456376 111946 456385
rect 111890 456311 111946 456320
rect 111798 455696 111854 455705
rect 111798 455631 111854 455640
rect 111812 455462 111840 455631
rect 111904 455530 111932 456311
rect 111892 455524 111944 455530
rect 111892 455466 111944 455472
rect 111800 455456 111852 455462
rect 111800 455398 111852 455404
rect 111798 455016 111854 455025
rect 111798 454951 111854 454960
rect 111812 454578 111840 454951
rect 111800 454572 111852 454578
rect 111800 454514 111852 454520
rect 111798 454336 111854 454345
rect 111798 454271 111854 454280
rect 111812 454102 111840 454271
rect 111800 454096 111852 454102
rect 111800 454038 111852 454044
rect 111890 453656 111946 453665
rect 111890 453591 111946 453600
rect 111798 452976 111854 452985
rect 111798 452911 111854 452920
rect 111812 452742 111840 452911
rect 111800 452736 111852 452742
rect 111800 452678 111852 452684
rect 111904 452674 111932 453591
rect 111892 452668 111944 452674
rect 111892 452610 111944 452616
rect 111890 452296 111946 452305
rect 111890 452231 111946 452240
rect 111798 451616 111854 451625
rect 111798 451551 111854 451560
rect 111812 451314 111840 451551
rect 111904 451382 111932 452231
rect 111892 451376 111944 451382
rect 111892 451318 111944 451324
rect 111800 451308 111852 451314
rect 111800 451250 111852 451256
rect 111890 450936 111946 450945
rect 111890 450871 111946 450880
rect 111798 450256 111854 450265
rect 111798 450191 111854 450200
rect 111812 450022 111840 450191
rect 111800 450016 111852 450022
rect 111800 449958 111852 449964
rect 111904 449954 111932 450871
rect 111892 449948 111944 449954
rect 111892 449890 111944 449896
rect 111890 449576 111946 449585
rect 111890 449511 111946 449520
rect 111798 448896 111854 448905
rect 111798 448831 111854 448840
rect 111812 448662 111840 448831
rect 111800 448656 111852 448662
rect 111800 448598 111852 448604
rect 111904 448594 111932 449511
rect 111892 448588 111944 448594
rect 111892 448530 111944 448536
rect 111798 448216 111854 448225
rect 111798 448151 111854 448160
rect 111812 447166 111840 448151
rect 111800 447160 111852 447166
rect 111800 447102 111852 447108
rect 112272 354686 112300 457671
rect 112260 354680 112312 354686
rect 112260 354622 112312 354628
rect 112364 354618 112392 459711
rect 112456 396030 112484 529790
rect 112444 396024 112496 396030
rect 112444 395966 112496 395972
rect 112548 387530 112576 529910
rect 112732 529802 112760 533831
rect 112640 529774 112760 529802
rect 112536 387524 112588 387530
rect 112536 387466 112588 387472
rect 112640 385014 112668 529774
rect 112718 525056 112774 525065
rect 112718 524991 112774 525000
rect 112628 385008 112680 385014
rect 112628 384950 112680 384956
rect 112732 380866 112760 524991
rect 112824 519586 112852 547431
rect 112902 544776 112958 544785
rect 112902 544711 112958 544720
rect 112916 521218 112944 544711
rect 112904 521212 112956 521218
rect 112904 521154 112956 521160
rect 112812 519580 112864 519586
rect 112812 519522 112864 519528
rect 112810 518256 112866 518265
rect 112810 518191 112866 518200
rect 112720 380860 112772 380866
rect 112720 380802 112772 380808
rect 112824 378146 112852 518191
rect 112902 510096 112958 510105
rect 112902 510031 112958 510040
rect 112812 378140 112864 378146
rect 112812 378082 112864 378088
rect 112916 375358 112944 510031
rect 113008 508570 113036 563751
rect 113088 552696 113140 552702
rect 113088 552638 113140 552644
rect 113100 541686 113128 552638
rect 113088 541680 113140 541686
rect 113088 541622 113140 541628
rect 113086 541376 113142 541385
rect 113086 541311 113142 541320
rect 113100 534750 113128 541311
rect 113088 534744 113140 534750
rect 113088 534686 113140 534692
rect 113086 533216 113142 533225
rect 113086 533151 113142 533160
rect 113100 532778 113128 533151
rect 113088 532772 113140 532778
rect 113088 532714 113140 532720
rect 113086 531856 113142 531865
rect 113086 531791 113142 531800
rect 113100 531418 113128 531791
rect 113088 531412 113140 531418
rect 113088 531354 113140 531360
rect 113086 531176 113142 531185
rect 113086 531111 113142 531120
rect 113100 530058 113128 531111
rect 113088 530052 113140 530058
rect 113088 529994 113140 530000
rect 113086 529136 113142 529145
rect 113086 529071 113142 529080
rect 113100 526538 113128 529071
rect 113100 526510 113220 526538
rect 113086 526416 113142 526425
rect 113086 526351 113142 526360
rect 113100 525842 113128 526351
rect 113088 525836 113140 525842
rect 113088 525778 113140 525784
rect 113192 525722 113220 526510
rect 113100 525694 113220 525722
rect 113100 520946 113128 525694
rect 113180 521212 113232 521218
rect 113180 521154 113232 521160
rect 113088 520940 113140 520946
rect 113088 520882 113140 520888
rect 113192 520826 113220 521154
rect 113100 520798 113220 520826
rect 113100 515438 113128 520798
rect 113088 515432 113140 515438
rect 113088 515374 113140 515380
rect 112996 508564 113048 508570
rect 112996 508506 113048 508512
rect 113086 493096 113142 493105
rect 113086 493031 113142 493040
rect 112994 485616 113050 485625
rect 112994 485551 113050 485560
rect 112904 375352 112956 375358
rect 112904 375294 112956 375300
rect 113008 365430 113036 485551
rect 113100 485110 113128 493031
rect 113088 485104 113140 485110
rect 113088 485046 113140 485052
rect 113086 477456 113142 477465
rect 113086 477391 113142 477400
rect 112996 365424 113048 365430
rect 112996 365366 113048 365372
rect 113100 362914 113128 477391
rect 113836 405686 113864 585346
rect 113916 583908 113968 583914
rect 113916 583850 113968 583856
rect 113824 405680 113876 405686
rect 113824 405622 113876 405628
rect 113928 405618 113956 583850
rect 117964 583772 118016 583778
rect 117964 583714 118016 583720
rect 115204 582412 115256 582418
rect 115204 582354 115256 582360
rect 114008 574388 114060 574394
rect 114008 574330 114060 574336
rect 113916 405612 113968 405618
rect 113916 405554 113968 405560
rect 114020 401402 114048 574330
rect 114100 527264 114152 527270
rect 114100 527206 114152 527212
rect 114008 401396 114060 401402
rect 114008 401338 114060 401344
rect 114112 382226 114140 527206
rect 114192 514888 114244 514894
rect 114192 514830 114244 514836
rect 114100 382220 114152 382226
rect 114100 382162 114152 382168
rect 114204 376718 114232 514830
rect 114284 503940 114336 503946
rect 114284 503882 114336 503888
rect 114192 376712 114244 376718
rect 114192 376654 114244 376660
rect 114296 372570 114324 503882
rect 114376 495100 114428 495106
rect 114376 495042 114428 495048
rect 114284 372564 114336 372570
rect 114284 372506 114336 372512
rect 114388 369850 114416 495042
rect 114468 477692 114520 477698
rect 114468 477634 114520 477640
rect 114376 369844 114428 369850
rect 114376 369786 114428 369792
rect 113088 362908 113140 362914
rect 113088 362850 113140 362856
rect 114480 362846 114508 477634
rect 115112 469396 115164 469402
rect 115112 469338 115164 469344
rect 115020 454572 115072 454578
rect 115020 454514 115072 454520
rect 114468 362840 114520 362846
rect 114468 362782 114520 362788
rect 112352 354612 112404 354618
rect 112352 354554 112404 354560
rect 115032 353258 115060 454514
rect 115124 358562 115152 469338
rect 115216 404326 115244 582354
rect 116768 579760 116820 579766
rect 116768 579702 116820 579708
rect 116584 565956 116636 565962
rect 116584 565898 116636 565904
rect 115296 561740 115348 561746
rect 115296 561682 115348 561688
rect 115204 404320 115256 404326
rect 115204 404262 115256 404268
rect 115308 395962 115336 561682
rect 115388 559020 115440 559026
rect 115388 558962 115440 558968
rect 115296 395956 115348 395962
rect 115296 395898 115348 395904
rect 115400 394670 115428 558962
rect 115480 554940 115532 554946
rect 115480 554882 115532 554888
rect 115388 394664 115440 394670
rect 115388 394606 115440 394612
rect 115492 393038 115520 554882
rect 115572 548140 115624 548146
rect 115572 548082 115624 548088
rect 115480 393032 115532 393038
rect 115480 392974 115532 392980
rect 115584 390250 115612 548082
rect 115664 499724 115716 499730
rect 115664 499666 115716 499672
rect 115572 390244 115624 390250
rect 115572 390186 115624 390192
rect 115676 371210 115704 499666
rect 115756 495780 115808 495786
rect 115756 495722 115808 495728
rect 115664 371204 115716 371210
rect 115664 371146 115716 371152
rect 115768 369782 115796 495722
rect 115848 474088 115900 474094
rect 115848 474030 115900 474036
rect 115756 369776 115808 369782
rect 115756 369718 115808 369724
rect 115860 361554 115888 474030
rect 116400 452736 116452 452742
rect 116400 452678 116452 452684
rect 115848 361548 115900 361554
rect 115848 361490 115900 361496
rect 115112 358556 115164 358562
rect 115112 358498 115164 358504
rect 116412 354550 116440 452678
rect 116492 448656 116544 448662
rect 116492 448598 116544 448604
rect 116400 354544 116452 354550
rect 116400 354486 116452 354492
rect 115020 353252 115072 353258
rect 115020 353194 115072 353200
rect 116504 350538 116532 448598
rect 116596 397458 116624 565898
rect 116676 550724 116728 550730
rect 116676 550666 116728 550672
rect 116584 397452 116636 397458
rect 116584 397394 116636 397400
rect 116688 391678 116716 550666
rect 116780 543046 116808 579702
rect 116768 543040 116820 543046
rect 116768 542982 116820 542988
rect 116860 542496 116912 542502
rect 116860 542438 116912 542444
rect 116768 541000 116820 541006
rect 116768 540942 116820 540948
rect 116676 391672 116728 391678
rect 116676 391614 116728 391620
rect 116780 387734 116808 540942
rect 116872 389162 116900 542438
rect 116952 533792 117004 533798
rect 116952 533734 117004 533740
rect 116860 389156 116912 389162
rect 116860 389098 116912 389104
rect 116768 387728 116820 387734
rect 116768 387670 116820 387676
rect 116964 384946 116992 533734
rect 117044 525768 117096 525774
rect 117044 525710 117096 525716
rect 116952 384940 117004 384946
rect 116952 384882 117004 384888
rect 117056 382158 117084 525710
rect 117136 510740 117188 510746
rect 117136 510682 117188 510688
rect 117044 382152 117096 382158
rect 117044 382094 117096 382100
rect 117148 375290 117176 510682
rect 117228 467968 117280 467974
rect 117228 467910 117280 467916
rect 117136 375284 117188 375290
rect 117136 375226 117188 375232
rect 117240 358698 117268 467910
rect 117976 407794 118004 583714
rect 118056 558952 118108 558958
rect 118056 558894 118108 558900
rect 117964 407788 118016 407794
rect 117964 407730 118016 407736
rect 118068 394602 118096 558894
rect 119344 554056 119396 554062
rect 119344 553998 119396 554004
rect 118148 545216 118200 545222
rect 118148 545158 118200 545164
rect 118056 394596 118108 394602
rect 118056 394538 118108 394544
rect 118160 390454 118188 545158
rect 118240 521756 118292 521762
rect 118240 521698 118292 521704
rect 118148 390448 118200 390454
rect 118148 390390 118200 390396
rect 118252 380798 118280 521698
rect 118332 519648 118384 519654
rect 118332 519590 118384 519596
rect 118240 380792 118292 380798
rect 118240 380734 118292 380740
rect 118344 379234 118372 519590
rect 118424 487280 118476 487286
rect 118424 487222 118476 487228
rect 118332 379228 118384 379234
rect 118332 379170 118384 379176
rect 118436 374678 118464 487222
rect 118516 478984 118568 478990
rect 118516 478926 118568 478932
rect 118424 374672 118476 374678
rect 118424 374614 118476 374620
rect 118528 367810 118556 478926
rect 119252 450016 119304 450022
rect 119252 449958 119304 449964
rect 118516 367804 118568 367810
rect 118516 367746 118568 367752
rect 117228 358692 117280 358698
rect 117228 358634 117280 358640
rect 119264 355366 119292 449958
rect 119356 393242 119384 553998
rect 119436 549364 119488 549370
rect 119436 549306 119488 549312
rect 119344 393236 119396 393242
rect 119344 393178 119396 393184
rect 119448 390386 119476 549306
rect 119528 542428 119580 542434
rect 119528 542370 119580 542376
rect 119436 390380 119488 390386
rect 119436 390322 119488 390328
rect 119540 389842 119568 542370
rect 119632 450566 119660 590718
rect 123484 589416 123536 589422
rect 123484 589358 123536 589364
rect 120724 584452 120776 584458
rect 120724 584394 120776 584400
rect 119712 516248 119764 516254
rect 119712 516190 119764 516196
rect 119620 450560 119672 450566
rect 119620 450502 119672 450508
rect 119528 389836 119580 389842
rect 119528 389778 119580 389784
rect 119724 378078 119752 516190
rect 119804 496936 119856 496942
rect 119804 496878 119856 496884
rect 119712 378072 119764 378078
rect 119712 378014 119764 378020
rect 119816 369714 119844 496878
rect 119896 462460 119948 462466
rect 119896 462402 119948 462408
rect 119804 369708 119856 369714
rect 119804 369650 119856 369656
rect 119908 355842 119936 462402
rect 119988 449948 120040 449954
rect 119988 449890 120040 449896
rect 119896 355836 119948 355842
rect 119896 355778 119948 355784
rect 119252 355360 119304 355366
rect 119252 355302 119304 355308
rect 120000 351898 120028 449890
rect 120736 405550 120764 584394
rect 122104 581052 122156 581058
rect 122104 580994 122156 581000
rect 120816 520396 120868 520402
rect 120816 520338 120868 520344
rect 120724 405544 120776 405550
rect 120724 405486 120776 405492
rect 120828 379438 120856 520338
rect 120908 514820 120960 514826
rect 120908 514762 120960 514768
rect 120816 379432 120868 379438
rect 120816 379374 120868 379380
rect 120920 378010 120948 514762
rect 121000 509924 121052 509930
rect 121000 509866 121052 509872
rect 120908 378004 120960 378010
rect 120908 377946 120960 377952
rect 121012 376650 121040 509866
rect 121092 503736 121144 503742
rect 121092 503678 121144 503684
rect 121000 376644 121052 376650
rect 121000 376586 121052 376592
rect 121104 372502 121132 503678
rect 121184 495508 121236 495514
rect 121184 495450 121236 495456
rect 121092 372496 121144 372502
rect 121092 372438 121144 372444
rect 121196 369646 121224 495450
rect 122116 404258 122144 580994
rect 122196 580304 122248 580310
rect 122196 580246 122248 580252
rect 122104 404252 122156 404258
rect 122104 404194 122156 404200
rect 122208 404190 122236 580246
rect 122288 570036 122340 570042
rect 122288 569978 122340 569984
rect 122196 404184 122248 404190
rect 122196 404126 122248 404132
rect 122300 400926 122328 569978
rect 122380 563712 122432 563718
rect 122380 563654 122432 563660
rect 122392 402694 122420 563654
rect 122656 508564 122708 508570
rect 122656 508506 122708 508512
rect 122472 491428 122524 491434
rect 122472 491370 122524 491376
rect 122380 402688 122432 402694
rect 122380 402630 122432 402636
rect 122288 400920 122340 400926
rect 122288 400862 122340 400868
rect 121184 369640 121236 369646
rect 121184 369582 121236 369588
rect 122484 368286 122512 491370
rect 122564 472116 122616 472122
rect 122564 472058 122616 472064
rect 122472 368280 122524 368286
rect 122472 368222 122524 368228
rect 122576 360194 122604 472058
rect 122668 397390 122696 508506
rect 122748 452668 122800 452674
rect 122748 452610 122800 452616
rect 122656 397384 122708 397390
rect 122656 397326 122708 397332
rect 122760 362234 122788 452610
rect 123496 406978 123524 589358
rect 123576 587920 123628 587926
rect 123576 587862 123628 587868
rect 123588 407114 123616 587862
rect 123760 586560 123812 586566
rect 123760 586502 123812 586508
rect 123668 585812 123720 585818
rect 123668 585754 123720 585760
rect 123576 407108 123628 407114
rect 123576 407050 123628 407056
rect 123680 407046 123708 585754
rect 123772 409154 123800 586502
rect 134524 579692 134576 579698
rect 134524 579634 134576 579640
rect 130384 578332 130436 578338
rect 130384 578274 130436 578280
rect 127624 569968 127676 569974
rect 127624 569910 127676 569916
rect 126244 552152 126296 552158
rect 126244 552094 126296 552100
rect 123852 529236 123904 529242
rect 123852 529178 123904 529184
rect 123760 409148 123812 409154
rect 123760 409090 123812 409096
rect 123668 407040 123720 407046
rect 123668 406982 123720 406988
rect 123484 406972 123536 406978
rect 123484 406914 123536 406920
rect 123864 405482 123892 529178
rect 124864 528624 124916 528630
rect 124864 528566 124916 528572
rect 123944 483132 123996 483138
rect 123944 483074 123996 483080
rect 123852 405476 123904 405482
rect 123852 405418 123904 405424
rect 123956 364342 123984 483074
rect 124036 480344 124088 480350
rect 124036 480286 124088 480292
rect 124048 366382 124076 480286
rect 124128 451376 124180 451382
rect 124128 451318 124180 451324
rect 124036 366376 124088 366382
rect 124036 366318 124088 366324
rect 123944 364336 123996 364342
rect 123944 364278 123996 364284
rect 122748 362228 122800 362234
rect 122748 362170 122800 362176
rect 122564 360188 122616 360194
rect 122564 360130 122616 360136
rect 119988 351892 120040 351898
rect 119988 351834 120040 351840
rect 124140 351830 124168 451318
rect 124876 383382 124904 528566
rect 124956 520328 125008 520334
rect 124956 520270 125008 520276
rect 124864 383376 124916 383382
rect 124864 383318 124916 383324
rect 124968 379370 124996 520270
rect 125048 513460 125100 513466
rect 125048 513402 125100 513408
rect 124956 379364 125008 379370
rect 124956 379306 125008 379312
rect 125060 376582 125088 513402
rect 125232 476808 125284 476814
rect 125232 476750 125284 476756
rect 125140 465180 125192 465186
rect 125140 465122 125192 465128
rect 125048 376576 125100 376582
rect 125048 376518 125100 376524
rect 125152 357134 125180 465122
rect 125244 373998 125272 476750
rect 126256 391882 126284 552094
rect 126520 547936 126572 547942
rect 126520 547878 126572 547884
rect 126336 521688 126388 521694
rect 126336 521630 126388 521636
rect 126244 391876 126296 391882
rect 126244 391818 126296 391824
rect 126348 380730 126376 521630
rect 126428 505164 126480 505170
rect 126428 505106 126480 505112
rect 126336 380724 126388 380730
rect 126336 380666 126388 380672
rect 125232 373992 125284 373998
rect 125232 373934 125284 373940
rect 126440 373930 126468 505106
rect 126532 504422 126560 547878
rect 126612 507952 126664 507958
rect 126612 507894 126664 507900
rect 126520 504416 126572 504422
rect 126520 504358 126572 504364
rect 126624 497486 126652 507894
rect 126612 497480 126664 497486
rect 126612 497422 126664 497428
rect 126796 496868 126848 496874
rect 126796 496810 126848 496816
rect 126704 491360 126756 491366
rect 126704 491302 126756 491308
rect 126520 488640 126572 488646
rect 126520 488582 126572 488588
rect 126428 373924 126480 373930
rect 126428 373866 126480 373872
rect 126532 367062 126560 488582
rect 126716 480962 126744 491302
rect 126704 480956 126756 480962
rect 126704 480898 126756 480904
rect 126612 480276 126664 480282
rect 126612 480218 126664 480224
rect 126520 367056 126572 367062
rect 126520 366998 126572 367004
rect 126624 364274 126652 480218
rect 126704 472048 126756 472054
rect 126704 471990 126756 471996
rect 126612 364268 126664 364274
rect 126612 364210 126664 364216
rect 126716 360126 126744 471990
rect 126808 385694 126836 496810
rect 126888 463820 126940 463826
rect 126888 463762 126940 463768
rect 126796 385688 126848 385694
rect 126796 385630 126848 385636
rect 126704 360120 126756 360126
rect 126704 360062 126756 360068
rect 126900 357338 126928 463762
rect 127636 400178 127664 569910
rect 127716 564528 127768 564534
rect 127716 564470 127768 564476
rect 127624 400172 127676 400178
rect 127624 400114 127676 400120
rect 127728 398138 127756 564470
rect 127808 557660 127860 557666
rect 127808 557602 127860 557608
rect 127716 398132 127768 398138
rect 127716 398074 127768 398080
rect 127820 395350 127848 557602
rect 127900 538348 127952 538354
rect 127900 538290 127952 538296
rect 127808 395344 127860 395350
rect 127808 395286 127860 395292
rect 127912 386170 127940 538290
rect 129004 536920 129056 536926
rect 129004 536862 129056 536868
rect 127992 498228 128044 498234
rect 127992 498170 128044 498176
rect 127900 386164 127952 386170
rect 127900 386106 127952 386112
rect 128004 371142 128032 498170
rect 128084 490000 128136 490006
rect 128084 489942 128136 489948
rect 127992 371136 128044 371142
rect 127992 371078 128044 371084
rect 128096 366994 128124 489942
rect 128176 481772 128228 481778
rect 128176 481714 128228 481720
rect 128084 366988 128136 366994
rect 128084 366930 128136 366936
rect 128188 364206 128216 481714
rect 128268 473476 128320 473482
rect 128268 473418 128320 473424
rect 128176 364200 128228 364206
rect 128176 364142 128228 364148
rect 128280 360058 128308 473418
rect 129016 393990 129044 536862
rect 129096 506524 129148 506530
rect 129096 506466 129148 506472
rect 129004 393984 129056 393990
rect 129004 393926 129056 393932
rect 129108 373862 129136 506466
rect 129188 489932 129240 489938
rect 129188 489874 129240 489880
rect 129096 373856 129148 373862
rect 129096 373798 129148 373804
rect 129200 368422 129228 489874
rect 129280 481704 129332 481710
rect 129280 481646 129332 481652
rect 129188 368416 129240 368422
rect 129188 368358 129240 368364
rect 129292 364138 129320 481646
rect 129372 473408 129424 473414
rect 129372 473350 129424 473356
rect 129280 364132 129332 364138
rect 129280 364074 129332 364080
rect 129384 361486 129412 473350
rect 130396 402898 130424 578274
rect 133144 578264 133196 578270
rect 133144 578206 133196 578212
rect 132040 575612 132092 575618
rect 132040 575554 132092 575560
rect 130476 571464 130528 571470
rect 130476 571406 130528 571412
rect 130384 402892 130436 402898
rect 130384 402834 130436 402840
rect 130488 400110 130516 571406
rect 130568 564460 130620 564466
rect 130568 564402 130620 564408
rect 130476 400104 130528 400110
rect 130476 400046 130528 400052
rect 130580 397322 130608 564402
rect 130660 557592 130712 557598
rect 130660 557534 130712 557540
rect 130568 397316 130620 397322
rect 130568 397258 130620 397264
rect 130672 394534 130700 557534
rect 130752 550656 130804 550662
rect 130752 550598 130804 550604
rect 130660 394528 130712 394534
rect 130660 394470 130712 394476
rect 130764 391814 130792 550598
rect 131764 545148 131816 545154
rect 131764 545090 131816 545096
rect 130844 515432 130896 515438
rect 130844 515374 130896 515380
rect 130752 391808 130804 391814
rect 130752 391750 130804 391756
rect 130856 389094 130884 515374
rect 130936 458312 130988 458318
rect 130936 458254 130988 458260
rect 130844 389088 130896 389094
rect 130844 389030 130896 389036
rect 129372 361480 129424 361486
rect 129372 361422 129424 361428
rect 128268 360052 128320 360058
rect 128268 359994 128320 360000
rect 126888 357332 126940 357338
rect 126888 357274 126940 357280
rect 125140 357128 125192 357134
rect 125140 357070 125192 357076
rect 130948 355434 130976 458254
rect 131776 389026 131804 545090
rect 131856 536852 131908 536858
rect 131856 536794 131908 536800
rect 131764 389020 131816 389026
rect 131764 388962 131816 388968
rect 131868 386306 131896 536794
rect 131948 530052 132000 530058
rect 131948 529994 132000 530000
rect 131856 386300 131908 386306
rect 131856 386242 131908 386248
rect 131960 383586 131988 529994
rect 132052 529242 132080 575554
rect 132040 529236 132092 529242
rect 132040 529178 132092 529184
rect 132040 523116 132092 523122
rect 132040 523058 132092 523064
rect 131948 383580 132000 383586
rect 131948 383522 132000 383528
rect 132052 380662 132080 523058
rect 132132 474836 132184 474842
rect 132132 474778 132184 474784
rect 132040 380656 132092 380662
rect 132040 380598 132092 380604
rect 132144 361418 132172 474778
rect 132224 466540 132276 466546
rect 132224 466482 132276 466488
rect 132132 361412 132184 361418
rect 132132 361354 132184 361360
rect 132236 357270 132264 466482
rect 132316 456816 132368 456822
rect 132316 456758 132368 456764
rect 132224 357264 132276 357270
rect 132224 357206 132276 357212
rect 130936 355428 130988 355434
rect 130936 355370 130988 355376
rect 132328 353122 132356 456758
rect 132408 455524 132460 455530
rect 132408 455466 132460 455472
rect 132420 353190 132448 455466
rect 133156 402830 133184 578206
rect 133236 571396 133288 571402
rect 133236 571338 133288 571344
rect 133144 402824 133196 402830
rect 133144 402766 133196 402772
rect 133248 400042 133276 571338
rect 133328 499588 133380 499594
rect 133328 499530 133380 499536
rect 133236 400036 133288 400042
rect 133236 399978 133288 399984
rect 133340 371074 133368 499530
rect 133420 483064 133472 483070
rect 133420 483006 133472 483012
rect 133328 371068 133380 371074
rect 133328 371010 133380 371016
rect 133432 365634 133460 483006
rect 133512 474768 133564 474774
rect 133512 474710 133564 474716
rect 133420 365628 133472 365634
rect 133420 365570 133472 365576
rect 133524 361350 133552 474710
rect 133604 458244 133656 458250
rect 133604 458186 133656 458192
rect 133512 361344 133564 361350
rect 133512 361286 133564 361292
rect 133616 354482 133644 458186
rect 134536 402762 134564 579634
rect 134616 572824 134668 572830
rect 134616 572766 134668 572772
rect 134524 402756 134576 402762
rect 134524 402698 134576 402704
rect 134628 399974 134656 572766
rect 134708 565888 134760 565894
rect 134708 565830 134760 565836
rect 134616 399968 134668 399974
rect 134616 399910 134668 399916
rect 134524 397520 134576 397526
rect 134524 397462 134576 397468
rect 133604 354476 133656 354482
rect 133604 354418 133656 354424
rect 132408 353184 132460 353190
rect 132408 353126 132460 353132
rect 132316 353116 132368 353122
rect 132316 353058 132368 353064
rect 124128 351824 124180 351830
rect 124128 351766 124180 351772
rect 116492 350532 116544 350538
rect 116492 350474 116544 350480
rect 126244 349172 126296 349178
rect 126244 349114 126296 349120
rect 122656 348016 122708 348022
rect 122656 347958 122708 347964
rect 119436 347948 119488 347954
rect 119436 347890 119488 347896
rect 116676 347812 116728 347818
rect 116676 347754 116728 347760
rect 116584 346520 116636 346526
rect 116584 346462 116636 346468
rect 113916 346452 113968 346458
rect 113916 346394 113968 346400
rect 113824 345160 113876 345166
rect 113824 345102 113876 345108
rect 112260 337068 112312 337074
rect 112260 337010 112312 337016
rect 30012 318844 30064 318850
rect 30012 318786 30064 318792
rect 29920 133816 29972 133822
rect 29920 133758 29972 133764
rect 30024 133482 30052 318786
rect 111800 314628 111852 314634
rect 111800 314570 111852 314576
rect 111812 314265 111840 314570
rect 111798 314256 111854 314265
rect 111798 314191 111854 314200
rect 111800 313268 111852 313274
rect 111800 313210 111852 313216
rect 111812 313177 111840 313210
rect 111892 313200 111944 313206
rect 111798 313168 111854 313177
rect 111892 313142 111944 313148
rect 111798 313103 111854 313112
rect 111904 312769 111932 313142
rect 111890 312760 111946 312769
rect 111890 312695 111946 312704
rect 111892 311840 111944 311846
rect 111798 311808 111854 311817
rect 111892 311782 111944 311788
rect 111798 311743 111800 311752
rect 111852 311743 111854 311752
rect 111800 311714 111852 311720
rect 111904 311409 111932 311782
rect 111890 311400 111946 311409
rect 111890 311335 111946 311344
rect 111800 310480 111852 310486
rect 111798 310448 111800 310457
rect 111852 310448 111854 310457
rect 111798 310383 111854 310392
rect 111892 310412 111944 310418
rect 111892 310354 111944 310360
rect 111904 310049 111932 310354
rect 111890 310040 111946 310049
rect 111890 309975 111946 309984
rect 111800 309120 111852 309126
rect 111798 309088 111800 309097
rect 111852 309088 111854 309097
rect 111798 309023 111854 309032
rect 111892 309052 111944 309058
rect 111892 308994 111944 309000
rect 111904 308689 111932 308994
rect 111890 308680 111946 308689
rect 111890 308615 111946 308624
rect 111800 307760 111852 307766
rect 111798 307728 111800 307737
rect 111852 307728 111854 307737
rect 111798 307663 111854 307672
rect 111800 307556 111852 307562
rect 111800 307498 111852 307504
rect 111812 307329 111840 307498
rect 111798 307320 111854 307329
rect 111798 307255 111854 307264
rect 112076 306400 112128 306406
rect 111798 306368 111854 306377
rect 112076 306342 112128 306348
rect 111798 306303 111800 306312
rect 111852 306303 111854 306312
rect 111800 306274 111852 306280
rect 111892 306264 111944 306270
rect 111892 306206 111944 306212
rect 111904 305969 111932 306206
rect 111890 305960 111946 305969
rect 111890 305895 111946 305904
rect 30104 305040 30156 305046
rect 30104 304982 30156 304988
rect 30116 133890 30144 304982
rect 111892 304972 111944 304978
rect 111892 304914 111944 304920
rect 111800 304904 111852 304910
rect 111798 304872 111800 304881
rect 111852 304872 111854 304881
rect 111798 304807 111854 304816
rect 111904 304609 111932 304914
rect 111890 304600 111946 304609
rect 111890 304535 111946 304544
rect 112088 304502 112116 306342
rect 112076 304496 112128 304502
rect 112076 304438 112128 304444
rect 111892 303612 111944 303618
rect 111892 303554 111944 303560
rect 111800 303544 111852 303550
rect 111798 303512 111800 303521
rect 111852 303512 111854 303521
rect 111798 303447 111854 303456
rect 111904 303249 111932 303554
rect 111890 303240 111946 303249
rect 111890 303175 111946 303184
rect 111800 302184 111852 302190
rect 111798 302152 111800 302161
rect 111852 302152 111854 302161
rect 111798 302087 111854 302096
rect 111892 302116 111944 302122
rect 111892 302058 111944 302064
rect 111904 301889 111932 302058
rect 111890 301880 111946 301889
rect 111890 301815 111946 301824
rect 111984 300824 112036 300830
rect 111890 300792 111946 300801
rect 111984 300766 112036 300772
rect 111890 300727 111892 300736
rect 111944 300727 111946 300736
rect 111892 300698 111944 300704
rect 111800 300688 111852 300694
rect 111800 300630 111852 300636
rect 111812 300393 111840 300630
rect 111798 300384 111854 300393
rect 111798 300319 111854 300328
rect 111996 299985 112024 300766
rect 111982 299976 112038 299985
rect 111982 299911 112038 299920
rect 111800 299192 111852 299198
rect 111800 299134 111852 299140
rect 111812 299033 111840 299134
rect 111798 299024 111854 299033
rect 111798 298959 111854 298968
rect 111800 298852 111852 298858
rect 111800 298794 111852 298800
rect 111812 298489 111840 298794
rect 111798 298480 111854 298489
rect 111798 298415 111854 298424
rect 111892 298104 111944 298110
rect 111892 298046 111944 298052
rect 111800 297968 111852 297974
rect 111800 297910 111852 297916
rect 111812 297673 111840 297910
rect 111798 297664 111854 297673
rect 111798 297599 111854 297608
rect 111904 297265 111932 298046
rect 111890 297256 111946 297265
rect 111890 297191 111946 297200
rect 112272 296714 112300 337010
rect 112352 328500 112404 328506
rect 112352 328442 112404 328448
rect 112088 296686 112300 296714
rect 111800 296676 111852 296682
rect 111800 296618 111852 296624
rect 111812 296449 111840 296618
rect 111892 296608 111944 296614
rect 111892 296550 111944 296556
rect 111798 296440 111854 296449
rect 111798 296375 111854 296384
rect 111904 295905 111932 296550
rect 111890 295896 111946 295905
rect 111890 295831 111946 295840
rect 111892 295316 111944 295322
rect 111892 295258 111944 295264
rect 111800 295248 111852 295254
rect 111800 295190 111852 295196
rect 111812 294953 111840 295190
rect 111798 294944 111854 294953
rect 111798 294879 111854 294888
rect 111904 294545 111932 295258
rect 111890 294536 111946 294545
rect 111890 294471 111946 294480
rect 111800 293956 111852 293962
rect 111800 293898 111852 293904
rect 111812 293729 111840 293898
rect 111892 293888 111944 293894
rect 111892 293830 111944 293836
rect 111798 293720 111854 293729
rect 111798 293655 111854 293664
rect 111904 293185 111932 293830
rect 111890 293176 111946 293185
rect 111890 293111 111946 293120
rect 111892 292528 111944 292534
rect 111892 292470 111944 292476
rect 111800 292460 111852 292466
rect 111800 292402 111852 292408
rect 111812 292233 111840 292402
rect 111798 292224 111854 292233
rect 111798 292159 111854 292168
rect 111904 291825 111932 292470
rect 111890 291816 111946 291825
rect 111890 291751 111946 291760
rect 111892 291168 111944 291174
rect 111892 291110 111944 291116
rect 111800 291100 111852 291106
rect 111800 291042 111852 291048
rect 111812 290873 111840 291042
rect 111798 290864 111854 290873
rect 111798 290799 111854 290808
rect 111904 290465 111932 291110
rect 111890 290456 111946 290465
rect 111890 290391 111946 290400
rect 111800 289808 111852 289814
rect 111800 289750 111852 289756
rect 111812 289513 111840 289750
rect 111892 289740 111944 289746
rect 111892 289682 111944 289688
rect 111798 289504 111854 289513
rect 111798 289439 111854 289448
rect 111904 289105 111932 289682
rect 111890 289096 111946 289105
rect 111890 289031 111946 289040
rect 111892 288380 111944 288386
rect 111892 288322 111944 288328
rect 111800 288312 111852 288318
rect 111800 288254 111852 288260
rect 111812 288153 111840 288254
rect 111798 288144 111854 288153
rect 111798 288079 111854 288088
rect 111904 287745 111932 288322
rect 111890 287736 111946 287745
rect 111890 287671 111946 287680
rect 111892 287020 111944 287026
rect 111892 286962 111944 286968
rect 111800 286952 111852 286958
rect 111800 286894 111852 286900
rect 111812 286793 111840 286894
rect 111798 286784 111854 286793
rect 111798 286719 111854 286728
rect 111904 286385 111932 286962
rect 111890 286376 111946 286385
rect 111890 286311 111946 286320
rect 111800 285660 111852 285666
rect 111800 285602 111852 285608
rect 111812 285433 111840 285602
rect 111892 285592 111944 285598
rect 111892 285534 111944 285540
rect 111798 285424 111854 285433
rect 111798 285359 111854 285368
rect 111904 285025 111932 285534
rect 111890 285016 111946 285025
rect 111890 284951 111946 284960
rect 111892 284300 111944 284306
rect 111892 284242 111944 284248
rect 111800 284232 111852 284238
rect 111800 284174 111852 284180
rect 111812 284073 111840 284174
rect 111798 284064 111854 284073
rect 111798 283999 111854 284008
rect 111904 283665 111932 284242
rect 111890 283656 111946 283665
rect 111890 283591 111946 283600
rect 111800 282872 111852 282878
rect 112088 282849 112116 296686
rect 111800 282814 111852 282820
rect 112074 282840 112130 282849
rect 111812 282305 111840 282814
rect 112074 282775 112130 282784
rect 111798 282296 111854 282305
rect 111798 282231 111854 282240
rect 111892 281512 111944 281518
rect 111892 281454 111944 281460
rect 111800 281444 111852 281450
rect 111800 281386 111852 281392
rect 111812 281353 111840 281386
rect 111798 281344 111854 281353
rect 111798 281279 111854 281288
rect 111904 280945 111932 281454
rect 111890 280936 111946 280945
rect 111890 280871 111946 280880
rect 111800 280152 111852 280158
rect 111800 280094 111852 280100
rect 111812 279993 111840 280094
rect 111892 280084 111944 280090
rect 111892 280026 111944 280032
rect 111798 279984 111854 279993
rect 111798 279919 111854 279928
rect 111904 279585 111932 280026
rect 111890 279576 111946 279585
rect 111890 279511 111946 279520
rect 111892 278724 111944 278730
rect 111892 278666 111944 278672
rect 111800 278656 111852 278662
rect 111800 278598 111852 278604
rect 111812 278497 111840 278598
rect 111798 278488 111854 278497
rect 111798 278423 111854 278432
rect 111904 278225 111932 278666
rect 111890 278216 111946 278225
rect 111890 278151 111946 278160
rect 112364 277394 112392 328442
rect 113088 325984 113140 325990
rect 113088 325926 113140 325932
rect 112996 325780 113048 325786
rect 112996 325722 113048 325728
rect 112904 324624 112956 324630
rect 112904 324566 112956 324572
rect 112812 323264 112864 323270
rect 112812 323206 112864 323212
rect 112720 320204 112772 320210
rect 112720 320146 112772 320152
rect 112628 313336 112680 313342
rect 112628 313278 112680 313284
rect 112536 304496 112588 304502
rect 112536 304438 112588 304444
rect 112444 294024 112496 294030
rect 112444 293966 112496 293972
rect 111800 277364 111852 277370
rect 111800 277306 111852 277312
rect 112180 277366 112392 277394
rect 111812 277273 111840 277306
rect 111892 277296 111944 277302
rect 111798 277264 111854 277273
rect 111892 277238 111944 277244
rect 111798 277199 111854 277208
rect 111904 276865 111932 277238
rect 111890 276856 111946 276865
rect 111890 276791 111946 276800
rect 111800 276004 111852 276010
rect 111800 275946 111852 275952
rect 111812 275913 111840 275946
rect 111892 275936 111944 275942
rect 111798 275904 111854 275913
rect 111892 275878 111944 275884
rect 111798 275839 111854 275848
rect 111904 275505 111932 275878
rect 111890 275496 111946 275505
rect 111890 275431 111946 275440
rect 111892 274644 111944 274650
rect 111892 274586 111944 274592
rect 111800 274576 111852 274582
rect 111800 274518 111852 274524
rect 111812 274417 111840 274518
rect 111798 274408 111854 274417
rect 111798 274343 111854 274352
rect 111904 274145 111932 274586
rect 111890 274136 111946 274145
rect 111890 274071 111946 274080
rect 111892 273216 111944 273222
rect 111892 273158 111944 273164
rect 111800 273080 111852 273086
rect 111798 273048 111800 273057
rect 111852 273048 111854 273057
rect 111798 272983 111854 272992
rect 111904 272785 111932 273158
rect 111890 272776 111946 272785
rect 111890 272711 111946 272720
rect 111892 271856 111944 271862
rect 111892 271798 111944 271804
rect 111800 271788 111852 271794
rect 111800 271730 111852 271736
rect 111812 271697 111840 271730
rect 111798 271688 111854 271697
rect 111798 271623 111854 271632
rect 111904 271425 111932 271798
rect 111890 271416 111946 271425
rect 111890 271351 111946 271360
rect 111800 270496 111852 270502
rect 111800 270438 111852 270444
rect 111812 270337 111840 270438
rect 111892 270428 111944 270434
rect 111892 270370 111944 270376
rect 111798 270328 111854 270337
rect 111798 270263 111854 270272
rect 111904 270065 111932 270370
rect 111890 270056 111946 270065
rect 111890 269991 111946 270000
rect 111892 269068 111944 269074
rect 111892 269010 111944 269016
rect 111800 269000 111852 269006
rect 111798 268968 111800 268977
rect 111852 268968 111854 268977
rect 111798 268903 111854 268912
rect 111904 268705 111932 269010
rect 111890 268696 111946 268705
rect 111890 268631 111946 268640
rect 111800 267708 111852 267714
rect 111800 267650 111852 267656
rect 111812 267617 111840 267650
rect 111892 267640 111944 267646
rect 111798 267608 111854 267617
rect 111892 267582 111944 267588
rect 111798 267543 111854 267552
rect 111904 267209 111932 267582
rect 111890 267200 111946 267209
rect 111890 267135 111946 267144
rect 30196 266416 30248 266422
rect 30196 266358 30248 266364
rect 30104 133884 30156 133890
rect 30104 133826 30156 133832
rect 30208 133618 30236 266358
rect 111892 266348 111944 266354
rect 111892 266290 111944 266296
rect 111800 266280 111852 266286
rect 111798 266248 111800 266257
rect 111852 266248 111854 266257
rect 111798 266183 111854 266192
rect 111904 265985 111932 266290
rect 111890 265976 111946 265985
rect 111890 265911 111946 265920
rect 111892 264920 111944 264926
rect 111798 264888 111854 264897
rect 111892 264862 111944 264868
rect 111798 264823 111800 264832
rect 111852 264823 111854 264832
rect 111800 264794 111852 264800
rect 111904 264489 111932 264862
rect 111890 264480 111946 264489
rect 111890 264415 111946 264424
rect 111892 263560 111944 263566
rect 111798 263528 111854 263537
rect 111892 263502 111944 263508
rect 111798 263463 111800 263472
rect 111852 263463 111854 263472
rect 111800 263434 111852 263440
rect 111904 263129 111932 263502
rect 111890 263120 111946 263129
rect 111890 263055 111946 263064
rect 111800 262200 111852 262206
rect 112180 262177 112208 277366
rect 111800 262142 111852 262148
rect 112166 262168 112222 262177
rect 111812 261769 111840 262142
rect 112166 262103 112222 262112
rect 111798 261760 111854 261769
rect 111798 261695 111854 261704
rect 111800 260840 111852 260846
rect 111798 260808 111800 260817
rect 111852 260808 111854 260817
rect 111798 260743 111854 260752
rect 111892 260772 111944 260778
rect 111892 260714 111944 260720
rect 111904 260409 111932 260714
rect 112260 260704 112312 260710
rect 112260 260646 112312 260652
rect 111890 260400 111946 260409
rect 111890 260335 111946 260344
rect 111892 259412 111944 259418
rect 111892 259354 111944 259360
rect 111800 259344 111852 259350
rect 111798 259312 111800 259321
rect 111852 259312 111854 259321
rect 111798 259247 111854 259256
rect 111904 259049 111932 259354
rect 111890 259040 111946 259049
rect 111890 258975 111946 258984
rect 111892 258052 111944 258058
rect 111892 257994 111944 258000
rect 111800 257984 111852 257990
rect 111798 257952 111800 257961
rect 111852 257952 111854 257961
rect 111798 257887 111854 257896
rect 111904 257689 111932 257994
rect 111890 257680 111946 257689
rect 111890 257615 111946 257624
rect 111800 256692 111852 256698
rect 111800 256634 111852 256640
rect 111812 256329 111840 256634
rect 111798 256320 111854 256329
rect 111798 256255 111854 256264
rect 111800 255264 111852 255270
rect 111800 255206 111852 255212
rect 111812 254969 111840 255206
rect 111798 254960 111854 254969
rect 111798 254895 111854 254904
rect 111800 253904 111852 253910
rect 111798 253872 111800 253881
rect 111852 253872 111854 253881
rect 111798 253807 111854 253816
rect 111892 253836 111944 253842
rect 111892 253778 111944 253784
rect 111800 253768 111852 253774
rect 111800 253710 111852 253716
rect 111812 253065 111840 253710
rect 111904 253609 111932 253778
rect 111890 253600 111946 253609
rect 111890 253535 111946 253544
rect 111798 253056 111854 253065
rect 111798 252991 111854 253000
rect 111800 252544 111852 252550
rect 111800 252486 111852 252492
rect 111812 252249 111840 252486
rect 111798 252240 111854 252249
rect 111798 252175 111854 252184
rect 112272 251705 112300 260646
rect 112352 253020 112404 253026
rect 112352 252962 112404 252968
rect 112258 251696 112314 251705
rect 112258 251631 112314 251640
rect 111800 251184 111852 251190
rect 111800 251126 111852 251132
rect 111812 250889 111840 251126
rect 111892 251116 111944 251122
rect 111892 251058 111944 251064
rect 111798 250880 111854 250889
rect 111798 250815 111854 250824
rect 111904 250345 111932 251058
rect 111890 250336 111946 250345
rect 111890 250271 111946 250280
rect 111800 249756 111852 249762
rect 111800 249698 111852 249704
rect 111812 249529 111840 249698
rect 111798 249520 111854 249529
rect 111798 249455 111854 249464
rect 111892 248396 111944 248402
rect 111892 248338 111944 248344
rect 111800 248328 111852 248334
rect 111800 248270 111852 248276
rect 111812 248033 111840 248270
rect 111798 248024 111854 248033
rect 111798 247959 111854 247968
rect 111904 247625 111932 248338
rect 111890 247616 111946 247625
rect 111890 247551 111946 247560
rect 111892 247036 111944 247042
rect 111892 246978 111944 246984
rect 111800 246968 111852 246974
rect 111800 246910 111852 246916
rect 111812 246673 111840 246910
rect 111798 246664 111854 246673
rect 111798 246599 111854 246608
rect 111904 246265 111932 246978
rect 111890 246256 111946 246265
rect 111890 246191 111946 246200
rect 111800 245608 111852 245614
rect 111800 245550 111852 245556
rect 111812 245313 111840 245550
rect 111892 245540 111944 245546
rect 111892 245482 111944 245488
rect 111798 245304 111854 245313
rect 111798 245239 111854 245248
rect 111904 244905 111932 245482
rect 111890 244896 111946 244905
rect 111890 244831 111946 244840
rect 111800 244248 111852 244254
rect 111800 244190 111852 244196
rect 111812 243953 111840 244190
rect 111798 243944 111854 243953
rect 111798 243879 111854 243888
rect 111984 243568 112036 243574
rect 112364 243545 112392 252962
rect 111984 243510 112036 243516
rect 112350 243536 112406 243545
rect 111800 242888 111852 242894
rect 111800 242830 111852 242836
rect 111812 242593 111840 242830
rect 111798 242584 111854 242593
rect 111798 242519 111854 242528
rect 111892 242208 111944 242214
rect 111996 242185 112024 243510
rect 112350 243471 112406 243480
rect 111892 242150 111944 242156
rect 111982 242176 112038 242185
rect 111904 241505 111932 242150
rect 111982 242111 112038 242120
rect 111890 241496 111946 241505
rect 111800 241460 111852 241466
rect 111890 241431 111946 241440
rect 111800 241402 111852 241408
rect 111812 240825 111840 241402
rect 111798 240816 111854 240825
rect 111798 240751 111854 240760
rect 112352 240780 112404 240786
rect 112352 240722 112404 240728
rect 111800 240100 111852 240106
rect 111800 240042 111852 240048
rect 111812 239873 111840 240042
rect 111892 240032 111944 240038
rect 111892 239974 111944 239980
rect 111798 239864 111854 239873
rect 111798 239799 111854 239808
rect 111904 239465 111932 239974
rect 111890 239456 111946 239465
rect 111890 239391 111946 239400
rect 111800 238740 111852 238746
rect 111800 238682 111852 238688
rect 111812 238513 111840 238682
rect 111892 238536 111944 238542
rect 111798 238504 111854 238513
rect 111892 238478 111944 238484
rect 111798 238439 111854 238448
rect 111904 238105 111932 238478
rect 111890 238096 111946 238105
rect 111890 238031 111946 238040
rect 111800 237380 111852 237386
rect 111800 237322 111852 237328
rect 111812 237153 111840 237322
rect 111798 237144 111854 237153
rect 111798 237079 111854 237088
rect 112364 236745 112392 240722
rect 112350 236736 112406 236745
rect 111892 236700 111944 236706
rect 112350 236671 112406 236680
rect 111892 236642 111944 236648
rect 111800 235952 111852 235958
rect 111800 235894 111852 235900
rect 111812 235793 111840 235894
rect 111798 235784 111854 235793
rect 111798 235719 111854 235728
rect 111904 235385 111932 236642
rect 111890 235376 111946 235385
rect 111890 235311 111946 235320
rect 111892 235272 111944 235278
rect 111892 235214 111944 235220
rect 111800 234592 111852 234598
rect 111800 234534 111852 234540
rect 111812 234433 111840 234534
rect 111798 234424 111854 234433
rect 111798 234359 111854 234368
rect 111904 234025 111932 235214
rect 111890 234016 111946 234025
rect 111890 233951 111946 233960
rect 112352 233980 112404 233986
rect 112352 233922 112404 233928
rect 111800 233912 111852 233918
rect 111800 233854 111852 233860
rect 111812 233209 111840 233854
rect 111798 233200 111854 233209
rect 111798 233135 111854 233144
rect 111800 232960 111852 232966
rect 111800 232902 111852 232908
rect 111812 232529 111840 232902
rect 111798 232520 111854 232529
rect 111798 232455 111854 232464
rect 111800 231804 111852 231810
rect 111800 231746 111852 231752
rect 111812 231305 111840 231746
rect 111798 231296 111854 231305
rect 111798 231231 111854 231240
rect 111800 230444 111852 230450
rect 111800 230386 111852 230392
rect 111812 230353 111840 230386
rect 111892 230376 111944 230382
rect 111798 230344 111854 230353
rect 111892 230318 111944 230324
rect 111798 230279 111854 230288
rect 111904 229945 111932 230318
rect 111890 229936 111946 229945
rect 111890 229871 111946 229880
rect 111800 229084 111852 229090
rect 111800 229026 111852 229032
rect 111812 228993 111840 229026
rect 111892 229016 111944 229022
rect 111798 228984 111854 228993
rect 111892 228958 111944 228964
rect 111798 228919 111854 228928
rect 111904 228585 111932 228958
rect 111890 228576 111946 228585
rect 111890 228511 111946 228520
rect 111800 227724 111852 227730
rect 111800 227666 111852 227672
rect 111812 227633 111840 227666
rect 111892 227656 111944 227662
rect 111798 227624 111854 227633
rect 111892 227598 111944 227604
rect 111798 227559 111854 227568
rect 111904 227225 111932 227598
rect 111890 227216 111946 227225
rect 111890 227151 111946 227160
rect 112364 226273 112392 233922
rect 112350 226264 112406 226273
rect 112350 226199 112406 226208
rect 111800 226024 111852 226030
rect 111800 225966 111852 225972
rect 111812 225729 111840 225966
rect 111798 225720 111854 225729
rect 111798 225655 111854 225664
rect 111800 224936 111852 224942
rect 111800 224878 111852 224884
rect 111812 224777 111840 224878
rect 111892 224868 111944 224874
rect 111892 224810 111944 224816
rect 111798 224768 111854 224777
rect 111798 224703 111854 224712
rect 111904 224505 111932 224810
rect 111890 224496 111946 224505
rect 111890 224431 111946 224440
rect 111800 223576 111852 223582
rect 111800 223518 111852 223524
rect 111812 223417 111840 223518
rect 111892 223508 111944 223514
rect 111892 223450 111944 223456
rect 111798 223408 111854 223417
rect 111798 223343 111854 223352
rect 111904 223145 111932 223450
rect 111890 223136 111946 223145
rect 111890 223071 111946 223080
rect 111800 222148 111852 222154
rect 111800 222090 111852 222096
rect 111812 222057 111840 222090
rect 111892 222080 111944 222086
rect 111798 222048 111854 222057
rect 111892 222022 111944 222028
rect 111798 221983 111854 221992
rect 111904 221649 111932 222022
rect 111890 221640 111946 221649
rect 111890 221575 111946 221584
rect 111800 220788 111852 220794
rect 111800 220730 111852 220736
rect 111812 220697 111840 220730
rect 111892 220720 111944 220726
rect 111798 220688 111854 220697
rect 111892 220662 111944 220668
rect 111798 220623 111854 220632
rect 111904 220289 111932 220662
rect 111890 220280 111946 220289
rect 111890 220215 111946 220224
rect 112456 219434 112484 293966
rect 112180 219406 112484 219434
rect 111892 218748 111944 218754
rect 111892 218690 111944 218696
rect 111800 218000 111852 218006
rect 111798 217968 111800 217977
rect 111852 217968 111854 217977
rect 111798 217903 111854 217912
rect 111904 217705 111932 218690
rect 111890 217696 111946 217705
rect 111890 217631 111946 217640
rect 111800 216640 111852 216646
rect 111800 216582 111852 216588
rect 111812 216209 111840 216582
rect 111798 216200 111854 216209
rect 111798 216135 111854 216144
rect 111800 215280 111852 215286
rect 111798 215248 111800 215257
rect 111852 215248 111854 215257
rect 111798 215183 111854 215192
rect 111892 215212 111944 215218
rect 111892 215154 111944 215160
rect 111904 214849 111932 215154
rect 111890 214840 111946 214849
rect 111890 214775 111946 214784
rect 30288 213988 30340 213994
rect 30288 213930 30340 213936
rect 30300 133686 30328 213930
rect 111800 213920 111852 213926
rect 111798 213888 111800 213897
rect 111852 213888 111854 213897
rect 111798 213823 111854 213832
rect 111892 213852 111944 213858
rect 111892 213794 111944 213800
rect 111904 213489 111932 213794
rect 111890 213480 111946 213489
rect 111890 213415 111946 213424
rect 111798 212528 111854 212537
rect 111798 212463 111800 212472
rect 111852 212463 111854 212472
rect 111800 212434 111852 212440
rect 111892 212424 111944 212430
rect 111892 212366 111944 212372
rect 111904 212129 111932 212366
rect 111890 212120 111946 212129
rect 111890 212055 111946 212064
rect 111798 211168 111854 211177
rect 111798 211103 111800 211112
rect 111852 211103 111854 211112
rect 111800 211074 111852 211080
rect 111892 211064 111944 211070
rect 111892 211006 111944 211012
rect 111904 210769 111932 211006
rect 111890 210760 111946 210769
rect 111890 210695 111946 210704
rect 111800 209772 111852 209778
rect 111800 209714 111852 209720
rect 111812 209681 111840 209714
rect 111798 209672 111854 209681
rect 111798 209607 111854 209616
rect 111800 209092 111852 209098
rect 111800 209034 111852 209040
rect 111812 208321 111840 209034
rect 111798 208312 111854 208321
rect 111798 208247 111854 208256
rect 111984 207732 112036 207738
rect 111984 207674 112036 207680
rect 111800 206984 111852 206990
rect 111798 206952 111800 206961
rect 111852 206952 111854 206961
rect 111798 206887 111854 206896
rect 111892 206916 111944 206922
rect 111892 206858 111944 206864
rect 111904 206689 111932 206858
rect 111890 206680 111946 206689
rect 111890 206615 111946 206624
rect 111996 206145 112024 207674
rect 112076 207664 112128 207670
rect 112076 207606 112128 207612
rect 111982 206136 112038 206145
rect 111982 206071 112038 206080
rect 111800 205624 111852 205630
rect 111800 205566 111852 205572
rect 111812 205057 111840 205566
rect 111892 205556 111944 205562
rect 111892 205498 111944 205504
rect 111798 205048 111854 205057
rect 111798 204983 111854 204992
rect 111904 204785 111932 205498
rect 111890 204776 111946 204785
rect 111890 204711 111946 204720
rect 111800 204264 111852 204270
rect 111800 204206 111852 204212
rect 111812 203697 111840 204206
rect 111892 204060 111944 204066
rect 111892 204002 111944 204008
rect 111798 203688 111854 203697
rect 111798 203623 111854 203632
rect 111904 203425 111932 204002
rect 111890 203416 111946 203425
rect 111890 203351 111946 203360
rect 111800 202836 111852 202842
rect 111800 202778 111852 202784
rect 111812 202609 111840 202778
rect 111892 202768 111944 202774
rect 111892 202710 111944 202716
rect 111798 202600 111854 202609
rect 111798 202535 111854 202544
rect 111904 202065 111932 202710
rect 111890 202056 111946 202065
rect 111890 201991 111946 202000
rect 111800 201408 111852 201414
rect 111800 201350 111852 201356
rect 111812 201113 111840 201350
rect 111798 201104 111854 201113
rect 111798 201039 111854 201048
rect 112088 200705 112116 207606
rect 112180 204966 112208 219406
rect 112548 214554 112576 304438
rect 112640 233986 112668 313278
rect 112732 253026 112760 320146
rect 112720 253020 112772 253026
rect 112720 252962 112772 252968
rect 112824 248985 112852 323206
rect 112916 261118 112944 324566
rect 112904 261112 112956 261118
rect 113008 261089 113036 325722
rect 112904 261054 112956 261060
rect 112994 261080 113050 261089
rect 113100 261050 113128 325926
rect 113836 304910 113864 345102
rect 113928 307562 113956 346394
rect 115204 342916 115256 342922
rect 115204 342858 115256 342864
rect 115112 334620 115164 334626
rect 115112 334562 115164 334568
rect 114468 332920 114520 332926
rect 114468 332862 114520 332868
rect 114376 323060 114428 323066
rect 114376 323002 114428 323008
rect 114284 318844 114336 318850
rect 114284 318786 114336 318792
rect 114192 310820 114244 310826
rect 114192 310762 114244 310768
rect 113916 307556 113968 307562
rect 113916 307498 113968 307504
rect 114100 305040 114152 305046
rect 114100 304982 114152 304988
rect 113824 304904 113876 304910
rect 113824 304846 113876 304852
rect 114008 302524 114060 302530
rect 114008 302466 114060 302472
rect 113916 299532 113968 299538
rect 113916 299474 113968 299480
rect 113824 295384 113876 295390
rect 113824 295326 113876 295332
rect 112994 261015 113050 261024
rect 113088 261044 113140 261050
rect 113088 260986 113140 260992
rect 112996 260976 113048 260982
rect 112996 260918 113048 260924
rect 112904 260908 112956 260914
rect 112904 260850 112956 260856
rect 112916 260726 112944 260850
rect 113008 260834 113036 260918
rect 113008 260806 113220 260834
rect 112916 260698 113128 260726
rect 113192 260710 113220 260806
rect 112994 260536 113050 260545
rect 112994 260471 113050 260480
rect 113008 255241 113036 260471
rect 113100 256601 113128 260698
rect 113180 260704 113232 260710
rect 113180 260646 113232 260652
rect 113086 256592 113142 256601
rect 113086 256527 113142 256536
rect 112994 255232 113050 255241
rect 112994 255167 113050 255176
rect 112810 248976 112866 248985
rect 112810 248911 112866 248920
rect 112904 246356 112956 246362
rect 112904 246298 112956 246304
rect 112628 233980 112680 233986
rect 112628 233922 112680 233928
rect 112812 232552 112864 232558
rect 112812 232494 112864 232500
rect 112824 224466 112852 232494
rect 112916 231849 112944 246298
rect 112902 231840 112958 231849
rect 112902 231775 112958 231784
rect 112904 231124 112956 231130
rect 112904 231066 112956 231072
rect 112812 224460 112864 224466
rect 112812 224402 112864 224408
rect 112916 224210 112944 231066
rect 112996 224460 113048 224466
rect 112996 224402 113048 224408
rect 112824 224182 112944 224210
rect 112628 220108 112680 220114
rect 112628 220050 112680 220056
rect 112640 219337 112668 220050
rect 112626 219328 112682 219337
rect 112626 219263 112682 219272
rect 112824 219065 112852 224182
rect 113008 219434 113036 224402
rect 112916 219406 113036 219434
rect 112810 219056 112866 219065
rect 112810 218991 112866 219000
rect 112628 217320 112680 217326
rect 112628 217262 112680 217268
rect 112364 214526 112576 214554
rect 112364 208185 112392 214526
rect 112640 213602 112668 217262
rect 112916 216617 112944 219406
rect 112902 216608 112958 216617
rect 112902 216543 112958 216552
rect 112720 215960 112772 215966
rect 112720 215902 112772 215908
rect 112456 213574 112668 213602
rect 112456 209409 112484 213574
rect 112732 209774 112760 215902
rect 112732 209746 112944 209774
rect 112442 209400 112498 209409
rect 112442 209335 112498 209344
rect 112350 208176 112406 208185
rect 112350 208111 112406 208120
rect 112628 207800 112680 207806
rect 112628 207742 112680 207748
rect 112180 204938 112392 204966
rect 112260 202156 112312 202162
rect 112260 202098 112312 202104
rect 112074 200696 112130 200705
rect 112074 200631 112130 200640
rect 111892 200116 111944 200122
rect 111892 200058 111944 200064
rect 111800 200048 111852 200054
rect 111800 199990 111852 199996
rect 111812 199753 111840 199990
rect 111798 199744 111854 199753
rect 111798 199679 111854 199688
rect 111904 199345 111932 200058
rect 111890 199336 111946 199345
rect 111890 199271 111946 199280
rect 111800 198688 111852 198694
rect 111800 198630 111852 198636
rect 111812 198393 111840 198630
rect 111798 198384 111854 198393
rect 111798 198319 111854 198328
rect 111800 197328 111852 197334
rect 112272 197305 112300 202098
rect 112364 200114 112392 204938
rect 112364 200086 112484 200114
rect 111800 197270 111852 197276
rect 112258 197296 112314 197305
rect 111812 196625 111840 197270
rect 112258 197231 112314 197240
rect 111798 196616 111854 196625
rect 111798 196551 111854 196560
rect 111800 195968 111852 195974
rect 111800 195910 111852 195916
rect 111812 195673 111840 195910
rect 111892 195900 111944 195906
rect 111892 195842 111944 195848
rect 111798 195664 111854 195673
rect 111798 195599 111854 195608
rect 111904 195265 111932 195842
rect 111890 195256 111946 195265
rect 111890 195191 111946 195200
rect 111800 194540 111852 194546
rect 111800 194482 111852 194488
rect 111812 194313 111840 194482
rect 111892 194472 111944 194478
rect 111892 194414 111944 194420
rect 111798 194304 111854 194313
rect 111798 194239 111854 194248
rect 111904 193769 111932 194414
rect 111890 193760 111946 193769
rect 111890 193695 111946 193704
rect 111892 193180 111944 193186
rect 111892 193122 111944 193128
rect 111800 193112 111852 193118
rect 111800 193054 111852 193060
rect 111812 192953 111840 193054
rect 111798 192944 111854 192953
rect 111798 192879 111854 192888
rect 111904 192545 111932 193122
rect 111890 192536 111946 192545
rect 111890 192471 111946 192480
rect 111800 191752 111852 191758
rect 111800 191694 111852 191700
rect 111812 191593 111840 191694
rect 111798 191584 111854 191593
rect 111798 191519 111854 191528
rect 111800 191208 111852 191214
rect 111800 191150 111852 191156
rect 111812 190913 111840 191150
rect 111798 190904 111854 190913
rect 111798 190839 111854 190848
rect 111892 190460 111944 190466
rect 111892 190402 111944 190408
rect 111800 190392 111852 190398
rect 111800 190334 111852 190340
rect 111812 190233 111840 190334
rect 111798 190224 111854 190233
rect 111798 190159 111854 190168
rect 111904 189825 111932 190402
rect 111890 189816 111946 189825
rect 111890 189751 111946 189760
rect 111892 189032 111944 189038
rect 111892 188974 111944 188980
rect 111800 188964 111852 188970
rect 111800 188906 111852 188912
rect 111812 188873 111840 188906
rect 111798 188864 111854 188873
rect 111798 188799 111854 188808
rect 111904 188465 111932 188974
rect 111890 188456 111946 188465
rect 111890 188391 111946 188400
rect 111892 187672 111944 187678
rect 111892 187614 111944 187620
rect 111800 187604 111852 187610
rect 111800 187546 111852 187552
rect 111812 187513 111840 187546
rect 111798 187504 111854 187513
rect 111798 187439 111854 187448
rect 111904 187105 111932 187614
rect 111890 187096 111946 187105
rect 111890 187031 111946 187040
rect 111800 186312 111852 186318
rect 111800 186254 111852 186260
rect 111812 185745 111840 186254
rect 111798 185736 111854 185745
rect 111798 185671 111854 185680
rect 111892 184884 111944 184890
rect 111892 184826 111944 184832
rect 111800 184816 111852 184822
rect 111800 184758 111852 184764
rect 111812 184657 111840 184758
rect 111798 184648 111854 184657
rect 111798 184583 111854 184592
rect 111904 184385 111932 184826
rect 111890 184376 111946 184385
rect 111890 184311 111946 184320
rect 111800 183524 111852 183530
rect 111800 183466 111852 183472
rect 111812 183025 111840 183466
rect 111798 183016 111854 183025
rect 111798 182951 111854 182960
rect 111800 182164 111852 182170
rect 111800 182106 111852 182112
rect 111812 182073 111840 182106
rect 111798 182064 111854 182073
rect 111798 181999 111854 182008
rect 111800 181824 111852 181830
rect 111800 181766 111852 181772
rect 111812 181529 111840 181766
rect 111798 181520 111854 181529
rect 111798 181455 111854 181464
rect 111892 180804 111944 180810
rect 111892 180746 111944 180752
rect 111800 180736 111852 180742
rect 111800 180678 111852 180684
rect 111812 180577 111840 180678
rect 111798 180568 111854 180577
rect 111798 180503 111854 180512
rect 111904 180305 111932 180746
rect 111890 180296 111946 180305
rect 111890 180231 111946 180240
rect 111892 179376 111944 179382
rect 111892 179318 111944 179324
rect 111800 179308 111852 179314
rect 111800 179250 111852 179256
rect 111812 179217 111840 179250
rect 111798 179208 111854 179217
rect 111798 179143 111854 179152
rect 111904 178945 111932 179318
rect 111890 178936 111946 178945
rect 111890 178871 111946 178880
rect 111984 177336 112036 177342
rect 111984 177278 112036 177284
rect 111800 176656 111852 176662
rect 111800 176598 111852 176604
rect 111812 176497 111840 176598
rect 111892 176588 111944 176594
rect 111892 176530 111944 176536
rect 111798 176488 111854 176497
rect 111798 176423 111854 176432
rect 111904 176225 111932 176530
rect 111890 176216 111946 176225
rect 111890 176151 111946 176160
rect 111996 175273 112024 177278
rect 111982 175264 112038 175273
rect 111982 175199 112038 175208
rect 112456 174865 112484 200086
rect 112536 195288 112588 195294
rect 112536 195230 112588 195236
rect 112548 183569 112576 195230
rect 112640 190454 112668 207742
rect 112916 197985 112944 209746
rect 112996 200796 113048 200802
rect 112996 200738 113048 200744
rect 112902 197976 112958 197985
rect 112902 197911 112958 197920
rect 113008 195294 113036 200738
rect 112996 195288 113048 195294
rect 112996 195230 113048 195236
rect 112904 193860 112956 193866
rect 112904 193802 112956 193808
rect 112640 190426 112760 190454
rect 112534 183560 112590 183569
rect 112534 183495 112590 183504
rect 112732 177993 112760 190426
rect 112916 186289 112944 193802
rect 112902 186280 112958 186289
rect 112902 186215 112958 186224
rect 112812 184204 112864 184210
rect 112812 184146 112864 184152
rect 112718 177984 112774 177993
rect 112718 177919 112774 177928
rect 112824 177585 112852 184146
rect 113836 181830 113864 295326
rect 113928 191214 113956 299474
rect 114020 198694 114048 302466
rect 114112 204066 114140 304982
rect 114204 218006 114232 310762
rect 114296 238542 114324 318786
rect 114388 248334 114416 323002
rect 114480 273086 114508 332862
rect 115124 297974 115152 334562
rect 115216 299198 115244 342858
rect 115848 342304 115900 342310
rect 115848 342246 115900 342252
rect 115756 331288 115808 331294
rect 115756 331230 115808 331236
rect 115664 329860 115716 329866
rect 115664 329802 115716 329808
rect 115572 321632 115624 321638
rect 115572 321574 115624 321580
rect 115480 316328 115532 316334
rect 115480 316270 115532 316276
rect 115388 313404 115440 313410
rect 115388 313346 115440 313352
rect 115296 303884 115348 303890
rect 115296 303826 115348 303832
rect 115204 299192 115256 299198
rect 115204 299134 115256 299140
rect 115112 297968 115164 297974
rect 115112 297910 115164 297916
rect 115204 296744 115256 296750
rect 115204 296686 115256 296692
rect 114468 273080 114520 273086
rect 114468 273022 114520 273028
rect 114376 248328 114428 248334
rect 114376 248270 114428 248276
rect 114284 238536 114336 238542
rect 114284 238478 114336 238484
rect 114192 218000 114244 218006
rect 114192 217942 114244 217948
rect 114100 204060 114152 204066
rect 114100 204002 114152 204008
rect 114008 198688 114060 198694
rect 114008 198630 114060 198636
rect 113916 191208 113968 191214
rect 113916 191150 113968 191156
rect 115216 184822 115244 296686
rect 115308 201414 115336 303826
rect 115400 226030 115428 313346
rect 115492 232966 115520 316270
rect 115584 246974 115612 321574
rect 115676 266286 115704 329802
rect 115768 269006 115796 331230
rect 115860 298858 115888 342246
rect 116596 309058 116624 346462
rect 116688 311778 116716 347754
rect 118240 347064 118292 347070
rect 118240 347006 118292 347012
rect 117136 340944 117188 340950
rect 117136 340886 117188 340892
rect 117044 327140 117096 327146
rect 117044 327082 117096 327088
rect 116952 321700 117004 321706
rect 116952 321642 117004 321648
rect 116676 311772 116728 311778
rect 116676 311714 116728 311720
rect 116860 311160 116912 311166
rect 116860 311102 116912 311108
rect 116584 309052 116636 309058
rect 116584 308994 116636 309000
rect 116768 303748 116820 303754
rect 116768 303690 116820 303696
rect 115848 298852 115900 298858
rect 115848 298794 115900 298800
rect 116676 296812 116728 296818
rect 116676 296754 116728 296760
rect 116584 292596 116636 292602
rect 116584 292538 116636 292544
rect 115756 269000 115808 269006
rect 115756 268942 115808 268948
rect 115664 266280 115716 266286
rect 115664 266222 115716 266228
rect 115572 246968 115624 246974
rect 115572 246910 115624 246916
rect 115480 232960 115532 232966
rect 115480 232902 115532 232908
rect 115388 226024 115440 226030
rect 115388 225966 115440 225972
rect 115296 201408 115348 201414
rect 115296 201350 115348 201356
rect 115204 184816 115256 184822
rect 115204 184758 115256 184764
rect 113824 181824 113876 181830
rect 113824 181766 113876 181772
rect 112810 177576 112866 177585
rect 112810 177511 112866 177520
rect 112442 174856 112498 174865
rect 112442 174791 112498 174800
rect 111800 173868 111852 173874
rect 111800 173810 111852 173816
rect 111812 173777 111840 173810
rect 111892 173800 111944 173806
rect 111798 173768 111854 173777
rect 111892 173742 111944 173748
rect 111798 173703 111854 173712
rect 111904 173369 111932 173742
rect 111890 173360 111946 173369
rect 111890 173295 111946 173304
rect 111800 172508 111852 172514
rect 111800 172450 111852 172456
rect 111812 172145 111840 172450
rect 111798 172136 111854 172145
rect 111798 172071 111854 172080
rect 111892 171080 111944 171086
rect 111798 171048 111854 171057
rect 111892 171022 111944 171028
rect 111798 170983 111800 170992
rect 111852 170983 111854 170992
rect 111800 170954 111852 170960
rect 111904 170649 111932 171022
rect 116596 171018 116624 292538
rect 116688 184890 116716 296754
rect 116780 202774 116808 303690
rect 116872 227662 116900 311102
rect 116964 245546 116992 321642
rect 117056 260778 117084 327082
rect 117148 293894 117176 340886
rect 117228 338768 117280 338774
rect 117228 338710 117280 338716
rect 117240 303550 117268 338710
rect 117964 333260 118016 333266
rect 117964 333202 118016 333208
rect 117976 313206 118004 333202
rect 118056 327208 118108 327214
rect 118056 327150 118108 327156
rect 117964 313200 118016 313206
rect 117964 313142 118016 313148
rect 117964 307828 118016 307834
rect 117964 307770 118016 307776
rect 117228 303544 117280 303550
rect 117228 303486 117280 303492
rect 117136 293888 117188 293894
rect 117136 293830 117188 293836
rect 117044 260772 117096 260778
rect 117044 260714 117096 260720
rect 116952 245540 117004 245546
rect 116952 245482 117004 245488
rect 116860 227656 116912 227662
rect 116860 227598 116912 227604
rect 117976 211070 118004 307770
rect 118068 259418 118096 327150
rect 118148 319456 118200 319462
rect 118148 319398 118200 319404
rect 118056 259412 118108 259418
rect 118056 259354 118108 259360
rect 118160 259350 118188 319398
rect 118252 309126 118280 347006
rect 119344 343664 119396 343670
rect 119344 343606 119396 343612
rect 118240 309120 118292 309126
rect 118240 309062 118292 309068
rect 119356 300694 119384 343606
rect 119448 310418 119476 347890
rect 119528 347880 119580 347886
rect 119528 347822 119580 347828
rect 119540 310486 119568 347822
rect 122104 345704 122156 345710
rect 122104 345646 122156 345652
rect 120724 343732 120776 343738
rect 120724 343674 120776 343680
rect 119896 337408 119948 337414
rect 119896 337350 119948 337356
rect 119804 335640 119856 335646
rect 119804 335582 119856 335588
rect 119712 317484 119764 317490
rect 119712 317426 119764 317432
rect 119620 310616 119672 310622
rect 119620 310558 119672 310564
rect 119528 310480 119580 310486
rect 119528 310422 119580 310428
rect 119436 310412 119488 310418
rect 119436 310354 119488 310360
rect 119528 304292 119580 304298
rect 119528 304234 119580 304240
rect 119436 300892 119488 300898
rect 119436 300834 119488 300840
rect 119344 300688 119396 300694
rect 119344 300630 119396 300636
rect 119344 292664 119396 292670
rect 119344 292606 119396 292612
rect 118148 259344 118200 259350
rect 118148 259286 118200 259292
rect 117964 211064 118016 211070
rect 117964 211006 118016 211012
rect 116768 202768 116820 202774
rect 116768 202710 116820 202716
rect 116676 184884 116728 184890
rect 116676 184826 116728 184832
rect 119356 173806 119384 292606
rect 119448 194478 119476 300834
rect 119540 202842 119568 304234
rect 119632 231130 119660 310558
rect 119724 240786 119752 317426
rect 119816 281450 119844 335582
rect 119908 292466 119936 337350
rect 120736 302122 120764 343674
rect 121184 341012 121236 341018
rect 121184 340954 121236 340960
rect 121092 327276 121144 327282
rect 121092 327218 121144 327224
rect 121000 324420 121052 324426
rect 121000 324362 121052 324368
rect 120724 302116 120776 302122
rect 120724 302058 120776 302064
rect 120816 300960 120868 300966
rect 120816 300902 120868 300908
rect 120724 292732 120776 292738
rect 120724 292674 120776 292680
rect 119896 292460 119948 292466
rect 119896 292402 119948 292408
rect 119804 281444 119856 281450
rect 119804 281386 119856 281392
rect 119712 240780 119764 240786
rect 119712 240722 119764 240728
rect 119620 231124 119672 231130
rect 119620 231066 119672 231072
rect 119528 202836 119580 202842
rect 119528 202778 119580 202784
rect 119436 194472 119488 194478
rect 119436 194414 119488 194420
rect 120736 173874 120764 292674
rect 120828 194546 120856 300902
rect 120908 294092 120960 294098
rect 120908 294034 120960 294040
rect 120920 207806 120948 294034
rect 121012 253774 121040 324362
rect 121104 257990 121132 327218
rect 121196 293962 121224 340954
rect 122116 306270 122144 345646
rect 122564 329928 122616 329934
rect 122564 329870 122616 329876
rect 122472 324488 122524 324494
rect 122472 324430 122524 324436
rect 122380 318096 122432 318102
rect 122380 318038 122432 318044
rect 122288 317552 122340 317558
rect 122288 317494 122340 317500
rect 122196 314696 122248 314702
rect 122196 314638 122248 314644
rect 122104 306264 122156 306270
rect 122104 306206 122156 306212
rect 122104 294160 122156 294166
rect 122104 294102 122156 294108
rect 121184 293956 121236 293962
rect 121184 293898 121236 293904
rect 121092 257984 121144 257990
rect 121092 257926 121144 257932
rect 121000 253768 121052 253774
rect 121000 253710 121052 253716
rect 120908 207800 120960 207806
rect 120908 207742 120960 207748
rect 120816 194540 120868 194546
rect 120816 194482 120868 194488
rect 122116 176594 122144 294102
rect 122208 227730 122236 314638
rect 122300 235958 122328 317494
rect 122392 244254 122420 318038
rect 122484 252550 122512 324430
rect 122576 267646 122604 329870
rect 122668 311846 122696 347958
rect 123484 343800 123536 343806
rect 123484 343742 123536 343748
rect 122656 311840 122708 311846
rect 122656 311782 122708 311788
rect 123496 300762 123524 343742
rect 124036 341080 124088 341086
rect 124036 341022 124088 341028
rect 123944 324556 123996 324562
rect 123944 324498 123996 324504
rect 123852 314764 123904 314770
rect 123852 314706 123904 314712
rect 123760 312180 123812 312186
rect 123760 312122 123812 312128
rect 123576 307896 123628 307902
rect 123576 307838 123628 307844
rect 123484 300756 123536 300762
rect 123484 300698 123536 300704
rect 123484 298172 123536 298178
rect 123484 298114 123536 298120
rect 122564 267640 122616 267646
rect 122564 267582 122616 267588
rect 122472 252544 122524 252550
rect 122472 252486 122524 252492
rect 122380 244248 122432 244254
rect 122380 244190 122432 244196
rect 122288 235952 122340 235958
rect 122288 235894 122340 235900
rect 122196 227724 122248 227730
rect 122196 227666 122248 227672
rect 123496 187610 123524 298114
rect 123588 212430 123616 307838
rect 123668 298784 123720 298790
rect 123668 298726 123720 298732
rect 123576 212424 123628 212430
rect 123576 212366 123628 212372
rect 123680 204270 123708 298726
rect 123772 220726 123800 312122
rect 123864 229022 123892 314706
rect 123956 253842 123984 324498
rect 124048 295254 124076 341022
rect 125140 338156 125192 338162
rect 125140 338098 125192 338104
rect 125048 314832 125100 314838
rect 125048 314774 125100 314780
rect 124956 309188 125008 309194
rect 124956 309130 125008 309136
rect 124864 305108 124916 305114
rect 124864 305050 124916 305056
rect 124036 295248 124088 295254
rect 124036 295190 124088 295196
rect 123944 253836 123996 253842
rect 123944 253778 123996 253784
rect 123852 229016 123904 229022
rect 123852 228958 123904 228964
rect 123760 220720 123812 220726
rect 123760 220662 123812 220668
rect 124876 205562 124904 305050
rect 124968 212498 124996 309130
rect 125060 229090 125088 314774
rect 125152 286958 125180 338098
rect 126256 313274 126284 349114
rect 131764 343868 131816 343874
rect 131764 343810 131816 343816
rect 128176 341148 128228 341154
rect 128176 341090 128228 341096
rect 126796 338224 126848 338230
rect 126796 338166 126848 338172
rect 126704 321768 126756 321774
rect 126704 321710 126756 321716
rect 126612 316124 126664 316130
rect 126612 316066 126664 316072
rect 126244 313268 126296 313274
rect 126244 313210 126296 313216
rect 126520 311976 126572 311982
rect 126520 311918 126572 311924
rect 126428 309256 126480 309262
rect 126428 309198 126480 309204
rect 126336 306468 126388 306474
rect 126336 306410 126388 306416
rect 126244 302320 126296 302326
rect 126244 302262 126296 302268
rect 125140 286952 125192 286958
rect 125140 286894 125192 286900
rect 125048 229084 125100 229090
rect 125048 229026 125100 229032
rect 124956 212492 125008 212498
rect 124956 212434 125008 212440
rect 124864 205556 124916 205562
rect 124864 205498 124916 205504
rect 123668 204264 123720 204270
rect 123668 204206 123720 204212
rect 126256 197334 126284 302262
rect 126348 205630 126376 306410
rect 126440 213858 126468 309198
rect 126532 222086 126560 311918
rect 126624 230382 126652 316066
rect 126716 247042 126744 321710
rect 126808 288318 126836 338166
rect 128084 335436 128136 335442
rect 128084 335378 128136 335384
rect 127992 318912 128044 318918
rect 127992 318854 128044 318860
rect 127900 314900 127952 314906
rect 127900 314842 127952 314848
rect 127808 312044 127860 312050
rect 127808 311986 127860 311992
rect 127716 309324 127768 309330
rect 127716 309266 127768 309272
rect 127624 305176 127676 305182
rect 127624 305118 127676 305124
rect 126796 288312 126848 288318
rect 126796 288254 126848 288260
rect 126704 247036 126756 247042
rect 126704 246978 126756 246984
rect 126612 230376 126664 230382
rect 126612 230318 126664 230324
rect 126520 222080 126572 222086
rect 126520 222022 126572 222028
rect 126428 213852 126480 213858
rect 126428 213794 126480 213800
rect 127636 207738 127664 305118
rect 127728 213926 127756 309266
rect 127820 222154 127848 311986
rect 127912 230450 127940 314842
rect 128004 238746 128032 318854
rect 128096 281518 128124 335378
rect 128188 295322 128216 341090
rect 129372 332716 129424 332722
rect 129372 332658 129424 332664
rect 129280 331356 129332 331362
rect 129280 331298 129332 331304
rect 129188 302388 129240 302394
rect 129188 302330 129240 302336
rect 129096 295520 129148 295526
rect 129096 295462 129148 295468
rect 129004 295452 129056 295458
rect 129004 295394 129056 295400
rect 128176 295316 128228 295322
rect 128176 295258 128228 295264
rect 128084 281512 128136 281518
rect 128084 281454 128136 281460
rect 127992 238740 128044 238746
rect 127992 238682 128044 238688
rect 127900 230444 127952 230450
rect 127900 230386 127952 230392
rect 127808 222148 127860 222154
rect 127808 222090 127860 222096
rect 127716 213920 127768 213926
rect 127716 213862 127768 213868
rect 127624 207732 127676 207738
rect 127624 207674 127676 207680
rect 126336 205624 126388 205630
rect 126336 205566 126388 205572
rect 126244 197328 126296 197334
rect 126244 197270 126296 197276
rect 123484 187604 123536 187610
rect 123484 187546 123536 187552
rect 129016 180810 129044 295394
rect 129004 180804 129056 180810
rect 129004 180746 129056 180752
rect 129108 180742 129136 295462
rect 129200 215966 129228 302330
rect 129292 267714 129320 331298
rect 129384 274582 129412 332658
rect 130844 323128 130896 323134
rect 130844 323070 130896 323076
rect 130752 318980 130804 318986
rect 130752 318922 130804 318928
rect 130660 316192 130712 316198
rect 130660 316134 130712 316140
rect 130568 313472 130620 313478
rect 130568 313414 130620 313420
rect 130476 309392 130528 309398
rect 130476 309334 130528 309340
rect 130384 306536 130436 306542
rect 130384 306478 130436 306484
rect 129372 274576 129424 274582
rect 129372 274518 129424 274524
rect 129280 267708 129332 267714
rect 129280 267650 129332 267656
rect 129188 215960 129240 215966
rect 129188 215902 129240 215908
rect 130396 206922 130424 306478
rect 130488 215218 130516 309334
rect 130580 223514 130608 313414
rect 130672 231810 130700 316134
rect 130764 240038 130792 318922
rect 130856 248402 130884 323070
rect 131776 300830 131804 343810
rect 133236 339516 133288 339522
rect 133236 339458 133288 339464
rect 132224 334144 132276 334150
rect 132224 334086 132276 334092
rect 132132 331424 132184 331430
rect 132132 331366 132184 331372
rect 132040 328568 132092 328574
rect 132040 328510 132092 328516
rect 131948 325848 132000 325854
rect 131948 325790 132000 325796
rect 131764 300824 131816 300830
rect 131764 300766 131816 300772
rect 131856 299600 131908 299606
rect 131856 299542 131908 299548
rect 131764 295588 131816 295594
rect 131764 295530 131816 295536
rect 130844 248396 130896 248402
rect 130844 248338 130896 248344
rect 130752 240032 130804 240038
rect 130752 239974 130804 239980
rect 130660 231804 130712 231810
rect 130660 231746 130712 231752
rect 130568 223508 130620 223514
rect 130568 223450 130620 223456
rect 130476 215212 130528 215218
rect 130476 215154 130528 215160
rect 130384 206916 130436 206922
rect 130384 206858 130436 206864
rect 129096 180736 129148 180742
rect 129096 180678 129148 180684
rect 131776 177342 131804 295530
rect 131868 190398 131896 299542
rect 131960 253910 131988 325790
rect 132052 260846 132080 328510
rect 132144 269074 132172 331366
rect 132236 275942 132264 334086
rect 133144 312112 133196 312118
rect 133144 312054 133196 312060
rect 132224 275936 132276 275942
rect 132224 275878 132276 275884
rect 132132 269068 132184 269074
rect 132132 269010 132184 269016
rect 132040 260840 132092 260846
rect 132040 260782 132092 260788
rect 131948 253904 132000 253910
rect 131948 253846 132000 253852
rect 133156 220794 133184 312054
rect 133248 291106 133276 339458
rect 133604 336864 133656 336870
rect 133604 336806 133656 336812
rect 133512 335504 133564 335510
rect 133512 335446 133564 335452
rect 133420 320340 133472 320346
rect 133420 320282 133472 320288
rect 133328 320272 133380 320278
rect 133328 320214 133380 320220
rect 133236 291100 133288 291106
rect 133236 291042 133288 291048
rect 133236 282192 133288 282198
rect 133236 282134 133288 282140
rect 133144 220788 133196 220794
rect 133144 220730 133196 220736
rect 133248 191758 133276 282134
rect 133340 241466 133368 320214
rect 133432 242894 133460 320282
rect 133524 280090 133552 335446
rect 133616 282878 133644 336806
rect 133604 282872 133656 282878
rect 133604 282814 133656 282820
rect 133512 280084 133564 280090
rect 133512 280026 133564 280032
rect 133420 242888 133472 242894
rect 133420 242830 133472 242836
rect 133328 241460 133380 241466
rect 133328 241402 133380 241408
rect 133236 191752 133288 191758
rect 133236 191694 133288 191700
rect 131856 190392 131908 190398
rect 131856 190334 131908 190340
rect 131764 177336 131816 177342
rect 131764 177278 131816 177284
rect 122104 176588 122156 176594
rect 122104 176530 122156 176536
rect 120724 173868 120776 173874
rect 120724 173810 120776 173816
rect 119344 173800 119396 173806
rect 119344 173742 119396 173748
rect 116584 171012 116636 171018
rect 116584 170954 116636 170960
rect 111890 170640 111946 170649
rect 111890 170575 111946 170584
rect 30288 133680 30340 133686
rect 30288 133622 30340 133628
rect 30196 133612 30248 133618
rect 30196 133554 30248 133560
rect 30012 133476 30064 133482
rect 30012 133418 30064 133424
rect 29828 133340 29880 133346
rect 29828 133282 29880 133288
rect 29644 133272 29696 133278
rect 29644 133214 29696 133220
rect 6920 133204 6972 133210
rect 6920 133146 6972 133152
rect 3422 110664 3478 110673
rect 3422 110599 3478 110608
rect 3436 110498 3464 110599
rect 3424 110492 3476 110498
rect 3424 110434 3476 110440
rect 22744 110492 22796 110498
rect 22744 110434 22796 110440
rect 3422 97608 3478 97617
rect 3422 97543 3478 97552
rect 3436 96694 3464 97543
rect 3424 96688 3476 96694
rect 3424 96630 3476 96636
rect 3422 84688 3478 84697
rect 3422 84623 3478 84632
rect 3436 25770 3464 84623
rect 3514 71632 3570 71641
rect 3514 71567 3570 71576
rect 3424 25764 3476 25770
rect 3424 25706 3476 25712
rect 3528 25702 3556 71567
rect 3606 58576 3662 58585
rect 3606 58511 3662 58520
rect 3516 25696 3568 25702
rect 3516 25638 3568 25644
rect 3620 25498 3648 58511
rect 3698 45520 3754 45529
rect 3698 45455 3754 45464
rect 3712 25566 3740 45455
rect 3790 32464 3846 32473
rect 3790 32399 3846 32408
rect 3804 25634 3832 32399
rect 3792 25628 3844 25634
rect 3792 25570 3844 25576
rect 3700 25560 3752 25566
rect 3700 25502 3752 25508
rect 3608 25492 3660 25498
rect 3608 25434 3660 25440
rect 22756 24857 22784 110434
rect 24124 96688 24176 96694
rect 24124 96630 24176 96636
rect 24136 25430 24164 96630
rect 134536 50522 134564 397462
rect 134720 397254 134748 565830
rect 134800 484424 134852 484430
rect 134800 484366 134852 484372
rect 134708 397248 134760 397254
rect 134708 397190 134760 397196
rect 134812 365566 134840 484366
rect 134800 365560 134852 365566
rect 134800 365502 134852 365508
rect 134708 339584 134760 339590
rect 134708 339526 134760 339532
rect 134616 313540 134668 313546
rect 134616 313482 134668 313488
rect 134628 224874 134656 313482
rect 134720 289746 134748 339526
rect 134708 289740 134760 289746
rect 134708 289682 134760 289688
rect 134616 224868 134668 224874
rect 134616 224810 134668 224816
rect 134616 160812 134668 160818
rect 134616 160754 134668 160760
rect 134524 50516 134576 50522
rect 134524 50458 134576 50464
rect 134628 48385 134656 160754
rect 134708 136672 134760 136678
rect 134708 136614 134760 136620
rect 134720 51338 134748 136614
rect 135260 121440 135312 121446
rect 135260 121382 135312 121388
rect 135272 120873 135300 121382
rect 135258 120864 135314 120873
rect 135258 120799 135314 120808
rect 135444 118652 135496 118658
rect 135444 118594 135496 118600
rect 135456 118289 135484 118594
rect 135442 118280 135498 118289
rect 135442 118215 135498 118224
rect 135812 87372 135864 87378
rect 135812 87314 135864 87320
rect 135260 86896 135312 86902
rect 135258 86864 135260 86873
rect 135312 86864 135314 86873
rect 135258 86799 135314 86808
rect 135824 84833 135852 87314
rect 135810 84824 135866 84833
rect 135810 84759 135866 84768
rect 135720 72480 135772 72486
rect 135720 72422 135772 72428
rect 135352 71664 135404 71670
rect 135350 71632 135352 71641
rect 135404 71632 135406 71641
rect 135350 71567 135406 71576
rect 135732 68921 135760 72422
rect 135718 68912 135774 68921
rect 135718 68847 135774 68856
rect 135628 62076 135680 62082
rect 135628 62018 135680 62024
rect 135640 61577 135668 62018
rect 135626 61568 135682 61577
rect 135626 61503 135682 61512
rect 135260 56432 135312 56438
rect 135258 56400 135260 56409
rect 135312 56400 135314 56409
rect 135258 56335 135314 56344
rect 135916 51406 135944 605814
rect 135996 496120 136048 496126
rect 135996 496062 136048 496068
rect 136008 371006 136036 496062
rect 136088 476128 136140 476134
rect 136088 476070 136140 476076
rect 135996 371000 136048 371006
rect 135996 370942 136048 370948
rect 136100 361282 136128 476070
rect 136088 361276 136140 361282
rect 136088 361218 136140 361224
rect 136180 346588 136232 346594
rect 136180 346530 136232 346536
rect 135996 345092 136048 345098
rect 135996 345034 136048 345040
rect 136008 51474 136036 345034
rect 136192 306338 136220 346530
rect 136180 306332 136232 306338
rect 136180 306274 136232 306280
rect 136088 305652 136140 305658
rect 136088 305594 136140 305600
rect 136100 237386 136128 305594
rect 136088 237380 136140 237386
rect 136088 237322 136140 237328
rect 136546 130520 136602 130529
rect 136546 130455 136602 130464
rect 136560 130422 136588 130455
rect 136548 130416 136600 130422
rect 136548 130358 136600 130364
rect 136546 127936 136602 127945
rect 136546 127871 136602 127880
rect 136560 127634 136588 127871
rect 136548 127628 136600 127634
rect 136548 127570 136600 127576
rect 136548 125588 136600 125594
rect 136548 125530 136600 125536
rect 136560 125497 136588 125530
rect 136546 125488 136602 125497
rect 136546 125423 136602 125432
rect 136180 124160 136232 124166
rect 136180 124102 136232 124108
rect 136192 123593 136220 124102
rect 136178 123584 136234 123593
rect 136178 123519 136234 123528
rect 136548 115932 136600 115938
rect 136548 115874 136600 115880
rect 136560 115569 136588 115874
rect 136546 115560 136602 115569
rect 136546 115495 136602 115504
rect 136548 113144 136600 113150
rect 136548 113086 136600 113092
rect 136560 112849 136588 113086
rect 136546 112840 136602 112849
rect 136546 112775 136602 112784
rect 136548 110424 136600 110430
rect 136548 110366 136600 110372
rect 136560 110265 136588 110366
rect 136546 110256 136602 110265
rect 136546 110191 136602 110200
rect 136548 107636 136600 107642
rect 136548 107578 136600 107584
rect 136560 107545 136588 107578
rect 136546 107536 136602 107545
rect 136546 107471 136602 107480
rect 136548 104848 136600 104854
rect 136546 104816 136548 104825
rect 136600 104816 136602 104825
rect 136546 104751 136602 104760
rect 136180 103488 136232 103494
rect 136180 103430 136232 103436
rect 136192 102921 136220 103430
rect 136178 102912 136234 102921
rect 136178 102847 136234 102856
rect 136180 100700 136232 100706
rect 136180 100642 136232 100648
rect 136192 100201 136220 100642
rect 136178 100192 136234 100201
rect 136178 100127 136234 100136
rect 136548 96280 136600 96286
rect 136548 96222 136600 96228
rect 136560 95169 136588 96222
rect 136546 95160 136602 95169
rect 136546 95095 136602 95104
rect 136088 92472 136140 92478
rect 136086 92440 136088 92449
rect 136140 92440 136142 92449
rect 136086 92375 136142 92384
rect 136548 89684 136600 89690
rect 136548 89626 136600 89632
rect 136560 89593 136588 89626
rect 136546 89584 136602 89593
rect 136546 89519 136602 89528
rect 136548 82272 136600 82278
rect 136546 82240 136548 82249
rect 136600 82240 136602 82249
rect 136546 82175 136602 82184
rect 136088 79756 136140 79762
rect 136088 79698 136140 79704
rect 136100 79665 136128 79698
rect 136086 79656 136142 79665
rect 136086 79591 136142 79600
rect 136548 77104 136600 77110
rect 136546 77072 136548 77081
rect 136600 77072 136602 77081
rect 136546 77007 136602 77016
rect 136546 73808 136602 73817
rect 136546 73743 136548 73752
rect 136600 73743 136602 73752
rect 136548 73714 136600 73720
rect 136088 66224 136140 66230
rect 136086 66192 136088 66201
rect 136140 66192 136142 66201
rect 136086 66127 136142 66136
rect 136548 64184 136600 64190
rect 136546 64152 136548 64161
rect 136600 64152 136602 64161
rect 136546 64087 136602 64096
rect 136548 59016 136600 59022
rect 136546 58984 136548 58993
rect 136600 58984 136602 58993
rect 136546 58919 136602 58928
rect 136548 53780 136600 53786
rect 136548 53722 136600 53728
rect 136560 53553 136588 53722
rect 136546 53544 136602 53553
rect 136546 53479 136602 53488
rect 136652 52018 136680 703582
rect 137664 703474 137692 703582
rect 137806 703520 137918 704960
rect 154090 703520 154202 704960
rect 170282 703520 170394 704960
rect 186474 703520 186586 704960
rect 202758 703520 202870 704960
rect 218072 703582 218836 703610
rect 137848 703474 137876 703520
rect 137664 703446 137876 703474
rect 154132 702434 154160 703520
rect 170324 702434 170352 703520
rect 153212 702406 154160 702434
rect 169772 702406 170352 702434
rect 142804 700596 142856 700602
rect 142804 700538 142856 700544
rect 138664 700392 138716 700398
rect 138664 700334 138716 700340
rect 137284 568676 137336 568682
rect 137284 568618 137336 568624
rect 137296 398546 137324 568618
rect 137376 539640 137428 539646
rect 137376 539582 137428 539588
rect 137284 398540 137336 398546
rect 137284 398482 137336 398488
rect 137388 387666 137416 539582
rect 137468 488572 137520 488578
rect 137468 488514 137520 488520
rect 137376 387660 137428 387666
rect 137376 387602 137428 387608
rect 137480 366926 137508 488514
rect 137560 485920 137612 485926
rect 137560 485862 137612 485868
rect 137468 366920 137520 366926
rect 137468 366862 137520 366868
rect 137572 365498 137600 485862
rect 137652 466472 137704 466478
rect 137652 466414 137704 466420
rect 137560 365492 137612 365498
rect 137560 365434 137612 365440
rect 137664 358630 137692 466414
rect 137744 461032 137796 461038
rect 137744 460974 137796 460980
rect 137652 358624 137704 358630
rect 137652 358566 137704 358572
rect 137756 355978 137784 460974
rect 137744 355972 137796 355978
rect 137744 355914 137796 355920
rect 137284 339652 137336 339658
rect 137284 339594 137336 339600
rect 137296 292534 137324 339594
rect 137652 329996 137704 330002
rect 137652 329938 137704 329944
rect 137560 325916 137612 325922
rect 137560 325858 137612 325864
rect 137468 323196 137520 323202
rect 137468 323138 137520 323144
rect 137376 301028 137428 301034
rect 137376 300970 137428 300976
rect 137284 292528 137336 292534
rect 137284 292470 137336 292476
rect 137284 290488 137336 290494
rect 137284 290430 137336 290436
rect 137296 183530 137324 290430
rect 137388 195906 137416 300970
rect 137480 251122 137508 323138
rect 137572 256698 137600 325858
rect 137664 266354 137692 329938
rect 137652 266348 137704 266354
rect 137652 266290 137704 266296
rect 137560 256692 137612 256698
rect 137560 256634 137612 256640
rect 137468 251116 137520 251122
rect 137468 251058 137520 251064
rect 137376 195900 137428 195906
rect 137376 195842 137428 195848
rect 137284 183524 137336 183530
rect 137284 183466 137336 183472
rect 136732 104916 136784 104922
rect 136732 104858 136784 104864
rect 136744 97753 136772 104858
rect 136730 97744 136786 97753
rect 136730 97679 136786 97688
rect 137284 94512 137336 94518
rect 137284 94454 137336 94460
rect 137296 86902 137324 94454
rect 137284 86896 137336 86902
rect 137284 86838 137336 86844
rect 137376 85604 137428 85610
rect 137376 85546 137428 85552
rect 137284 74588 137336 74594
rect 137284 74530 137336 74536
rect 137296 56438 137324 74530
rect 137388 71670 137416 85546
rect 137376 71664 137428 71670
rect 137376 71606 137428 71612
rect 137376 68332 137428 68338
rect 137376 68274 137428 68280
rect 137284 56432 137336 56438
rect 137284 56374 137336 56380
rect 136640 52012 136692 52018
rect 136640 51954 136692 51960
rect 135996 51468 136048 51474
rect 135996 51410 136048 51416
rect 135904 51400 135956 51406
rect 135904 51342 135956 51348
rect 134708 51332 134760 51338
rect 134708 51274 134760 51280
rect 137388 50998 137416 68274
rect 135352 50992 135404 50998
rect 135350 50960 135352 50969
rect 137376 50992 137428 50998
rect 135404 50960 135406 50969
rect 137376 50934 137428 50940
rect 135350 50895 135406 50904
rect 138676 50114 138704 700334
rect 141424 670744 141476 670750
rect 141424 670686 141476 670692
rect 140044 590708 140096 590714
rect 140044 590650 140096 590656
rect 138756 581664 138808 581670
rect 138756 581606 138808 581612
rect 138768 404122 138796 581606
rect 138848 553444 138900 553450
rect 138848 553386 138900 553392
rect 138756 404116 138808 404122
rect 138756 404058 138808 404064
rect 138860 393174 138888 553386
rect 138940 531412 138992 531418
rect 138940 531354 138992 531360
rect 138848 393168 138900 393174
rect 138848 393110 138900 393116
rect 138952 383518 138980 531354
rect 139032 525904 139084 525910
rect 139032 525846 139084 525852
rect 138940 383512 138992 383518
rect 138940 383454 138992 383460
rect 139044 382090 139072 525846
rect 139124 512032 139176 512038
rect 139124 511974 139176 511980
rect 139032 382084 139084 382090
rect 139032 382026 139084 382032
rect 139136 378826 139164 511974
rect 139216 455456 139268 455462
rect 139216 455398 139268 455404
rect 139124 378820 139176 378826
rect 139124 378762 139176 378768
rect 139228 353054 139256 455398
rect 140056 408474 140084 590650
rect 140136 563100 140188 563106
rect 140136 563042 140188 563048
rect 140044 408468 140096 408474
rect 140044 408410 140096 408416
rect 140148 395894 140176 563042
rect 140228 560312 140280 560318
rect 140228 560254 140280 560260
rect 140136 395888 140188 395894
rect 140136 395830 140188 395836
rect 140240 395826 140268 560254
rect 140320 516180 140372 516186
rect 140320 516122 140372 516128
rect 140228 395820 140280 395826
rect 140228 395762 140280 395768
rect 140332 377942 140360 516122
rect 140412 502444 140464 502450
rect 140412 502386 140464 502392
rect 140320 377936 140372 377942
rect 140320 377878 140372 377884
rect 140424 372434 140452 502386
rect 140504 502376 140556 502382
rect 140504 502318 140556 502324
rect 140412 372428 140464 372434
rect 140412 372370 140464 372376
rect 140516 372366 140544 502318
rect 140596 485104 140648 485110
rect 140596 485046 140648 485052
rect 140504 372360 140556 372366
rect 140504 372302 140556 372308
rect 140608 368354 140636 485046
rect 140688 447160 140740 447166
rect 140688 447102 140740 447108
rect 140596 368348 140648 368354
rect 140596 368290 140648 368296
rect 139216 353048 139268 353054
rect 139216 352990 139268 352996
rect 140700 350470 140728 447102
rect 140688 350464 140740 350470
rect 140688 350406 140740 350412
rect 138756 349240 138808 349246
rect 138756 349182 138808 349188
rect 138768 314634 138796 349182
rect 140136 345092 140188 345098
rect 140136 345034 140188 345040
rect 139216 342372 139268 342378
rect 139216 342314 139268 342320
rect 139124 336932 139176 336938
rect 139124 336874 139176 336880
rect 139032 317620 139084 317626
rect 139032 317562 139084 317568
rect 138756 314628 138808 314634
rect 138756 314570 138808 314576
rect 138940 310684 138992 310690
rect 138940 310626 138992 310632
rect 138756 302456 138808 302462
rect 138756 302398 138808 302404
rect 138768 195974 138796 302398
rect 138848 296880 138900 296886
rect 138848 296822 138900 296828
rect 138860 200802 138888 296822
rect 138952 216646 138980 310626
rect 139044 236706 139072 317562
rect 139136 285598 139164 336874
rect 139228 296614 139256 342314
rect 140044 324964 140096 324970
rect 140044 324906 140096 324912
rect 139216 296608 139268 296614
rect 139216 296550 139268 296556
rect 139124 285592 139176 285598
rect 139124 285534 139176 285540
rect 139032 236700 139084 236706
rect 139032 236642 139084 236648
rect 138940 216640 138992 216646
rect 138940 216582 138992 216588
rect 138848 200796 138900 200802
rect 138848 200738 138900 200744
rect 138756 195968 138808 195974
rect 138756 195910 138808 195916
rect 139400 102196 139452 102202
rect 139400 102138 139452 102144
rect 138848 100768 138900 100774
rect 138848 100710 138900 100716
rect 138860 92478 138888 100710
rect 139412 96286 139440 102138
rect 139400 96280 139452 96286
rect 139400 96222 139452 96228
rect 138848 92472 138900 92478
rect 138848 92414 138900 92420
rect 138756 91112 138808 91118
rect 138756 91054 138808 91060
rect 138768 79762 138796 91054
rect 138848 81456 138900 81462
rect 138848 81398 138900 81404
rect 138756 79756 138808 79762
rect 138756 79698 138808 79704
rect 138756 66292 138808 66298
rect 138756 66234 138808 66240
rect 138664 50108 138716 50114
rect 138664 50050 138716 50056
rect 134614 48376 134670 48385
rect 134614 48311 134670 48320
rect 134524 47728 134576 47734
rect 134524 47670 134576 47676
rect 136546 47696 136602 47705
rect 133144 47592 133196 47598
rect 133144 47534 133196 47540
rect 133326 47560 133382 47569
rect 24124 25424 24176 25430
rect 24124 25366 24176 25372
rect 22742 24848 22798 24857
rect 22742 24783 22798 24792
rect 89720 24812 89772 24818
rect 89720 24754 89772 24760
rect 81440 24676 81492 24682
rect 81440 24618 81492 24624
rect 71780 24608 71832 24614
rect 71780 24550 71832 24556
rect 64880 24540 64932 24546
rect 64880 24482 64932 24488
rect 60740 24472 60792 24478
rect 60740 24414 60792 24420
rect 57980 24404 58032 24410
rect 57980 24346 58032 24352
rect 46940 24336 46992 24342
rect 46940 24278 46992 24284
rect 45560 24268 45612 24274
rect 45560 24210 45612 24216
rect 38660 24200 38712 24206
rect 18602 24168 18658 24177
rect 38660 24142 38712 24148
rect 18602 24103 18658 24112
rect 35900 24132 35952 24138
rect 13820 22840 13872 22846
rect 13820 22782 13872 22788
rect 9680 22772 9732 22778
rect 9680 22714 9732 22720
rect 4160 21412 4212 21418
rect 4160 21354 4212 21360
rect 1398 21312 1454 21321
rect 1398 21247 1454 21256
rect 572 3460 624 3466
rect 572 3402 624 3408
rect 584 480 612 3402
rect 542 -960 654 480
rect 1412 354 1440 21247
rect 3424 20664 3476 20670
rect 3424 20606 3476 20612
rect 3436 19417 3464 20606
rect 3422 19408 3478 19417
rect 3422 19343 3478 19352
rect 4172 16574 4200 21354
rect 6920 18624 6972 18630
rect 6920 18566 6972 18572
rect 6932 16574 6960 18566
rect 4172 16546 5304 16574
rect 6932 16546 7696 16574
rect 2872 15904 2924 15910
rect 2872 15846 2924 15852
rect 2884 480 2912 15846
rect 3606 11656 3662 11665
rect 3606 11591 3662 11600
rect 3424 6860 3476 6866
rect 3424 6802 3476 6808
rect 3436 6497 3464 6802
rect 3422 6488 3478 6497
rect 3422 6423 3478 6432
rect 1646 354 1758 480
rect 1412 326 1758 354
rect 1646 -960 1758 326
rect 2842 -960 2954 480
rect 3620 354 3648 11591
rect 5276 480 5304 16546
rect 6460 3664 6512 3670
rect 6460 3606 6512 3612
rect 6472 480 6500 3606
rect 7668 480 7696 16546
rect 8760 11756 8812 11762
rect 8760 11698 8812 11704
rect 8772 480 8800 11698
rect 4038 354 4150 480
rect 3620 326 4150 354
rect 4038 -960 4150 326
rect 5234 -960 5346 480
rect 6430 -960 6542 480
rect 7626 -960 7738 480
rect 8730 -960 8842 480
rect 9692 354 9720 22714
rect 11060 18692 11112 18698
rect 11060 18634 11112 18640
rect 11072 16574 11100 18634
rect 13832 16574 13860 22782
rect 15200 21480 15252 21486
rect 15200 21422 15252 21428
rect 15212 16574 15240 21422
rect 11072 16546 11928 16574
rect 13832 16546 14320 16574
rect 15212 16546 15976 16574
rect 11152 3732 11204 3738
rect 11152 3674 11204 3680
rect 11164 480 11192 3674
rect 9926 354 10038 480
rect 9692 326 10038 354
rect 9926 -960 10038 326
rect 11122 -960 11234 480
rect 11900 354 11928 16546
rect 13544 14476 13596 14482
rect 13544 14418 13596 14424
rect 13556 480 13584 14418
rect 12318 354 12430 480
rect 11900 326 12430 354
rect 12318 -960 12430 326
rect 13514 -960 13626 480
rect 14292 354 14320 16546
rect 15948 480 15976 16546
rect 18236 5024 18288 5030
rect 18236 4966 18288 4972
rect 17040 3528 17092 3534
rect 17040 3470 17092 3476
rect 17052 480 17080 3470
rect 18248 480 18276 4966
rect 18616 3534 18644 24103
rect 35900 24074 35952 24080
rect 31760 22908 31812 22914
rect 31760 22850 31812 22856
rect 19338 22672 19394 22681
rect 19338 22607 19394 22616
rect 19352 16574 19380 22607
rect 20718 18592 20774 18601
rect 20718 18527 20774 18536
rect 20732 16574 20760 18527
rect 31772 16574 31800 22850
rect 34520 19984 34572 19990
rect 34520 19926 34572 19932
rect 33140 17264 33192 17270
rect 33140 17206 33192 17212
rect 33152 16574 33180 17206
rect 19352 16546 20208 16574
rect 20732 16546 21864 16574
rect 31772 16546 31984 16574
rect 33152 16546 33640 16574
rect 18604 3528 18656 3534
rect 18604 3470 18656 3476
rect 19432 3528 19484 3534
rect 19432 3470 19484 3476
rect 19444 480 19472 3470
rect 14710 354 14822 480
rect 14292 326 14822 354
rect 14710 -960 14822 326
rect 15906 -960 16018 480
rect 17010 -960 17122 480
rect 18206 -960 18318 480
rect 19402 -960 19514 480
rect 20180 354 20208 16546
rect 21836 480 21864 16546
rect 28448 15972 28500 15978
rect 28448 15914 28500 15920
rect 26240 13116 26292 13122
rect 26240 13058 26292 13064
rect 23018 8936 23074 8945
rect 23018 8871 23074 8880
rect 23032 480 23060 8871
rect 25320 3868 25372 3874
rect 25320 3810 25372 3816
rect 24216 3596 24268 3602
rect 24216 3538 24268 3544
rect 24228 480 24256 3538
rect 25332 480 25360 3810
rect 20598 354 20710 480
rect 20180 326 20710 354
rect 20598 -960 20710 326
rect 21794 -960 21906 480
rect 22990 -960 23102 480
rect 24186 -960 24298 480
rect 25290 -960 25402 480
rect 26252 354 26280 13058
rect 27712 7608 27764 7614
rect 27712 7550 27764 7556
rect 27724 480 27752 7550
rect 26486 354 26598 480
rect 26252 326 26598 354
rect 26486 -960 26598 326
rect 27682 -960 27794 480
rect 28460 354 28488 15914
rect 30104 13184 30156 13190
rect 30104 13126 30156 13132
rect 30116 480 30144 13126
rect 31300 4888 31352 4894
rect 31300 4830 31352 4836
rect 31312 480 31340 4830
rect 28878 354 28990 480
rect 28460 326 28990 354
rect 28878 -960 28990 326
rect 30074 -960 30186 480
rect 31270 -960 31382 480
rect 31956 354 31984 16546
rect 33612 480 33640 16546
rect 32374 354 32486 480
rect 31956 326 32486 354
rect 32374 -960 32486 326
rect 33570 -960 33682 480
rect 34532 354 34560 19926
rect 35912 16574 35940 24074
rect 38672 16574 38700 24142
rect 45572 16574 45600 24210
rect 46952 16574 46980 24278
rect 53840 21616 53892 21622
rect 53840 21558 53892 21564
rect 49700 21548 49752 21554
rect 49700 21490 49752 21496
rect 49712 16574 49740 21490
rect 51080 17332 51132 17338
rect 51080 17274 51132 17280
rect 35912 16546 36032 16574
rect 38672 16546 39160 16574
rect 45572 16546 46704 16574
rect 46952 16546 47440 16574
rect 49712 16546 50200 16574
rect 36004 480 36032 16546
rect 36726 10296 36782 10305
rect 36726 10231 36782 10240
rect 34766 354 34878 480
rect 34532 326 34878 354
rect 34766 -960 34878 326
rect 35962 -960 36074 480
rect 36740 354 36768 10231
rect 38382 6216 38438 6225
rect 38382 6151 38438 6160
rect 38396 480 38424 6151
rect 37158 354 37270 480
rect 36740 326 37270 354
rect 37158 -960 37270 326
rect 38354 -960 38466 480
rect 39132 354 39160 16546
rect 41878 15872 41934 15881
rect 41878 15807 41934 15816
rect 40682 6352 40738 6361
rect 40682 6287 40738 6296
rect 40696 480 40724 6287
rect 41892 480 41920 15807
rect 45468 8968 45520 8974
rect 45468 8910 45520 8916
rect 44272 4956 44324 4962
rect 44272 4898 44324 4904
rect 43076 3800 43128 3806
rect 43076 3742 43128 3748
rect 43088 480 43116 3742
rect 44284 480 44312 4898
rect 45480 480 45508 8910
rect 46676 480 46704 16546
rect 39550 354 39662 480
rect 39132 326 39662 354
rect 39550 -960 39662 326
rect 40654 -960 40766 480
rect 41850 -960 41962 480
rect 43046 -960 43158 480
rect 44242 -960 44354 480
rect 45438 -960 45550 480
rect 46634 -960 46746 480
rect 47412 354 47440 16546
rect 48964 7676 49016 7682
rect 48964 7618 49016 7624
rect 48976 480 49004 7618
rect 50172 480 50200 16546
rect 47830 354 47942 480
rect 47412 326 47942 354
rect 47830 -960 47942 326
rect 48934 -960 49046 480
rect 50130 -960 50242 480
rect 51092 354 51120 17274
rect 53852 16574 53880 21558
rect 57992 16574 58020 24346
rect 53852 16546 54984 16574
rect 57992 16546 58480 16574
rect 53288 11824 53340 11830
rect 53288 11766 53340 11772
rect 52552 6180 52604 6186
rect 52552 6122 52604 6128
rect 52564 480 52592 6122
rect 51326 354 51438 480
rect 51092 326 51438 354
rect 51326 -960 51438 326
rect 52522 -960 52634 480
rect 53300 354 53328 11766
rect 54956 480 54984 16546
rect 56046 4856 56102 4865
rect 56046 4791 56102 4800
rect 56060 480 56088 4791
rect 57244 3936 57296 3942
rect 57244 3878 57296 3884
rect 57256 480 57284 3878
rect 58452 480 58480 16546
rect 59636 7744 59688 7750
rect 59636 7686 59688 7692
rect 59648 480 59676 7686
rect 60752 3398 60780 24414
rect 60832 17400 60884 17406
rect 60832 17342 60884 17348
rect 60740 3392 60792 3398
rect 60740 3334 60792 3340
rect 60844 480 60872 17342
rect 64892 16574 64920 24482
rect 67640 20052 67692 20058
rect 67640 19994 67692 20000
rect 64892 16546 65104 16574
rect 63224 13252 63276 13258
rect 63224 13194 63276 13200
rect 61660 3392 61712 3398
rect 61660 3334 61712 3340
rect 53718 354 53830 480
rect 53300 326 53830 354
rect 53718 -960 53830 326
rect 54914 -960 55026 480
rect 56018 -960 56130 480
rect 57214 -960 57326 480
rect 58410 -960 58522 480
rect 59606 -960 59718 480
rect 60802 -960 60914 480
rect 61672 354 61700 3334
rect 63236 480 63264 13194
rect 64328 7812 64380 7818
rect 64328 7754 64380 7760
rect 64340 480 64368 7754
rect 61998 354 62110 480
rect 61672 326 62110 354
rect 61998 -960 62110 326
rect 63194 -960 63306 480
rect 64298 -960 64410 480
rect 65076 354 65104 16546
rect 66720 6248 66772 6254
rect 66720 6190 66772 6196
rect 66732 480 66760 6190
rect 65494 354 65606 480
rect 65076 326 65606 354
rect 65494 -960 65606 326
rect 66690 -960 66802 480
rect 67652 354 67680 19994
rect 69020 18828 69072 18834
rect 69020 18770 69072 18776
rect 69032 6914 69060 18770
rect 69112 18760 69164 18766
rect 69112 18702 69164 18708
rect 69124 16574 69152 18702
rect 71792 16574 71820 24550
rect 78680 21684 78732 21690
rect 78680 21626 78732 21632
rect 75918 17232 75974 17241
rect 75918 17167 75974 17176
rect 69124 16546 69888 16574
rect 71792 16546 72648 16574
rect 69032 6886 69152 6914
rect 69124 480 69152 6886
rect 67886 354 67998 480
rect 67652 326 67998 354
rect 67886 -960 67998 326
rect 69082 -960 69194 480
rect 69860 354 69888 16546
rect 71504 9036 71556 9042
rect 71504 8978 71556 8984
rect 71516 480 71544 8978
rect 72620 480 72648 16546
rect 74998 13016 75054 13025
rect 74998 12951 75054 12960
rect 73802 4992 73858 5001
rect 73802 4927 73858 4936
rect 73816 480 73844 4927
rect 75012 480 75040 12951
rect 70278 354 70390 480
rect 69860 326 70390 354
rect 70278 -960 70390 326
rect 71474 -960 71586 480
rect 72578 -960 72690 480
rect 73774 -960 73886 480
rect 74970 -960 75082 480
rect 75932 354 75960 17167
rect 78692 16574 78720 21626
rect 81452 16574 81480 24618
rect 85580 22976 85632 22982
rect 85580 22918 85632 22924
rect 82820 20120 82872 20126
rect 82820 20062 82872 20068
rect 82832 16574 82860 20062
rect 85592 16574 85620 22918
rect 89732 16574 89760 24754
rect 95240 24744 95292 24750
rect 95240 24686 95292 24692
rect 93858 21448 93914 21457
rect 93858 21383 93914 21392
rect 93872 16574 93900 21383
rect 95252 16574 95280 24686
rect 107660 24064 107712 24070
rect 107660 24006 107712 24012
rect 102140 20188 102192 20194
rect 102140 20130 102192 20136
rect 78692 16546 79272 16574
rect 81452 16546 81664 16574
rect 82832 16546 83320 16574
rect 85592 16546 85712 16574
rect 89732 16546 89944 16574
rect 93872 16546 93992 16574
rect 95252 16546 95832 16574
rect 77298 14512 77354 14521
rect 77298 14447 77354 14456
rect 77312 3398 77340 14447
rect 77392 11892 77444 11898
rect 77392 11834 77444 11840
rect 77300 3392 77352 3398
rect 77300 3334 77352 3340
rect 77404 480 77432 11834
rect 78220 3392 78272 3398
rect 78220 3334 78272 3340
rect 76166 354 76278 480
rect 75932 326 76278 354
rect 76166 -960 76278 326
rect 77362 -960 77474 480
rect 78232 354 78260 3334
rect 78558 354 78670 480
rect 78232 326 78670 354
rect 79244 354 79272 16546
rect 80888 14544 80940 14550
rect 80888 14486 80940 14492
rect 80900 480 80928 14486
rect 79662 354 79774 480
rect 79244 326 79774 354
rect 78558 -960 78670 326
rect 79662 -960 79774 326
rect 80858 -960 80970 480
rect 81636 354 81664 16546
rect 83292 480 83320 16546
rect 84476 7880 84528 7886
rect 84476 7822 84528 7828
rect 84488 480 84516 7822
rect 85684 480 85712 16546
rect 87512 14612 87564 14618
rect 87512 14554 87564 14560
rect 86408 10328 86460 10334
rect 86408 10270 86460 10276
rect 82054 354 82166 480
rect 81636 326 82166 354
rect 82054 -960 82166 326
rect 83250 -960 83362 480
rect 84446 -960 84558 480
rect 85642 -960 85754 480
rect 86420 354 86448 10270
rect 86838 354 86950 480
rect 86420 326 86950 354
rect 87524 354 87552 14554
rect 89168 4004 89220 4010
rect 89168 3946 89220 3952
rect 89180 480 89208 3946
rect 87942 354 88054 480
rect 87524 326 88054 354
rect 86838 -960 86950 326
rect 87942 -960 88054 326
rect 89138 -960 89250 480
rect 89916 354 89944 16546
rect 91558 14648 91614 14657
rect 91558 14583 91614 14592
rect 91572 480 91600 14583
rect 92756 4072 92808 4078
rect 92756 4014 92808 4020
rect 92768 480 92796 4014
rect 93964 480 93992 16546
rect 94686 13152 94742 13161
rect 94686 13087 94742 13096
rect 90334 354 90446 480
rect 89916 326 90446 354
rect 90334 -960 90446 326
rect 91530 -960 91642 480
rect 92726 -960 92838 480
rect 93922 -960 94034 480
rect 94700 354 94728 13087
rect 95118 354 95230 480
rect 94700 326 95230 354
rect 95804 354 95832 16546
rect 98184 16040 98236 16046
rect 98184 15982 98236 15988
rect 97448 10396 97500 10402
rect 97448 10338 97500 10344
rect 97460 480 97488 10338
rect 96222 354 96334 480
rect 95804 326 96334 354
rect 95118 -960 95230 326
rect 96222 -960 96334 326
rect 97418 -960 97530 480
rect 98196 354 98224 15982
rect 99840 11960 99892 11966
rect 99840 11902 99892 11908
rect 99852 480 99880 11902
rect 100760 10464 100812 10470
rect 100760 10406 100812 10412
rect 98614 354 98726 480
rect 98196 326 98726 354
rect 98614 -960 98726 326
rect 99810 -960 99922 480
rect 100772 354 100800 10406
rect 102152 3398 102180 20130
rect 107672 16574 107700 24006
rect 120080 23996 120132 24002
rect 120080 23938 120132 23944
rect 110420 23928 110472 23934
rect 110420 23870 110472 23876
rect 110432 16574 110460 23870
rect 120092 16574 120120 23938
rect 121460 21752 121512 21758
rect 121460 21694 121512 21700
rect 121472 16574 121500 21694
rect 122840 20256 122892 20262
rect 122840 20198 122892 20204
rect 122852 16574 122880 20198
rect 131118 18864 131174 18873
rect 131118 18799 131174 18808
rect 129738 18728 129794 18737
rect 129738 18663 129794 18672
rect 126980 17536 127032 17542
rect 126980 17478 127032 17484
rect 125600 17468 125652 17474
rect 125600 17410 125652 17416
rect 107672 16546 108160 16574
rect 110432 16546 110552 16574
rect 120092 16546 120672 16574
rect 121472 16546 122328 16574
rect 122852 16546 123064 16574
rect 104072 16176 104124 16182
rect 104072 16118 104124 16124
rect 102232 16108 102284 16114
rect 102232 16050 102284 16056
rect 102140 3392 102192 3398
rect 102140 3334 102192 3340
rect 102244 480 102272 16050
rect 103336 3392 103388 3398
rect 103336 3334 103388 3340
rect 103348 480 103376 3334
rect 101006 354 101118 480
rect 100772 326 101118 354
rect 101006 -960 101118 326
rect 102202 -960 102314 480
rect 103306 -960 103418 480
rect 104084 354 104112 16118
rect 105728 6316 105780 6322
rect 105728 6258 105780 6264
rect 105740 480 105768 6258
rect 106924 3392 106976 3398
rect 106924 3334 106976 3340
rect 106936 480 106964 3334
rect 108132 480 108160 16546
rect 109314 9072 109370 9081
rect 109314 9007 109370 9016
rect 109328 480 109356 9007
rect 110524 480 110552 16546
rect 116400 16244 116452 16250
rect 116400 16186 116452 16192
rect 114008 14680 114060 14686
rect 114008 14622 114060 14628
rect 112810 9208 112866 9217
rect 112810 9143 112866 9152
rect 111614 5128 111670 5137
rect 111614 5063 111670 5072
rect 111628 480 111656 5063
rect 112824 480 112852 9143
rect 114020 480 114048 14622
rect 114744 13320 114796 13326
rect 114744 13262 114796 13268
rect 104502 354 104614 480
rect 104084 326 104614 354
rect 104502 -960 104614 326
rect 105698 -960 105810 480
rect 106894 -960 107006 480
rect 108090 -960 108202 480
rect 109286 -960 109398 480
rect 110482 -960 110594 480
rect 111586 -960 111698 480
rect 112782 -960 112894 480
rect 113978 -960 114090 480
rect 114756 354 114784 13262
rect 116412 480 116440 16186
rect 118792 10532 118844 10538
rect 118792 10474 118844 10480
rect 117596 3324 117648 3330
rect 117596 3266 117648 3272
rect 117608 480 117636 3266
rect 118804 480 118832 10474
rect 119896 9104 119948 9110
rect 119896 9046 119948 9052
rect 119908 480 119936 9046
rect 115174 354 115286 480
rect 114756 326 115286 354
rect 115174 -960 115286 326
rect 116370 -960 116482 480
rect 117566 -960 117678 480
rect 118762 -960 118874 480
rect 119866 -960 119978 480
rect 120644 354 120672 16546
rect 122300 480 122328 16546
rect 121062 354 121174 480
rect 120644 326 121174 354
rect 121062 -960 121174 326
rect 122258 -960 122370 480
rect 123036 354 123064 16546
rect 124680 4140 124732 4146
rect 124680 4082 124732 4088
rect 124692 480 124720 4082
rect 123454 354 123566 480
rect 123036 326 123566 354
rect 123454 -960 123566 326
rect 124650 -960 124762 480
rect 125612 354 125640 17410
rect 126992 480 127020 17478
rect 127070 17368 127126 17377
rect 127070 17303 127126 17312
rect 127084 16574 127112 17303
rect 129752 16574 129780 18663
rect 131132 16574 131160 18799
rect 127084 16546 128216 16574
rect 129752 16546 130608 16574
rect 131132 16546 131344 16574
rect 128188 480 128216 16546
rect 128912 12028 128964 12034
rect 128912 11970 128964 11976
rect 125846 354 125958 480
rect 125612 326 125958 354
rect 125846 -960 125958 326
rect 126950 -960 127062 480
rect 128146 -960 128258 480
rect 128924 354 128952 11970
rect 130580 480 130608 16546
rect 129342 354 129454 480
rect 128924 326 129454 354
rect 129342 -960 129454 326
rect 130538 -960 130650 480
rect 131316 354 131344 16546
rect 133156 4010 133184 47534
rect 133326 47495 133382 47504
rect 133340 26234 133368 47495
rect 133248 26206 133368 26234
rect 133144 4004 133196 4010
rect 133144 3946 133196 3952
rect 133248 3942 133276 26206
rect 133236 3936 133288 3942
rect 133236 3878 133288 3884
rect 134156 3936 134208 3942
rect 134156 3878 134208 3884
rect 132960 3120 133012 3126
rect 132960 3062 133012 3068
rect 132972 480 133000 3062
rect 134168 480 134196 3878
rect 134536 3738 134564 47670
rect 134616 47660 134668 47666
rect 136546 47631 136602 47640
rect 134616 47602 134668 47608
rect 134524 3732 134576 3738
rect 134524 3674 134576 3680
rect 134628 3398 134656 47602
rect 136560 47462 136588 47631
rect 136548 47456 136600 47462
rect 136548 47398 136600 47404
rect 138664 46504 138716 46510
rect 138664 46446 138716 46452
rect 134708 46368 134760 46374
rect 134708 46310 134760 46316
rect 137282 46336 137338 46345
rect 134616 3392 134668 3398
rect 134616 3334 134668 3340
rect 134720 3330 134748 46310
rect 137282 46271 137338 46280
rect 135996 46232 136048 46238
rect 134798 46200 134854 46209
rect 135996 46174 136048 46180
rect 134798 46135 134854 46144
rect 134812 4078 134840 46135
rect 135628 45552 135680 45558
rect 135626 45520 135628 45529
rect 135680 45520 135682 45529
rect 135626 45455 135682 45464
rect 135902 44840 135958 44849
rect 135902 44775 135958 44784
rect 135442 29472 135498 29481
rect 135442 29407 135498 29416
rect 135456 29102 135484 29407
rect 135444 29096 135496 29102
rect 135444 29038 135496 29044
rect 135260 26920 135312 26926
rect 135260 26862 135312 26868
rect 134800 4072 134852 4078
rect 134800 4014 134852 4020
rect 134708 3324 134760 3330
rect 134708 3266 134760 3272
rect 135272 480 135300 26862
rect 135916 3126 135944 44775
rect 136008 6866 136036 46174
rect 136548 43512 136600 43518
rect 136546 43480 136548 43489
rect 136600 43480 136602 43489
rect 136546 43415 136602 43424
rect 136640 43444 136692 43450
rect 136640 43386 136692 43392
rect 136088 41336 136140 41342
rect 136088 41278 136140 41284
rect 136100 40905 136128 41278
rect 136086 40896 136142 40905
rect 136086 40831 136142 40840
rect 136548 38072 136600 38078
rect 136548 38014 136600 38020
rect 136560 37913 136588 38014
rect 136546 37904 136602 37913
rect 136546 37839 136602 37848
rect 136548 35896 136600 35902
rect 136548 35838 136600 35844
rect 136560 35465 136588 35838
rect 136546 35456 136602 35465
rect 136546 35391 136602 35400
rect 136548 33040 136600 33046
rect 136546 33008 136548 33017
rect 136600 33008 136602 33017
rect 136546 32943 136602 32952
rect 136548 28280 136600 28286
rect 136548 28222 136600 28228
rect 136560 27577 136588 28222
rect 136546 27568 136602 27577
rect 136546 27503 136602 27512
rect 136652 16574 136680 43386
rect 136652 16546 137232 16574
rect 135996 6860 136048 6866
rect 135996 6802 136048 6808
rect 136456 3732 136508 3738
rect 136456 3674 136508 3680
rect 135904 3120 135956 3126
rect 135904 3062 135956 3068
rect 136468 480 136496 3674
rect 131734 354 131846 480
rect 131316 326 131846 354
rect 131734 -960 131846 326
rect 132930 -960 133042 480
rect 134126 -960 134238 480
rect 135230 -960 135342 480
rect 136426 -960 136538 480
rect 137204 354 137232 16546
rect 137296 3874 137324 46271
rect 138020 35216 138072 35222
rect 138020 35158 138072 35164
rect 138032 16574 138060 35158
rect 138032 16546 138612 16574
rect 137284 3868 137336 3874
rect 137284 3810 137336 3816
rect 138584 3482 138612 16546
rect 138676 3670 138704 46446
rect 138768 45558 138796 66234
rect 138860 66230 138888 81398
rect 138848 66224 138900 66230
rect 138848 66166 138900 66172
rect 138848 62144 138900 62150
rect 138848 62086 138900 62092
rect 138756 45552 138808 45558
rect 138756 45494 138808 45500
rect 138860 41342 138888 62086
rect 140056 49337 140084 324906
rect 140148 302190 140176 345034
rect 140596 334688 140648 334694
rect 140596 334630 140648 334636
rect 140504 332784 140556 332790
rect 140504 332726 140556 332732
rect 140412 328636 140464 328642
rect 140412 328578 140464 328584
rect 140320 303816 140372 303822
rect 140320 303758 140372 303764
rect 140136 302184 140188 302190
rect 140136 302126 140188 302132
rect 140228 301096 140280 301102
rect 140228 301038 140280 301044
rect 140136 294228 140188 294234
rect 140136 294170 140188 294176
rect 140148 184210 140176 294170
rect 140240 193118 140268 301038
rect 140332 200054 140360 303758
rect 140424 263498 140452 328578
rect 140516 274650 140544 332726
rect 140608 285666 140636 334630
rect 140596 285660 140648 285666
rect 140596 285602 140648 285608
rect 140504 274644 140556 274650
rect 140504 274586 140556 274592
rect 140412 263492 140464 263498
rect 140412 263434 140464 263440
rect 140320 200048 140372 200054
rect 140320 199990 140372 199996
rect 140228 193112 140280 193118
rect 140228 193054 140280 193060
rect 140136 184204 140188 184210
rect 140136 184146 140188 184152
rect 140136 92540 140188 92546
rect 140136 92482 140188 92488
rect 140148 82278 140176 92482
rect 140136 82272 140188 82278
rect 140136 82214 140188 82220
rect 140228 80096 140280 80102
rect 140228 80038 140280 80044
rect 140136 64932 140188 64938
rect 140136 64874 140188 64880
rect 140042 49328 140098 49337
rect 140042 49263 140098 49272
rect 139400 44872 139452 44878
rect 139400 44814 139452 44820
rect 138848 41336 138900 41342
rect 138848 41278 138900 41284
rect 139412 16574 139440 44814
rect 140148 43518 140176 64874
rect 140240 64190 140268 80038
rect 140228 64184 140280 64190
rect 140228 64126 140280 64132
rect 141436 50250 141464 670686
rect 141516 575544 141568 575550
rect 141516 575486 141568 575492
rect 141528 401538 141556 575486
rect 141608 567248 141660 567254
rect 141608 567190 141660 567196
rect 141516 401532 141568 401538
rect 141516 401474 141568 401480
rect 141620 398750 141648 567190
rect 141700 510672 141752 510678
rect 141700 510614 141752 510620
rect 141608 398744 141660 398750
rect 141608 398686 141660 398692
rect 141712 375222 141740 510614
rect 141792 507884 141844 507890
rect 141792 507826 141844 507832
rect 141700 375216 141752 375222
rect 141700 375158 141752 375164
rect 141804 373794 141832 507826
rect 141884 498840 141936 498846
rect 141884 498782 141936 498788
rect 141792 373788 141844 373794
rect 141792 373730 141844 373736
rect 141896 370938 141924 498782
rect 141976 470688 142028 470694
rect 141976 470630 142028 470636
rect 141884 370932 141936 370938
rect 141884 370874 141936 370880
rect 141988 359990 142016 470630
rect 142068 454096 142120 454102
rect 142068 454038 142120 454044
rect 141976 359984 142028 359990
rect 141976 359926 142028 359932
rect 142080 352986 142108 454038
rect 142068 352980 142120 352986
rect 142068 352922 142120 352928
rect 141516 345228 141568 345234
rect 141516 345170 141568 345176
rect 141528 304978 141556 345170
rect 141792 339720 141844 339726
rect 141792 339662 141844 339668
rect 141700 307964 141752 307970
rect 141700 307906 141752 307912
rect 141516 304972 141568 304978
rect 141516 304914 141568 304920
rect 141608 302932 141660 302938
rect 141608 302874 141660 302880
rect 141516 299668 141568 299674
rect 141516 299610 141568 299616
rect 141528 188970 141556 299610
rect 141620 200122 141648 302874
rect 141712 211138 141740 307906
rect 141804 289814 141832 339662
rect 141792 289808 141844 289814
rect 141792 289750 141844 289756
rect 141700 211132 141752 211138
rect 141700 211074 141752 211080
rect 141608 200116 141660 200122
rect 141608 200058 141660 200064
rect 141516 188964 141568 188970
rect 141516 188906 141568 188912
rect 142160 95260 142212 95266
rect 142160 95202 142212 95208
rect 141608 89752 141660 89758
rect 141608 89694 141660 89700
rect 141620 77110 141648 89694
rect 142172 87378 142200 95202
rect 142160 87372 142212 87378
rect 142160 87314 142212 87320
rect 141608 77104 141660 77110
rect 141608 77046 141660 77052
rect 141516 75948 141568 75954
rect 141516 75890 141568 75896
rect 141528 59022 141556 75890
rect 141516 59016 141568 59022
rect 141516 58958 141568 58964
rect 141516 56636 141568 56642
rect 141516 56578 141568 56584
rect 141424 50244 141476 50250
rect 141424 50186 141476 50192
rect 140136 43512 140188 43518
rect 140136 43454 140188 43460
rect 140780 37936 140832 37942
rect 140780 37878 140832 37884
rect 140792 16574 140820 37878
rect 141528 33046 141556 56578
rect 142816 52834 142844 700538
rect 151084 700528 151136 700534
rect 151084 700470 151136 700476
rect 148324 700460 148376 700466
rect 148324 700402 148376 700408
rect 144184 656940 144236 656946
rect 144184 656882 144236 656888
rect 142896 589348 142948 589354
rect 142896 589290 142948 589296
rect 142908 406910 142936 589290
rect 142988 572756 143040 572762
rect 142988 572698 143040 572704
rect 142896 406904 142948 406910
rect 142896 406846 142948 406852
rect 143000 401470 143028 572698
rect 143080 548548 143132 548554
rect 143080 548490 143132 548496
rect 142988 401464 143040 401470
rect 142988 401406 143040 401412
rect 143092 393106 143120 548490
rect 143172 534132 143224 534138
rect 143172 534074 143224 534080
rect 143080 393100 143132 393106
rect 143080 393042 143132 393048
rect 143184 384878 143212 534074
rect 143264 523048 143316 523054
rect 143264 522990 143316 522996
rect 143172 384872 143224 384878
rect 143172 384814 143224 384820
rect 143276 380594 143304 522990
rect 143356 509312 143408 509318
rect 143356 509254 143408 509260
rect 143264 380588 143316 380594
rect 143264 380530 143316 380536
rect 143368 376038 143396 509254
rect 143448 477556 143500 477562
rect 143448 477498 143500 477504
rect 143356 376032 143408 376038
rect 143356 375974 143408 375980
rect 143460 362778 143488 477498
rect 143448 362772 143500 362778
rect 143448 362714 143500 362720
rect 142988 346656 143040 346662
rect 142988 346598 143040 346604
rect 142896 322312 142948 322318
rect 142896 322254 142948 322260
rect 142804 52828 142856 52834
rect 142804 52770 142856 52776
rect 142908 48521 142936 322254
rect 143000 307766 143028 346598
rect 143356 337000 143408 337006
rect 143356 336942 143408 336948
rect 143264 327344 143316 327350
rect 143264 327286 143316 327292
rect 143172 320408 143224 320414
rect 143172 320350 143224 320356
rect 142988 307760 143040 307766
rect 142988 307702 143040 307708
rect 143080 306604 143132 306610
rect 143080 306546 143132 306552
rect 142988 299736 143040 299742
rect 142988 299678 143040 299684
rect 143000 190466 143028 299678
rect 143092 206990 143120 306546
rect 143184 242214 143212 320350
rect 143276 258058 143304 327286
rect 143368 284238 143396 336942
rect 143356 284232 143408 284238
rect 143356 284174 143408 284180
rect 143264 258052 143316 258058
rect 143264 257994 143316 258000
rect 143172 242208 143224 242214
rect 143172 242150 143224 242156
rect 143080 206984 143132 206990
rect 143080 206926 143132 206932
rect 142988 190460 143040 190466
rect 142988 190402 143040 190408
rect 143080 69080 143132 69086
rect 143080 69022 143132 69028
rect 142988 55276 143040 55282
rect 142988 55218 143040 55224
rect 142894 48512 142950 48521
rect 142894 48447 142950 48456
rect 141516 33040 141568 33046
rect 141516 32982 141568 32988
rect 143000 29102 143028 55218
rect 143092 47462 143120 69022
rect 144196 50318 144224 656882
rect 146944 618316 146996 618322
rect 146944 618258 146996 618264
rect 144276 562352 144328 562358
rect 144276 562294 144328 562300
rect 144288 398682 144316 562294
rect 144368 543788 144420 543794
rect 144368 543730 144420 543736
rect 144276 398676 144328 398682
rect 144276 398618 144328 398624
rect 144380 388958 144408 543730
rect 145564 534744 145616 534750
rect 145564 534686 145616 534692
rect 144460 525836 144512 525842
rect 144460 525778 144512 525784
rect 144368 388952 144420 388958
rect 144368 388894 144420 388900
rect 144472 382022 144500 525778
rect 144552 517540 144604 517546
rect 144552 517482 144604 517488
rect 144460 382016 144512 382022
rect 144460 381958 144512 381964
rect 144564 377874 144592 517482
rect 144644 487212 144696 487218
rect 144644 487154 144696 487160
rect 144552 377868 144604 377874
rect 144552 377810 144604 377816
rect 144656 366858 144684 487154
rect 144736 460964 144788 460970
rect 144736 460906 144788 460912
rect 144644 366852 144696 366858
rect 144644 366794 144696 366800
rect 144748 355910 144776 460906
rect 145576 387598 145604 534686
rect 145748 519580 145800 519586
rect 145748 519522 145800 519528
rect 145656 513392 145708 513398
rect 145656 513334 145708 513340
rect 145564 387592 145616 387598
rect 145564 387534 145616 387540
rect 145668 376514 145696 513334
rect 145760 390318 145788 519522
rect 145840 478916 145892 478922
rect 145840 478858 145892 478864
rect 145748 390312 145800 390318
rect 145748 390254 145800 390260
rect 145656 376508 145708 376514
rect 145656 376450 145708 376456
rect 145852 362710 145880 478858
rect 145932 448588 145984 448594
rect 145932 448530 145984 448536
rect 145840 362704 145892 362710
rect 145840 362646 145892 362652
rect 144736 355904 144788 355910
rect 144736 355846 144788 355852
rect 145944 351762 145972 448530
rect 145932 351756 145984 351762
rect 145932 351698 145984 351704
rect 144552 342440 144604 342446
rect 144552 342382 144604 342388
rect 144460 320476 144512 320482
rect 144460 320418 144512 320424
rect 144368 309460 144420 309466
rect 144368 309402 144420 309408
rect 144276 298240 144328 298246
rect 144276 298182 144328 298188
rect 144288 187678 144316 298182
rect 144380 215286 144408 309402
rect 144472 243574 144500 320418
rect 144564 298110 144592 342382
rect 144736 338292 144788 338298
rect 144736 338234 144788 338240
rect 144644 330064 144696 330070
rect 144644 330006 144696 330012
rect 144552 298104 144604 298110
rect 144552 298046 144604 298052
rect 144552 291848 144604 291854
rect 144552 291790 144604 291796
rect 144460 243568 144512 243574
rect 144460 243510 144512 243516
rect 144564 224942 144592 291790
rect 144656 264858 144684 330006
rect 144748 288386 144776 338234
rect 145932 335572 145984 335578
rect 145932 335514 145984 335520
rect 145840 332852 145892 332858
rect 145840 332794 145892 332800
rect 145656 317688 145708 317694
rect 145656 317630 145708 317636
rect 145564 295656 145616 295662
rect 145564 295598 145616 295604
rect 144736 288380 144788 288386
rect 144736 288322 144788 288328
rect 144644 264852 144696 264858
rect 144644 264794 144696 264800
rect 144552 224936 144604 224942
rect 144552 224878 144604 224884
rect 144368 215280 144420 215286
rect 144368 215222 144420 215228
rect 144276 187672 144328 187678
rect 144276 187614 144328 187620
rect 145576 179314 145604 295598
rect 145668 235278 145696 317630
rect 145748 310752 145800 310758
rect 145748 310694 145800 310700
rect 145656 235272 145708 235278
rect 145656 235214 145708 235220
rect 145760 232558 145788 310694
rect 145852 271794 145880 332794
rect 145944 280158 145972 335514
rect 145932 280152 145984 280158
rect 145932 280094 145984 280100
rect 145840 271788 145892 271794
rect 145840 271730 145892 271736
rect 145748 232552 145800 232558
rect 145748 232494 145800 232500
rect 145564 179308 145616 179314
rect 145564 179250 145616 179256
rect 144276 87032 144328 87038
rect 144276 86974 144328 86980
rect 144288 73778 144316 86974
rect 144276 73772 144328 73778
rect 144276 73714 144328 73720
rect 144276 60784 144328 60790
rect 144276 60726 144328 60732
rect 144184 50312 144236 50318
rect 144184 50254 144236 50260
rect 143080 47456 143132 47462
rect 143080 47398 143132 47404
rect 143540 46300 143592 46306
rect 143540 46242 143592 46248
rect 142988 29096 143040 29102
rect 142988 29038 143040 29044
rect 139412 16546 139624 16574
rect 140792 16546 141280 16574
rect 138664 3664 138716 3670
rect 138664 3606 138716 3612
rect 138584 3454 138888 3482
rect 138860 480 138888 3454
rect 137622 354 137734 480
rect 137204 326 137734 354
rect 137622 -960 137734 326
rect 138818 -960 138930 480
rect 139596 354 139624 16546
rect 141252 480 141280 16546
rect 143552 11694 143580 46242
rect 143632 44940 143684 44946
rect 143632 44882 143684 44888
rect 143540 11688 143592 11694
rect 143540 11630 143592 11636
rect 143644 6914 143672 44882
rect 144288 38078 144316 60726
rect 146956 48006 146984 618258
rect 147036 556232 147088 556238
rect 147036 556174 147088 556180
rect 147048 394466 147076 556174
rect 147128 532772 147180 532778
rect 147128 532714 147180 532720
rect 147036 394460 147088 394466
rect 147036 394402 147088 394408
rect 147140 384810 147168 532714
rect 147220 524476 147272 524482
rect 147220 524418 147272 524424
rect 147232 387122 147260 524418
rect 147312 512644 147364 512650
rect 147312 512586 147364 512592
rect 147220 387116 147272 387122
rect 147220 387058 147272 387064
rect 147128 384804 147180 384810
rect 147128 384746 147180 384752
rect 147324 379302 147352 512586
rect 147404 505776 147456 505782
rect 147404 505718 147456 505724
rect 147312 379296 147364 379302
rect 147312 379238 147364 379244
rect 147416 373726 147444 505718
rect 147496 470620 147548 470626
rect 147496 470562 147548 470568
rect 147404 373720 147456 373726
rect 147404 373662 147456 373668
rect 147508 359922 147536 470562
rect 147496 359916 147548 359922
rect 147496 359858 147548 359864
rect 147496 339788 147548 339794
rect 147496 339730 147548 339736
rect 147404 330540 147456 330546
rect 147404 330482 147456 330488
rect 147312 321836 147364 321842
rect 147312 321778 147364 321784
rect 147220 316260 147272 316266
rect 147220 316202 147272 316208
rect 147128 313608 147180 313614
rect 147128 313550 147180 313556
rect 147036 297424 147088 297430
rect 147036 297366 147088 297372
rect 147048 186318 147076 297366
rect 147140 223582 147168 313550
rect 147232 233918 147260 316202
rect 147324 245614 147352 321778
rect 147416 271862 147444 330482
rect 147508 291174 147536 339730
rect 147496 291168 147548 291174
rect 147496 291110 147548 291116
rect 147404 271856 147456 271862
rect 147404 271798 147456 271804
rect 147312 245608 147364 245614
rect 147312 245550 147364 245556
rect 147220 233912 147272 233918
rect 147220 233854 147272 233860
rect 147128 223576 147180 223582
rect 147128 223518 147180 223524
rect 147036 186312 147088 186318
rect 147036 186254 147088 186260
rect 147036 99408 147088 99414
rect 147036 99350 147088 99356
rect 147048 89690 147076 99350
rect 147036 89684 147088 89690
rect 147036 89626 147088 89632
rect 147036 77308 147088 77314
rect 147036 77250 147088 77256
rect 147048 62082 147076 77250
rect 147036 62076 147088 62082
rect 147036 62018 147088 62024
rect 147036 59424 147088 59430
rect 147036 59366 147088 59372
rect 146944 48000 146996 48006
rect 146944 47942 146996 47948
rect 146298 44976 146354 44985
rect 146298 44911 146354 44920
rect 144918 43480 144974 43489
rect 144918 43415 144974 43424
rect 144276 38072 144328 38078
rect 144276 38014 144328 38020
rect 144932 16574 144960 43415
rect 146312 16574 146340 44911
rect 147048 35902 147076 59366
rect 148336 50726 148364 700402
rect 148416 556844 148468 556850
rect 148416 556786 148468 556792
rect 148428 395758 148456 556786
rect 149704 552084 149756 552090
rect 149704 552026 149756 552032
rect 148508 535560 148560 535566
rect 148508 535502 148560 535508
rect 148416 395752 148468 395758
rect 148416 395694 148468 395700
rect 148520 386238 148548 535502
rect 148600 531344 148652 531350
rect 148600 531286 148652 531292
rect 148508 386232 148560 386238
rect 148508 386174 148560 386180
rect 148612 384742 148640 531286
rect 148692 501016 148744 501022
rect 148692 500958 148744 500964
rect 148600 384736 148652 384742
rect 148600 384678 148652 384684
rect 148704 372298 148732 500958
rect 148784 494080 148836 494086
rect 148784 494022 148836 494028
rect 148692 372292 148744 372298
rect 148692 372234 148744 372240
rect 148796 369578 148824 494022
rect 148876 451308 148928 451314
rect 148876 451250 148928 451256
rect 148784 369572 148836 369578
rect 148784 369514 148836 369520
rect 148888 351694 148916 451250
rect 149716 391746 149744 552026
rect 149796 541680 149848 541686
rect 149796 541622 149848 541628
rect 149808 398614 149836 541622
rect 149888 520940 149940 520946
rect 149888 520882 149940 520888
rect 149796 398608 149848 398614
rect 149796 398550 149848 398556
rect 149704 391740 149756 391746
rect 149704 391682 149756 391688
rect 149900 383450 149928 520882
rect 149980 463752 150032 463758
rect 149980 463694 150032 463700
rect 149888 383444 149940 383450
rect 149888 383386 149940 383392
rect 149992 357202 150020 463694
rect 150072 459604 150124 459610
rect 150072 459546 150124 459552
rect 150084 367878 150112 459546
rect 150072 367872 150124 367878
rect 150072 367814 150124 367820
rect 149980 357196 150032 357202
rect 149980 357138 150032 357144
rect 148876 351688 148928 351694
rect 148876 351630 148928 351636
rect 148876 338360 148928 338366
rect 148876 338302 148928 338308
rect 148784 334076 148836 334082
rect 148784 334018 148836 334024
rect 148692 319048 148744 319054
rect 148692 318990 148744 318996
rect 148600 317756 148652 317762
rect 148600 317698 148652 317704
rect 148508 306672 148560 306678
rect 148508 306614 148560 306620
rect 148416 298376 148468 298382
rect 148416 298318 148468 298324
rect 148428 189038 148456 298318
rect 148520 209098 148548 306614
rect 148612 234598 148640 317698
rect 148704 240106 148732 318990
rect 148796 277302 148824 334018
rect 148888 287026 148916 338302
rect 150072 331492 150124 331498
rect 150072 331434 150124 331440
rect 149980 328704 150032 328710
rect 149980 328646 150032 328652
rect 149888 324352 149940 324358
rect 149888 324294 149940 324300
rect 149796 308032 149848 308038
rect 149796 307974 149848 307980
rect 149704 298308 149756 298314
rect 149704 298250 149756 298256
rect 148876 287020 148928 287026
rect 148876 286962 148928 286968
rect 148784 277296 148836 277302
rect 148784 277238 148836 277244
rect 148692 240100 148744 240106
rect 148692 240042 148744 240048
rect 148600 234592 148652 234598
rect 148600 234534 148652 234540
rect 148508 209092 148560 209098
rect 148508 209034 148560 209040
rect 149716 193866 149744 298250
rect 149808 217326 149836 307974
rect 149900 251190 149928 324294
rect 149992 262206 150020 328646
rect 150084 270434 150112 331434
rect 150072 270428 150124 270434
rect 150072 270370 150124 270376
rect 149980 262200 150032 262206
rect 149980 262142 150032 262148
rect 149888 251184 149940 251190
rect 149888 251126 149940 251132
rect 149796 217320 149848 217326
rect 149796 217262 149848 217268
rect 149704 193860 149756 193866
rect 149704 193802 149756 193808
rect 148416 189032 148468 189038
rect 148416 188974 148468 188980
rect 149060 120148 149112 120154
rect 149060 120090 149112 120096
rect 149072 118658 149100 120090
rect 149060 118652 149112 118658
rect 149060 118594 149112 118600
rect 149060 117360 149112 117366
rect 149060 117302 149112 117308
rect 149072 115938 149100 117302
rect 149060 115932 149112 115938
rect 149060 115874 149112 115880
rect 148416 52488 148468 52494
rect 148416 52430 148468 52436
rect 148324 50720 148376 50726
rect 148324 50662 148376 50668
rect 147678 37904 147734 37913
rect 147678 37839 147734 37848
rect 147036 35896 147088 35902
rect 147036 35838 147088 35844
rect 147692 16574 147720 37839
rect 148428 28286 148456 52430
rect 151096 51542 151124 700470
rect 152556 576904 152608 576910
rect 152556 576846 152608 576852
rect 151176 554804 151228 554810
rect 151176 554746 151228 554752
rect 151188 393310 151216 554746
rect 151268 538280 151320 538286
rect 151268 538222 151320 538228
rect 151176 393304 151228 393310
rect 151176 393246 151228 393252
rect 151280 387802 151308 538222
rect 151360 535492 151412 535498
rect 151360 535434 151412 535440
rect 151268 387796 151320 387802
rect 151268 387738 151320 387744
rect 151372 386374 151400 535434
rect 151452 492720 151504 492726
rect 151452 492662 151504 492668
rect 151360 386368 151412 386374
rect 151360 386310 151412 386316
rect 151464 368490 151492 492662
rect 151544 485852 151596 485858
rect 151544 485794 151596 485800
rect 151452 368484 151504 368490
rect 151452 368426 151504 368432
rect 151556 365702 151584 485794
rect 151636 465112 151688 465118
rect 151636 465054 151688 465060
rect 151544 365696 151596 365702
rect 151544 365638 151596 365644
rect 151648 357406 151676 465054
rect 152464 409896 152516 409902
rect 152464 409838 152516 409844
rect 151636 357400 151688 357406
rect 151636 357342 151688 357348
rect 151544 336796 151596 336802
rect 151544 336738 151596 336744
rect 151452 335368 151504 335374
rect 151452 335310 151504 335316
rect 151360 325712 151412 325718
rect 151360 325654 151412 325660
rect 151268 310548 151320 310554
rect 151268 310490 151320 310496
rect 151176 294296 151228 294302
rect 151176 294238 151228 294244
rect 151188 176662 151216 294238
rect 151280 218754 151308 310490
rect 151372 255270 151400 325654
rect 151464 278662 151492 335310
rect 151556 284306 151584 336738
rect 151636 297220 151688 297226
rect 151636 297162 151688 297168
rect 151544 284300 151596 284306
rect 151544 284242 151596 284248
rect 151452 278656 151504 278662
rect 151452 278598 151504 278604
rect 151648 263566 151676 297162
rect 151636 263560 151688 263566
rect 151636 263502 151688 263508
rect 151360 255264 151412 255270
rect 151360 255206 151412 255212
rect 151268 218748 151320 218754
rect 151268 218690 151320 218696
rect 151176 176656 151228 176662
rect 151176 176598 151228 176604
rect 151268 133884 151320 133890
rect 151268 133826 151320 133832
rect 151176 133816 151228 133822
rect 151176 133758 151228 133764
rect 151084 51536 151136 51542
rect 151084 51478 151136 51484
rect 151188 46646 151216 133758
rect 151280 46782 151308 133826
rect 151360 133748 151412 133754
rect 151360 133690 151412 133696
rect 151372 50658 151400 133690
rect 151452 133408 151504 133414
rect 151452 133350 151504 133356
rect 151464 51610 151492 133350
rect 151636 84244 151688 84250
rect 151636 84186 151688 84192
rect 151648 72486 151676 84186
rect 151636 72480 151688 72486
rect 151636 72422 151688 72428
rect 151544 71800 151596 71806
rect 151544 71742 151596 71748
rect 151556 53786 151584 71742
rect 151544 53780 151596 53786
rect 151544 53722 151596 53728
rect 151452 51604 151504 51610
rect 151452 51546 151504 51552
rect 151360 50652 151412 50658
rect 151360 50594 151412 50600
rect 152476 47530 152504 409838
rect 152568 402490 152596 576846
rect 152648 574116 152700 574122
rect 152648 574058 152700 574064
rect 152556 402484 152608 402490
rect 152556 402426 152608 402432
rect 152660 401606 152688 574058
rect 152740 568608 152792 568614
rect 152740 568550 152792 568556
rect 152648 401600 152700 401606
rect 152648 401542 152700 401548
rect 152752 398818 152780 568550
rect 152832 546508 152884 546514
rect 152832 546450 152884 546456
rect 152740 398812 152792 398818
rect 152740 398754 152792 398760
rect 152844 390522 152872 546450
rect 152924 467900 152976 467906
rect 152924 467842 152976 467848
rect 152832 390516 152884 390522
rect 152832 390458 152884 390464
rect 152936 358766 152964 467842
rect 153016 462392 153068 462398
rect 153016 462334 153068 462340
rect 152924 358760 152976 358766
rect 152924 358702 152976 358708
rect 153028 356046 153056 462334
rect 153016 356040 153068 356046
rect 153016 355982 153068 355988
rect 153016 334008 153068 334014
rect 153016 333950 153068 333956
rect 152924 328772 152976 328778
rect 152924 328714 152976 328720
rect 152556 322244 152608 322250
rect 152556 322186 152608 322192
rect 152568 49201 152596 322186
rect 152832 316396 152884 316402
rect 152832 316338 152884 316344
rect 152740 311908 152792 311914
rect 152740 311850 152792 311856
rect 152648 303680 152700 303686
rect 152648 303622 152700 303628
rect 152660 207670 152688 303622
rect 152752 220114 152780 311850
rect 152844 246362 152872 316338
rect 152936 264926 152964 328714
rect 153028 276010 153056 333950
rect 153016 276004 153068 276010
rect 153016 275946 153068 275952
rect 152924 264920 152976 264926
rect 152924 264862 152976 264868
rect 152832 246356 152884 246362
rect 152832 246298 152884 246304
rect 152740 220108 152792 220114
rect 152740 220050 152792 220056
rect 152648 207664 152700 207670
rect 152648 207606 152700 207612
rect 153212 51746 153240 702406
rect 157984 700324 158036 700330
rect 157984 700266 158036 700272
rect 153844 549296 153896 549302
rect 153844 549238 153896 549244
rect 153856 390833 153884 549238
rect 155224 543040 155276 543046
rect 155224 542982 155276 542988
rect 153936 529984 153988 529990
rect 153936 529926 153988 529932
rect 153842 390824 153898 390833
rect 153842 390759 153898 390768
rect 153948 382945 153976 529926
rect 154028 518220 154080 518226
rect 154028 518162 154080 518168
rect 153934 382936 153990 382945
rect 153934 382871 153990 382880
rect 154040 378593 154068 518162
rect 154120 469260 154172 469266
rect 154120 469202 154172 469208
rect 154026 378584 154082 378593
rect 154026 378519 154082 378528
rect 154132 375358 154160 469202
rect 154672 409148 154724 409154
rect 154672 409090 154724 409096
rect 154580 406904 154632 406910
rect 154578 406872 154580 406881
rect 154632 406872 154634 406881
rect 154578 406807 154634 406816
rect 154684 405793 154712 409090
rect 154948 408468 155000 408474
rect 154948 408410 155000 408416
rect 154960 407425 154988 408410
rect 154946 407416 155002 407425
rect 154946 407351 155002 407360
rect 154856 407108 154908 407114
rect 154856 407050 154908 407056
rect 154764 407040 154816 407046
rect 154764 406982 154816 406988
rect 154776 406065 154804 406982
rect 154868 406337 154896 407050
rect 154948 406972 155000 406978
rect 154948 406914 155000 406920
rect 154960 406609 154988 406914
rect 154946 406600 155002 406609
rect 154946 406535 155002 406544
rect 154854 406328 154910 406337
rect 154854 406263 154910 406272
rect 154762 406056 154818 406065
rect 154762 405991 154818 406000
rect 154670 405784 154726 405793
rect 154670 405719 154726 405728
rect 154764 405680 154816 405686
rect 154764 405622 154816 405628
rect 154578 405512 154634 405521
rect 154578 405447 154580 405456
rect 154632 405447 154634 405456
rect 154580 405418 154632 405424
rect 154776 405249 154804 405622
rect 154856 405612 154908 405618
rect 154856 405554 154908 405560
rect 155040 405612 155092 405618
rect 155040 405554 155092 405560
rect 154762 405240 154818 405249
rect 154762 405175 154818 405184
rect 154868 404705 154896 405554
rect 154948 405544 155000 405550
rect 154948 405486 155000 405492
rect 154960 404977 154988 405486
rect 154946 404968 155002 404977
rect 154946 404903 155002 404912
rect 154854 404696 154910 404705
rect 154854 404631 154910 404640
rect 154672 404320 154724 404326
rect 154672 404262 154724 404268
rect 154684 404161 154712 404262
rect 154948 404252 155000 404258
rect 154948 404194 155000 404200
rect 154856 404184 154908 404190
rect 154670 404152 154726 404161
rect 154856 404126 154908 404132
rect 154670 404087 154726 404096
rect 154764 404116 154816 404122
rect 154764 404058 154816 404064
rect 154776 403889 154804 404058
rect 154762 403880 154818 403889
rect 154762 403815 154818 403824
rect 154868 403345 154896 404126
rect 154960 403617 154988 404194
rect 154946 403608 155002 403617
rect 154946 403543 155002 403552
rect 154854 403336 154910 403345
rect 154854 403271 154910 403280
rect 155052 402974 155080 405554
rect 155236 403073 155264 542982
rect 155316 529236 155368 529242
rect 155316 529178 155368 529184
rect 155328 405618 155356 529178
rect 155500 504416 155552 504422
rect 155500 504358 155552 504364
rect 155408 497480 155460 497486
rect 155408 497422 155460 497428
rect 155316 405612 155368 405618
rect 155316 405554 155368 405560
rect 155222 403064 155278 403073
rect 155222 402999 155278 403008
rect 155052 402946 155172 402974
rect 154764 402892 154816 402898
rect 154764 402834 154816 402840
rect 154670 402792 154726 402801
rect 154670 402727 154672 402736
rect 154724 402727 154726 402736
rect 154672 402698 154724 402704
rect 154776 402257 154804 402834
rect 154856 402824 154908 402830
rect 154856 402766 154908 402772
rect 154868 402529 154896 402766
rect 154948 402688 155000 402694
rect 154948 402630 155000 402636
rect 154854 402520 154910 402529
rect 154854 402455 154910 402464
rect 154762 402248 154818 402257
rect 154762 402183 154818 402192
rect 154960 401713 154988 402630
rect 154946 401704 155002 401713
rect 154946 401639 155002 401648
rect 154856 401532 154908 401538
rect 154856 401474 154908 401480
rect 154868 401169 154896 401474
rect 155040 401464 155092 401470
rect 155144 401441 155172 402946
rect 155224 402484 155276 402490
rect 155224 402426 155276 402432
rect 155236 401985 155264 402426
rect 155222 401976 155278 401985
rect 155222 401911 155278 401920
rect 155224 401600 155276 401606
rect 155224 401542 155276 401548
rect 155040 401406 155092 401412
rect 155130 401432 155186 401441
rect 154948 401396 155000 401402
rect 154948 401338 155000 401344
rect 154854 401160 154910 401169
rect 154854 401095 154910 401104
rect 154960 400897 154988 401338
rect 154946 400888 155002 400897
rect 154946 400823 155002 400832
rect 155052 400353 155080 401406
rect 155130 401367 155186 401376
rect 155132 400920 155184 400926
rect 155132 400862 155184 400868
rect 155038 400344 155094 400353
rect 155038 400279 155094 400288
rect 154764 400172 154816 400178
rect 154764 400114 154816 400120
rect 154776 399265 154804 400114
rect 155040 400104 155092 400110
rect 154946 400072 155002 400081
rect 154856 400036 154908 400042
rect 155040 400046 155092 400052
rect 154946 400007 155002 400016
rect 154856 399978 154908 399984
rect 154868 399809 154896 399978
rect 154960 399974 154988 400007
rect 154948 399968 155000 399974
rect 154948 399910 155000 399916
rect 154854 399800 154910 399809
rect 154854 399735 154910 399744
rect 155052 399537 155080 400046
rect 155038 399528 155094 399537
rect 155038 399463 155094 399472
rect 154762 399256 154818 399265
rect 154762 399191 154818 399200
rect 155144 398993 155172 400862
rect 155236 400625 155264 401542
rect 155222 400616 155278 400625
rect 155222 400551 155278 400560
rect 155130 398984 155186 398993
rect 155130 398919 155186 398928
rect 154580 398812 154632 398818
rect 154580 398754 154632 398760
rect 154592 398449 154620 398754
rect 154672 398744 154724 398750
rect 154672 398686 154724 398692
rect 154946 398712 155002 398721
rect 154578 398440 154634 398449
rect 154578 398375 154634 398384
rect 154684 397633 154712 398686
rect 154856 398676 154908 398682
rect 154946 398647 155002 398656
rect 154856 398618 154908 398624
rect 154868 398177 154896 398618
rect 154960 398546 154988 398647
rect 155040 398608 155092 398614
rect 155040 398550 155092 398556
rect 154948 398540 155000 398546
rect 154948 398482 155000 398488
rect 154854 398168 154910 398177
rect 154764 398132 154816 398138
rect 154854 398103 154910 398112
rect 154764 398074 154816 398080
rect 154670 397624 154726 397633
rect 154670 397559 154726 397568
rect 154776 396545 154804 398074
rect 155052 397905 155080 398550
rect 155038 397896 155094 397905
rect 155038 397831 155094 397840
rect 155040 397452 155092 397458
rect 155040 397394 155092 397400
rect 154946 397352 155002 397361
rect 154856 397316 154908 397322
rect 154946 397287 155002 397296
rect 154856 397258 154908 397264
rect 154868 396817 154896 397258
rect 154960 397254 154988 397287
rect 154948 397248 155000 397254
rect 154948 397190 155000 397196
rect 155052 397089 155080 397394
rect 155132 397384 155184 397390
rect 155132 397326 155184 397332
rect 155038 397080 155094 397089
rect 155038 397015 155094 397024
rect 154854 396808 154910 396817
rect 154854 396743 154910 396752
rect 154762 396536 154818 396545
rect 154762 396471 154818 396480
rect 155144 396273 155172 397326
rect 155130 396264 155186 396273
rect 155130 396199 155186 396208
rect 154764 396024 154816 396030
rect 155224 396024 155276 396030
rect 154764 395966 154816 395972
rect 154946 395992 155002 396001
rect 154672 395752 154724 395758
rect 154670 395720 154672 395729
rect 154724 395720 154726 395729
rect 154670 395655 154726 395664
rect 154776 395185 154804 395966
rect 154856 395956 154908 395962
rect 155224 395966 155276 395972
rect 154946 395927 155002 395936
rect 154856 395898 154908 395904
rect 154868 395457 154896 395898
rect 154960 395894 154988 395927
rect 154948 395888 155000 395894
rect 154948 395830 155000 395836
rect 155040 395820 155092 395826
rect 155040 395762 155092 395768
rect 154854 395448 154910 395457
rect 154854 395383 154910 395392
rect 154948 395344 155000 395350
rect 154948 395286 155000 395292
rect 154762 395176 154818 395185
rect 154762 395111 154818 395120
rect 154580 394664 154632 394670
rect 154580 394606 154632 394612
rect 154670 394632 154726 394641
rect 154592 394369 154620 394606
rect 154670 394567 154672 394576
rect 154724 394567 154726 394576
rect 154672 394538 154724 394544
rect 154764 394528 154816 394534
rect 154764 394470 154816 394476
rect 154578 394360 154634 394369
rect 154578 394295 154634 394304
rect 154776 394097 154804 394470
rect 154856 394460 154908 394466
rect 154856 394402 154908 394408
rect 154762 394088 154818 394097
rect 154762 394023 154818 394032
rect 154868 393553 154896 394402
rect 154960 393825 154988 395286
rect 155052 394913 155080 395762
rect 155038 394904 155094 394913
rect 155038 394839 155094 394848
rect 155132 393984 155184 393990
rect 155132 393926 155184 393932
rect 154946 393816 155002 393825
rect 154946 393751 155002 393760
rect 154854 393544 154910 393553
rect 154854 393479 154910 393488
rect 155040 393304 155092 393310
rect 154946 393272 155002 393281
rect 155040 393246 155092 393252
rect 154946 393207 154948 393216
rect 155000 393207 155002 393216
rect 154948 393178 155000 393184
rect 154764 393168 154816 393174
rect 154764 393110 154816 393116
rect 154776 392193 154804 393110
rect 154856 393100 154908 393106
rect 154856 393042 154908 393048
rect 154868 392465 154896 393042
rect 154948 393032 155000 393038
rect 155052 393009 155080 393246
rect 154948 392974 155000 392980
rect 155038 393000 155094 393009
rect 154960 392737 154988 392974
rect 155038 392935 155094 392944
rect 154946 392728 155002 392737
rect 154946 392663 155002 392672
rect 154854 392456 154910 392465
rect 154854 392391 154910 392400
rect 154762 392184 154818 392193
rect 154762 392119 154818 392128
rect 154946 391912 155002 391921
rect 154946 391847 154948 391856
rect 155000 391847 155002 391856
rect 154948 391818 155000 391824
rect 154764 391808 154816 391814
rect 154764 391750 154816 391756
rect 154672 391740 154724 391746
rect 154672 391682 154724 391688
rect 154684 391649 154712 391682
rect 154670 391640 154726 391649
rect 154670 391575 154726 391584
rect 154776 391377 154804 391750
rect 154948 391672 155000 391678
rect 154948 391614 155000 391620
rect 154762 391368 154818 391377
rect 154762 391303 154818 391312
rect 154960 391105 154988 391614
rect 154946 391096 155002 391105
rect 154946 391031 155002 391040
rect 154946 390552 155002 390561
rect 154580 390516 154632 390522
rect 154946 390487 155002 390496
rect 154580 390458 154632 390464
rect 154592 389473 154620 390458
rect 154960 390386 154988 390487
rect 155040 390448 155092 390454
rect 155040 390390 155092 390396
rect 154948 390380 155000 390386
rect 154948 390322 155000 390328
rect 154856 390312 154908 390318
rect 154856 390254 154908 390260
rect 154868 389745 154896 390254
rect 154948 390244 155000 390250
rect 154948 390186 155000 390192
rect 154960 390017 154988 390186
rect 154946 390008 155002 390017
rect 154946 389943 155002 389952
rect 154854 389736 154910 389745
rect 154854 389671 154910 389680
rect 154578 389464 154634 389473
rect 154578 389399 154634 389408
rect 155052 389201 155080 390390
rect 155144 389994 155172 393926
rect 155236 390289 155264 395966
rect 155222 390280 155278 390289
rect 155222 390215 155278 390224
rect 155144 389966 155356 389994
rect 155224 389836 155276 389842
rect 155224 389778 155276 389784
rect 155038 389192 155094 389201
rect 154856 389156 154908 389162
rect 155038 389127 155094 389136
rect 154856 389098 154908 389104
rect 154764 389088 154816 389094
rect 154764 389030 154816 389036
rect 154672 389020 154724 389026
rect 154672 388962 154724 388968
rect 154684 388929 154712 388962
rect 154670 388920 154726 388929
rect 154670 388855 154726 388864
rect 154776 388657 154804 389030
rect 154762 388648 154818 388657
rect 154762 388583 154818 388592
rect 154868 388113 154896 389098
rect 154948 388952 155000 388958
rect 154948 388894 155000 388900
rect 154960 388385 154988 388894
rect 154946 388376 155002 388385
rect 154946 388311 155002 388320
rect 154854 388104 154910 388113
rect 154854 388039 154910 388048
rect 155236 387841 155264 389778
rect 155222 387832 155278 387841
rect 155132 387796 155184 387802
rect 155222 387767 155278 387776
rect 155132 387738 155184 387744
rect 154948 387728 155000 387734
rect 154948 387670 155000 387676
rect 154764 387660 154816 387666
rect 154764 387602 154816 387608
rect 154776 386753 154804 387602
rect 154856 387592 154908 387598
rect 154960 387569 154988 387670
rect 154856 387534 154908 387540
rect 154946 387560 155002 387569
rect 154868 387297 154896 387534
rect 154946 387495 155002 387504
rect 155040 387524 155092 387530
rect 155040 387466 155092 387472
rect 154854 387288 154910 387297
rect 154854 387223 154910 387232
rect 155052 387025 155080 387466
rect 155038 387016 155094 387025
rect 155038 386951 155094 386960
rect 154762 386744 154818 386753
rect 154762 386679 154818 386688
rect 155144 386481 155172 387738
rect 155130 386472 155186 386481
rect 155130 386407 155186 386416
rect 155040 386368 155092 386374
rect 155040 386310 155092 386316
rect 154672 386300 154724 386306
rect 154672 386242 154724 386248
rect 154684 385937 154712 386242
rect 154856 386232 154908 386238
rect 154856 386174 154908 386180
rect 154946 386200 155002 386209
rect 154670 385928 154726 385937
rect 154670 385863 154726 385872
rect 154868 385393 154896 386174
rect 154946 386135 154948 386144
rect 155000 386135 155002 386144
rect 154948 386106 155000 386112
rect 154854 385384 154910 385393
rect 154854 385319 154910 385328
rect 155052 385121 155080 386310
rect 155224 385688 155276 385694
rect 155328 385665 155356 389966
rect 155224 385630 155276 385636
rect 155314 385656 155370 385665
rect 155038 385112 155094 385121
rect 155038 385047 155094 385056
rect 155132 385008 155184 385014
rect 155132 384950 155184 384956
rect 155040 384940 155092 384946
rect 155040 384882 155092 384888
rect 154948 384872 155000 384878
rect 154946 384840 154948 384849
rect 155000 384840 155002 384849
rect 154856 384804 154908 384810
rect 154946 384775 155002 384784
rect 154856 384746 154908 384752
rect 154672 384736 154724 384742
rect 154672 384678 154724 384684
rect 154684 383761 154712 384678
rect 154868 384033 154896 384746
rect 155052 384577 155080 384882
rect 155038 384568 155094 384577
rect 155038 384503 155094 384512
rect 155144 384305 155172 384950
rect 155130 384296 155186 384305
rect 155130 384231 155186 384240
rect 154854 384024 154910 384033
rect 154854 383959 154910 383968
rect 154670 383752 154726 383761
rect 154670 383687 154726 383696
rect 155236 383654 155264 385630
rect 155314 385591 155370 385600
rect 155236 383626 155356 383654
rect 154856 383580 154908 383586
rect 154856 383522 154908 383528
rect 154672 383444 154724 383450
rect 154672 383386 154724 383392
rect 154684 382401 154712 383386
rect 154868 383217 154896 383522
rect 154948 383512 155000 383518
rect 154946 383480 154948 383489
rect 155000 383480 155002 383489
rect 154946 383415 155002 383424
rect 154948 383376 155000 383382
rect 154948 383318 155000 383324
rect 154854 383208 154910 383217
rect 154854 383143 154910 383152
rect 154960 382673 154988 383318
rect 154946 382664 155002 382673
rect 154946 382599 155002 382608
rect 154670 382392 154726 382401
rect 154670 382327 154726 382336
rect 154948 382220 155000 382226
rect 154948 382162 155000 382168
rect 154580 382152 154632 382158
rect 154960 382129 154988 382162
rect 154580 382094 154632 382100
rect 154946 382120 155002 382129
rect 154592 381857 154620 382094
rect 154856 382084 154908 382090
rect 154946 382055 155002 382064
rect 154856 382026 154908 382032
rect 154578 381848 154634 381857
rect 154578 381783 154634 381792
rect 154868 381585 154896 382026
rect 154948 382016 155000 382022
rect 154948 381958 155000 381964
rect 154854 381576 154910 381585
rect 154854 381511 154910 381520
rect 154960 381313 154988 381958
rect 154946 381304 155002 381313
rect 154946 381239 155002 381248
rect 154948 380860 155000 380866
rect 154948 380802 155000 380808
rect 154764 380792 154816 380798
rect 154960 380769 154988 380802
rect 154764 380734 154816 380740
rect 154946 380760 155002 380769
rect 154776 379953 154804 380734
rect 154946 380695 155002 380704
rect 155040 380724 155092 380730
rect 155040 380666 155092 380672
rect 154856 380656 154908 380662
rect 154856 380598 154908 380604
rect 154868 380225 154896 380598
rect 154948 380588 155000 380594
rect 154948 380530 155000 380536
rect 154960 380497 154988 380530
rect 154946 380488 155002 380497
rect 154946 380423 155002 380432
rect 154854 380216 154910 380225
rect 154854 380151 154910 380160
rect 154762 379944 154818 379953
rect 154762 379879 154818 379888
rect 155052 379681 155080 380666
rect 155038 379672 155094 379681
rect 155038 379607 155094 379616
rect 154856 379432 154908 379438
rect 154856 379374 154908 379380
rect 154946 379400 155002 379409
rect 154868 379137 154896 379374
rect 154946 379335 154948 379344
rect 155000 379335 155002 379344
rect 154948 379306 155000 379312
rect 155040 379296 155092 379302
rect 155040 379238 155092 379244
rect 154948 379228 155000 379234
rect 154948 379170 155000 379176
rect 154854 379128 154910 379137
rect 154854 379063 154910 379072
rect 154960 378865 154988 379170
rect 154946 378856 155002 378865
rect 154672 378820 154724 378826
rect 154946 378791 155002 378800
rect 154672 378762 154724 378768
rect 154684 375601 154712 378762
rect 155052 378321 155080 379238
rect 155038 378312 155094 378321
rect 155038 378247 155094 378256
rect 154948 378140 155000 378146
rect 154948 378082 155000 378088
rect 154960 378049 154988 378082
rect 155040 378072 155092 378078
rect 154946 378040 155002 378049
rect 154764 378004 154816 378010
rect 155040 378014 155092 378020
rect 154946 377975 155002 377984
rect 154764 377946 154816 377952
rect 154776 377233 154804 377946
rect 154856 377936 154908 377942
rect 154856 377878 154908 377884
rect 154762 377224 154818 377233
rect 154762 377159 154818 377168
rect 154868 376961 154896 377878
rect 154948 377868 155000 377874
rect 154948 377810 155000 377816
rect 154960 377777 154988 377810
rect 154946 377768 155002 377777
rect 154946 377703 155002 377712
rect 155052 377505 155080 378014
rect 155038 377496 155094 377505
rect 155038 377431 155094 377440
rect 154854 376952 154910 376961
rect 154854 376887 154910 376896
rect 154948 376712 155000 376718
rect 154946 376680 154948 376689
rect 155000 376680 155002 376689
rect 154946 376615 155002 376624
rect 155040 376644 155092 376650
rect 155040 376586 155092 376592
rect 154856 376576 154908 376582
rect 154856 376518 154908 376524
rect 154868 376145 154896 376518
rect 154948 376508 155000 376514
rect 154948 376450 155000 376456
rect 154960 376417 154988 376450
rect 154946 376408 155002 376417
rect 154946 376343 155002 376352
rect 154854 376136 154910 376145
rect 154854 376071 154910 376080
rect 155052 375873 155080 376586
rect 155132 376032 155184 376038
rect 155132 375974 155184 375980
rect 155038 375864 155094 375873
rect 155038 375799 155094 375808
rect 154670 375592 154726 375601
rect 154670 375527 154726 375536
rect 154580 375420 154632 375426
rect 154580 375362 154632 375368
rect 154120 375352 154172 375358
rect 154120 375294 154172 375300
rect 154592 374785 154620 375362
rect 155040 375352 155092 375358
rect 154946 375320 155002 375329
rect 155040 375294 155092 375300
rect 154946 375255 154948 375264
rect 155000 375255 155002 375264
rect 154948 375226 155000 375232
rect 154856 375216 154908 375222
rect 154856 375158 154908 375164
rect 154868 375057 154896 375158
rect 154854 375048 154910 375057
rect 154854 374983 154910 374992
rect 154578 374776 154634 374785
rect 154578 374711 154634 374720
rect 154672 373992 154724 373998
rect 154578 373960 154634 373969
rect 154672 373934 154724 373940
rect 154578 373895 154634 373904
rect 154592 373862 154620 373895
rect 154580 373856 154632 373862
rect 154580 373798 154632 373804
rect 154684 372881 154712 373934
rect 154764 373924 154816 373930
rect 154764 373866 154816 373872
rect 154776 373153 154804 373866
rect 154948 373788 155000 373794
rect 154948 373730 155000 373736
rect 154856 373720 154908 373726
rect 154960 373697 154988 373730
rect 154856 373662 154908 373668
rect 154946 373688 155002 373697
rect 154868 373425 154896 373662
rect 154946 373623 155002 373632
rect 154854 373416 154910 373425
rect 154854 373351 154910 373360
rect 154762 373144 154818 373153
rect 154762 373079 154818 373088
rect 154670 372872 154726 372881
rect 154670 372807 154726 372816
rect 154946 372600 155002 372609
rect 154764 372564 154816 372570
rect 154946 372535 155002 372544
rect 154764 372506 154816 372512
rect 154776 372337 154804 372506
rect 154960 372502 154988 372535
rect 154948 372496 155000 372502
rect 154948 372438 155000 372444
rect 154948 372360 155000 372366
rect 154762 372328 154818 372337
rect 154948 372302 155000 372308
rect 154762 372263 154818 372272
rect 154856 372292 154908 372298
rect 154856 372234 154908 372240
rect 154868 371521 154896 372234
rect 154960 372065 154988 372302
rect 154946 372056 155002 372065
rect 154946 371991 155002 372000
rect 154854 371512 154910 371521
rect 154854 371447 154910 371456
rect 154764 371204 154816 371210
rect 154764 371146 154816 371152
rect 154672 371136 154724 371142
rect 154672 371078 154724 371084
rect 154684 370161 154712 371078
rect 154776 370433 154804 371146
rect 154948 371068 155000 371074
rect 154948 371010 155000 371016
rect 154856 371000 154908 371006
rect 154960 370977 154988 371010
rect 154856 370942 154908 370948
rect 154946 370968 155002 370977
rect 154868 370705 154896 370942
rect 154946 370903 155002 370912
rect 154854 370696 154910 370705
rect 154854 370631 154910 370640
rect 154762 370424 154818 370433
rect 154762 370359 154818 370368
rect 154670 370152 154726 370161
rect 154670 370087 154726 370096
rect 154672 369844 154724 369850
rect 154672 369786 154724 369792
rect 154684 368801 154712 369786
rect 154948 369708 155000 369714
rect 154948 369650 155000 369656
rect 154856 369640 154908 369646
rect 154960 369617 154988 369650
rect 154856 369582 154908 369588
rect 154946 369608 155002 369617
rect 154764 369572 154816 369578
rect 154764 369514 154816 369520
rect 154670 368792 154726 368801
rect 154670 368727 154726 368736
rect 154776 368529 154804 369514
rect 154868 369345 154896 369582
rect 154946 369543 155002 369552
rect 154854 369336 154910 369345
rect 154854 369271 154910 369280
rect 154762 368520 154818 368529
rect 154580 368484 154632 368490
rect 154762 368455 154818 368464
rect 154580 368426 154632 368432
rect 154592 368257 154620 368426
rect 154764 368416 154816 368422
rect 154764 368358 154816 368364
rect 154578 368248 154634 368257
rect 154578 368183 154634 368192
rect 154776 367441 154804 368358
rect 154948 368348 155000 368354
rect 154948 368290 155000 368296
rect 154856 368280 154908 368286
rect 154856 368222 154908 368228
rect 154762 367432 154818 367441
rect 154762 367367 154818 367376
rect 154868 367169 154896 368222
rect 154960 367985 154988 368290
rect 154946 367976 155002 367985
rect 154946 367911 155002 367920
rect 154854 367160 154910 367169
rect 154854 367095 154910 367104
rect 154948 366988 155000 366994
rect 154948 366930 155000 366936
rect 154672 366920 154724 366926
rect 154960 366897 154988 366930
rect 154672 366862 154724 366868
rect 154946 366888 155002 366897
rect 154684 366353 154712 366862
rect 154856 366852 154908 366858
rect 154946 366823 155002 366832
rect 154856 366794 154908 366800
rect 154670 366344 154726 366353
rect 154670 366279 154726 366288
rect 154868 366081 154896 366794
rect 154854 366072 154910 366081
rect 154854 366007 154910 366016
rect 154948 365696 155000 365702
rect 154948 365638 155000 365644
rect 154856 365560 154908 365566
rect 154670 365528 154726 365537
rect 154856 365502 154908 365508
rect 154670 365463 154672 365472
rect 154724 365463 154726 365472
rect 154672 365434 154724 365440
rect 154764 365424 154816 365430
rect 154764 365366 154816 365372
rect 154776 364993 154804 365366
rect 154762 364984 154818 364993
rect 154762 364919 154818 364928
rect 154868 364721 154896 365502
rect 154960 365265 154988 365638
rect 154946 365256 155002 365265
rect 154946 365191 155002 365200
rect 154854 364712 154910 364721
rect 154854 364647 154910 364656
rect 154764 364336 154816 364342
rect 155052 364334 155080 375294
rect 155144 374513 155172 375974
rect 155130 374504 155186 374513
rect 155130 374439 155186 374448
rect 155132 372428 155184 372434
rect 155132 372370 155184 372376
rect 155144 371793 155172 372370
rect 155130 371784 155186 371793
rect 155130 371719 155186 371728
rect 155130 371240 155186 371249
rect 155130 371175 155186 371184
rect 155144 370938 155172 371175
rect 155132 370932 155184 370938
rect 155132 370874 155184 370880
rect 155328 369889 155356 383626
rect 155420 374241 155448 497422
rect 155512 396030 155540 504358
rect 155592 480956 155644 480962
rect 155592 480898 155644 480904
rect 155500 396024 155552 396030
rect 155500 395966 155552 395972
rect 155500 387116 155552 387122
rect 155500 387058 155552 387064
rect 155512 381041 155540 387058
rect 155498 381032 155554 381041
rect 155498 380967 155554 380976
rect 155604 378842 155632 480898
rect 155684 450560 155736 450566
rect 155684 450502 155736 450508
rect 155696 407153 155724 450502
rect 156604 422340 156656 422346
rect 156604 422282 156656 422288
rect 155776 407788 155828 407794
rect 155776 407730 155828 407736
rect 155682 407144 155738 407153
rect 155682 407079 155738 407088
rect 155788 404433 155816 407730
rect 155774 404424 155830 404433
rect 155774 404359 155830 404368
rect 155512 378814 155632 378842
rect 155406 374232 155462 374241
rect 155406 374167 155462 374176
rect 155314 369880 155370 369889
rect 155314 369815 155370 369824
rect 155132 369776 155184 369782
rect 155132 369718 155184 369724
rect 155144 369073 155172 369718
rect 155130 369064 155186 369073
rect 155130 368999 155186 369008
rect 155316 367872 155368 367878
rect 155316 367814 155368 367820
rect 155132 367056 155184 367062
rect 155132 366998 155184 367004
rect 155144 366625 155172 366998
rect 155130 366616 155186 366625
rect 155130 366551 155186 366560
rect 155224 366376 155276 366382
rect 155224 366318 155276 366324
rect 155132 365628 155184 365634
rect 155132 365570 155184 365576
rect 155144 364449 155172 365570
rect 155130 364440 155186 364449
rect 155130 364375 155186 364384
rect 155052 364306 155172 364334
rect 154764 364278 154816 364284
rect 154776 363905 154804 364278
rect 155040 364268 155092 364274
rect 155040 364210 155092 364216
rect 154856 364200 154908 364206
rect 154856 364142 154908 364148
rect 154946 364168 155002 364177
rect 154762 363896 154818 363905
rect 154762 363831 154818 363840
rect 154868 363633 154896 364142
rect 154946 364103 154948 364112
rect 155000 364103 155002 364112
rect 154948 364074 155000 364080
rect 154854 363624 154910 363633
rect 154854 363559 154910 363568
rect 155052 363361 155080 364210
rect 155038 363352 155094 363361
rect 155038 363287 155094 363296
rect 154580 362908 154632 362914
rect 154580 362850 154632 362856
rect 154592 361729 154620 362850
rect 155040 362840 155092 362846
rect 154946 362808 155002 362817
rect 154856 362772 154908 362778
rect 155040 362782 155092 362788
rect 154946 362743 155002 362752
rect 154856 362714 154908 362720
rect 154868 362273 154896 362714
rect 154960 362710 154988 362743
rect 154948 362704 155000 362710
rect 154948 362646 155000 362652
rect 154854 362264 154910 362273
rect 154854 362199 154910 362208
rect 155052 362001 155080 362782
rect 155038 361992 155094 362001
rect 155038 361927 155094 361936
rect 154578 361720 154634 361729
rect 154578 361655 154634 361664
rect 155040 361548 155092 361554
rect 155040 361490 155092 361496
rect 154764 361480 154816 361486
rect 154764 361422 154816 361428
rect 154946 361448 155002 361457
rect 154580 361344 154632 361350
rect 154580 361286 154632 361292
rect 154592 361185 154620 361286
rect 154578 361176 154634 361185
rect 154578 361111 154634 361120
rect 154776 360641 154804 361422
rect 154856 361412 154908 361418
rect 154946 361383 155002 361392
rect 154856 361354 154908 361360
rect 154868 360913 154896 361354
rect 154960 361282 154988 361383
rect 154948 361276 155000 361282
rect 154948 361218 155000 361224
rect 154854 360904 154910 360913
rect 154854 360839 154910 360848
rect 154762 360632 154818 360641
rect 154762 360567 154818 360576
rect 155052 360369 155080 361490
rect 155038 360360 155094 360369
rect 155038 360295 155094 360304
rect 154580 360188 154632 360194
rect 154580 360130 154632 360136
rect 154592 359553 154620 360130
rect 155040 360120 155092 360126
rect 154946 360088 155002 360097
rect 155040 360062 155092 360068
rect 154946 360023 154948 360032
rect 155000 360023 155002 360032
rect 154948 359994 155000 360000
rect 154856 359984 154908 359990
rect 154856 359926 154908 359932
rect 154578 359544 154634 359553
rect 154578 359479 154634 359488
rect 154868 359281 154896 359926
rect 154948 359916 155000 359922
rect 154948 359858 155000 359864
rect 154854 359272 154910 359281
rect 154854 359207 154910 359216
rect 154960 359009 154988 359858
rect 155052 359825 155080 360062
rect 155038 359816 155094 359825
rect 155038 359751 155094 359760
rect 154946 359000 155002 359009
rect 154946 358935 155002 358944
rect 154578 358728 154634 358737
rect 154578 358663 154634 358672
rect 154948 358692 155000 358698
rect 154592 358562 154620 358663
rect 154948 358634 155000 358640
rect 154764 358624 154816 358630
rect 154764 358566 154816 358572
rect 154580 358556 154632 358562
rect 154580 358498 154632 358504
rect 154776 357649 154804 358566
rect 154960 357921 154988 358634
rect 155144 358465 155172 364306
rect 155236 363089 155264 366318
rect 155222 363080 155278 363089
rect 155222 363015 155278 363024
rect 155130 358456 155186 358465
rect 155130 358391 155186 358400
rect 154946 357912 155002 357921
rect 154946 357847 155002 357856
rect 154762 357640 154818 357649
rect 154762 357575 154818 357584
rect 155040 357400 155092 357406
rect 154946 357368 155002 357377
rect 154764 357332 154816 357338
rect 155040 357342 155092 357348
rect 154946 357303 155002 357312
rect 154764 357274 154816 357280
rect 154776 356289 154804 357274
rect 154960 357270 154988 357303
rect 154948 357264 155000 357270
rect 154948 357206 155000 357212
rect 154856 357196 154908 357202
rect 154856 357138 154908 357144
rect 154868 356561 154896 357138
rect 154948 357128 155000 357134
rect 155052 357105 155080 357342
rect 154948 357070 155000 357076
rect 155038 357096 155094 357105
rect 154960 356833 154988 357070
rect 155038 357031 155094 357040
rect 154946 356824 155002 356833
rect 154946 356759 155002 356768
rect 154854 356552 154910 356561
rect 154854 356487 154910 356496
rect 154762 356280 154818 356289
rect 154762 356215 154818 356224
rect 154580 356040 154632 356046
rect 154578 356008 154580 356017
rect 154632 356008 154634 356017
rect 154578 355943 154634 355952
rect 155040 355972 155092 355978
rect 155040 355914 155092 355920
rect 154856 355904 154908 355910
rect 154856 355846 154908 355852
rect 154868 355473 154896 355846
rect 154948 355836 155000 355842
rect 154948 355778 155000 355784
rect 154960 355745 154988 355778
rect 154946 355736 155002 355745
rect 154946 355671 155002 355680
rect 154854 355464 154910 355473
rect 154854 355399 154910 355408
rect 155052 355201 155080 355914
rect 155132 355360 155184 355366
rect 155132 355302 155184 355308
rect 155038 355192 155094 355201
rect 155038 355127 155094 355136
rect 154856 354680 154908 354686
rect 154578 354648 154634 354657
rect 154856 354622 154908 354628
rect 154578 354583 154580 354592
rect 154632 354583 154634 354592
rect 154580 354554 154632 354560
rect 154764 354476 154816 354482
rect 154764 354418 154816 354424
rect 154776 354113 154804 354418
rect 154762 354104 154818 354113
rect 154762 354039 154818 354048
rect 154868 353569 154896 354622
rect 154948 354544 155000 354550
rect 154948 354486 155000 354492
rect 154960 354385 154988 354486
rect 154946 354376 155002 354385
rect 154946 354311 155002 354320
rect 154854 353560 154910 353569
rect 154854 353495 154910 353504
rect 154854 353288 154910 353297
rect 154764 353252 154816 353258
rect 154854 353223 154910 353232
rect 154764 353194 154816 353200
rect 154776 352481 154804 353194
rect 154868 353122 154896 353223
rect 154948 353184 155000 353190
rect 154948 353126 155000 353132
rect 154856 353116 154908 353122
rect 154856 353058 154908 353064
rect 154960 353025 154988 353126
rect 155040 353048 155092 353054
rect 154946 353016 155002 353025
rect 154856 352980 154908 352986
rect 155040 352990 155092 352996
rect 154946 352951 155002 352960
rect 154856 352922 154908 352928
rect 154762 352472 154818 352481
rect 154762 352407 154818 352416
rect 154868 352209 154896 352922
rect 155052 352753 155080 352990
rect 155038 352744 155094 352753
rect 155038 352679 155094 352688
rect 154854 352200 154910 352209
rect 154854 352135 154910 352144
rect 154856 351892 154908 351898
rect 154856 351834 154908 351840
rect 154764 351688 154816 351694
rect 154764 351630 154816 351636
rect 154776 351393 154804 351630
rect 154762 351384 154818 351393
rect 154762 351319 154818 351328
rect 154868 351121 154896 351834
rect 154948 351824 155000 351830
rect 154948 351766 155000 351772
rect 154960 351665 154988 351766
rect 155040 351756 155092 351762
rect 155040 351698 155092 351704
rect 154946 351656 155002 351665
rect 154946 351591 155002 351600
rect 154854 351112 154910 351121
rect 154854 351047 154910 351056
rect 155052 350577 155080 351698
rect 155144 350849 155172 355302
rect 155328 354929 155356 367814
rect 155408 367804 155460 367810
rect 155408 367746 155460 367752
rect 155420 362545 155448 367746
rect 155512 367713 155540 378814
rect 155592 374672 155644 374678
rect 155592 374614 155644 374620
rect 155498 367704 155554 367713
rect 155498 367639 155554 367648
rect 155604 365809 155632 374614
rect 155590 365800 155646 365809
rect 155590 365735 155646 365744
rect 155406 362536 155462 362545
rect 155406 362471 155462 362480
rect 155408 362228 155460 362234
rect 155408 362170 155460 362176
rect 155314 354920 155370 354929
rect 155314 354855 155370 354864
rect 155420 351937 155448 362170
rect 155592 358760 155644 358766
rect 155592 358702 155644 358708
rect 155604 358193 155632 358702
rect 155590 358184 155646 358193
rect 155590 358119 155646 358128
rect 155592 355428 155644 355434
rect 155592 355370 155644 355376
rect 155604 353841 155632 355370
rect 155590 353832 155646 353841
rect 155590 353767 155646 353776
rect 155406 351928 155462 351937
rect 155406 351863 155462 351872
rect 155130 350840 155186 350849
rect 155130 350775 155186 350784
rect 155038 350568 155094 350577
rect 154580 350532 154632 350538
rect 155038 350503 155094 350512
rect 154580 350474 154632 350480
rect 154592 350305 154620 350474
rect 154948 350464 155000 350470
rect 154948 350406 155000 350412
rect 154578 350296 154634 350305
rect 154578 350231 154634 350240
rect 154960 350033 154988 350406
rect 154946 350024 155002 350033
rect 154946 349959 155002 349968
rect 154946 349752 155002 349761
rect 154946 349687 155002 349696
rect 154854 349480 154910 349489
rect 154854 349415 154910 349424
rect 154868 349178 154896 349415
rect 154960 349246 154988 349687
rect 154948 349240 155000 349246
rect 154948 349182 155000 349188
rect 155498 349208 155554 349217
rect 154856 349172 154908 349178
rect 155498 349143 155554 349152
rect 154856 349114 154908 349120
rect 155038 348936 155094 348945
rect 155038 348871 155094 348880
rect 154854 348664 154910 348673
rect 154854 348599 154910 348608
rect 154762 348392 154818 348401
rect 154762 348327 154818 348336
rect 154776 347886 154804 348327
rect 154868 348022 154896 348599
rect 154946 348120 155002 348129
rect 154946 348055 155002 348064
rect 154856 348016 154908 348022
rect 154856 347958 154908 347964
rect 154960 347954 154988 348055
rect 154948 347948 155000 347954
rect 154948 347890 155000 347896
rect 154764 347880 154816 347886
rect 154764 347822 154816 347828
rect 154946 347848 155002 347857
rect 155052 347818 155080 348871
rect 154946 347783 155002 347792
rect 155040 347812 155092 347818
rect 154854 347304 154910 347313
rect 154854 347239 154910 347248
rect 154578 347032 154634 347041
rect 154578 346967 154634 346976
rect 154592 346458 154620 346967
rect 154868 346662 154896 347239
rect 154960 347070 154988 347783
rect 155040 347754 155092 347760
rect 155038 347576 155094 347585
rect 155038 347511 155094 347520
rect 154948 347064 155000 347070
rect 154948 347006 155000 347012
rect 154946 346760 155002 346769
rect 154946 346695 155002 346704
rect 154856 346656 154908 346662
rect 154856 346598 154908 346604
rect 154960 346594 154988 346695
rect 154948 346588 155000 346594
rect 154948 346530 155000 346536
rect 155052 346526 155080 347511
rect 155040 346520 155092 346526
rect 154854 346488 154910 346497
rect 154580 346452 154632 346458
rect 155040 346462 155092 346468
rect 154854 346423 154910 346432
rect 154580 346394 154632 346400
rect 154868 345710 154896 346423
rect 155038 346216 155094 346225
rect 155038 346151 155094 346160
rect 154946 345944 155002 345953
rect 154946 345879 155002 345888
rect 154856 345704 154908 345710
rect 154856 345646 154908 345652
rect 154854 345536 154910 345545
rect 154854 345471 154910 345480
rect 154868 345014 154896 345471
rect 154960 345234 154988 345879
rect 154948 345228 155000 345234
rect 154948 345170 155000 345176
rect 155052 345166 155080 346151
rect 155040 345160 155092 345166
rect 154946 345128 155002 345137
rect 155040 345102 155092 345108
rect 154946 345063 154948 345072
rect 155000 345063 155002 345072
rect 154948 345034 155000 345040
rect 155512 345014 155540 349143
rect 155590 345400 155646 345409
rect 155590 345335 155646 345344
rect 154684 344986 154896 345014
rect 155420 344986 155540 345014
rect 154578 344040 154634 344049
rect 154578 343975 154634 343984
rect 154592 343874 154620 343975
rect 154580 343868 154632 343874
rect 154580 343810 154632 343816
rect 154578 343768 154634 343777
rect 154578 343703 154634 343712
rect 154592 342922 154620 343703
rect 154580 342916 154632 342922
rect 154580 342858 154632 342864
rect 154684 339538 154712 344986
rect 155038 344856 155094 344865
rect 155038 344791 155094 344800
rect 154946 344584 155002 344593
rect 154946 344519 155002 344528
rect 154854 344312 154910 344321
rect 154854 344247 154910 344256
rect 154868 343670 154896 344247
rect 154960 343806 154988 344519
rect 154948 343800 155000 343806
rect 154948 343742 155000 343748
rect 155052 343738 155080 344791
rect 155040 343732 155092 343738
rect 155040 343674 155092 343680
rect 154856 343664 154908 343670
rect 154856 343606 154908 343612
rect 155038 343496 155094 343505
rect 155038 343431 155094 343440
rect 154854 342952 154910 342961
rect 154854 342887 154910 342896
rect 154868 342446 154896 342887
rect 154856 342440 154908 342446
rect 154856 342382 154908 342388
rect 154946 342408 155002 342417
rect 154946 342343 154948 342352
rect 155000 342343 155002 342352
rect 154948 342314 155000 342320
rect 155052 342310 155080 343431
rect 155040 342304 155092 342310
rect 155040 342246 155092 342252
rect 154762 342136 154818 342145
rect 154762 342071 154818 342080
rect 154776 341086 154804 342071
rect 154946 341864 155002 341873
rect 154946 341799 155002 341808
rect 154854 341320 154910 341329
rect 154854 341255 154910 341264
rect 154764 341080 154816 341086
rect 154764 341022 154816 341028
rect 154868 340950 154896 341255
rect 154960 341154 154988 341799
rect 155038 341592 155094 341601
rect 155038 341527 155094 341536
rect 154948 341148 155000 341154
rect 154948 341090 155000 341096
rect 155052 341018 155080 341527
rect 155130 341048 155186 341057
rect 155040 341012 155092 341018
rect 155130 340983 155186 340992
rect 155040 340954 155092 340960
rect 154856 340944 154908 340950
rect 154856 340886 154908 340892
rect 155038 340776 155094 340785
rect 155038 340711 155094 340720
rect 154762 340504 154818 340513
rect 154762 340439 154818 340448
rect 154592 339510 154712 339538
rect 154776 339522 154804 340439
rect 154946 340232 155002 340241
rect 154946 340167 155002 340176
rect 154854 339960 154910 339969
rect 154854 339895 154910 339904
rect 154868 339726 154896 339895
rect 154960 339794 154988 340167
rect 154948 339788 155000 339794
rect 154948 339730 155000 339736
rect 154856 339720 154908 339726
rect 154856 339662 154908 339668
rect 154946 339688 155002 339697
rect 155052 339658 155080 340711
rect 154946 339623 155002 339632
rect 155040 339652 155092 339658
rect 154960 339590 154988 339623
rect 155040 339594 155092 339600
rect 154948 339584 155000 339590
rect 154948 339526 155000 339532
rect 154764 339516 154816 339522
rect 154592 338774 154620 339510
rect 154764 339458 154816 339464
rect 154670 339416 154726 339425
rect 154670 339351 154726 339360
rect 154580 338768 154632 338774
rect 154580 338710 154632 338716
rect 154684 338230 154712 339351
rect 154854 339144 154910 339153
rect 154854 339079 154910 339088
rect 154868 338298 154896 339079
rect 155038 338872 155094 338881
rect 155038 338807 155094 338816
rect 154946 338600 155002 338609
rect 154946 338535 155002 338544
rect 154960 338366 154988 338535
rect 154948 338360 155000 338366
rect 154948 338302 155000 338308
rect 154856 338292 154908 338298
rect 154856 338234 154908 338240
rect 154672 338224 154724 338230
rect 154672 338166 154724 338172
rect 155052 338162 155080 338807
rect 155040 338156 155092 338162
rect 155040 338098 155092 338104
rect 154762 338056 154818 338065
rect 154762 337991 154818 338000
rect 154578 337240 154634 337249
rect 154578 337175 154634 337184
rect 154592 337074 154620 337175
rect 154580 337068 154632 337074
rect 154580 337010 154632 337016
rect 154776 336938 154804 337991
rect 154854 337784 154910 337793
rect 154854 337719 154910 337728
rect 154868 337006 154896 337719
rect 155038 337512 155094 337521
rect 155038 337447 155094 337456
rect 154856 337000 154908 337006
rect 154856 336942 154908 336948
rect 154946 336968 155002 336977
rect 154764 336932 154816 336938
rect 154946 336903 155002 336912
rect 154764 336874 154816 336880
rect 154960 336870 154988 336903
rect 154948 336864 155000 336870
rect 154948 336806 155000 336812
rect 155052 336802 155080 337447
rect 155144 337414 155172 340983
rect 155316 340196 155368 340202
rect 155316 340138 155368 340144
rect 155222 338328 155278 338337
rect 155222 338263 155278 338272
rect 155132 337408 155184 337414
rect 155132 337350 155184 337356
rect 155040 336796 155092 336802
rect 155040 336738 155092 336744
rect 154762 336696 154818 336705
rect 154762 336631 154818 336640
rect 154670 336424 154726 336433
rect 154670 336359 154726 336368
rect 154684 335442 154712 336359
rect 154776 335646 154804 336631
rect 155038 336152 155094 336161
rect 155038 336087 155094 336096
rect 154854 335880 154910 335889
rect 154854 335815 154910 335824
rect 154764 335640 154816 335646
rect 154764 335582 154816 335588
rect 154868 335510 154896 335815
rect 154946 335608 155002 335617
rect 155052 335578 155080 336087
rect 154946 335543 155002 335552
rect 155040 335572 155092 335578
rect 154856 335504 154908 335510
rect 154856 335446 154908 335452
rect 154672 335436 154724 335442
rect 154672 335378 154724 335384
rect 154960 335374 154988 335543
rect 155040 335514 155092 335520
rect 155236 335458 155264 338263
rect 155052 335430 155264 335458
rect 154948 335368 155000 335374
rect 154948 335310 155000 335316
rect 154762 334792 154818 334801
rect 154762 334727 154818 334736
rect 154776 334082 154804 334727
rect 155052 334694 155080 335430
rect 155224 335368 155276 335374
rect 155224 335310 155276 335316
rect 155040 334688 155092 334694
rect 155040 334630 155092 334636
rect 155130 334520 155186 334529
rect 155130 334455 155186 334464
rect 154946 334248 155002 334257
rect 154946 334183 155002 334192
rect 154960 334150 154988 334183
rect 154948 334144 155000 334150
rect 154948 334086 155000 334092
rect 154764 334076 154816 334082
rect 154764 334018 154816 334024
rect 155144 334014 155172 334455
rect 155132 334008 155184 334014
rect 154854 333976 154910 333985
rect 155132 333950 155184 333956
rect 154854 333911 154910 333920
rect 154762 333432 154818 333441
rect 154762 333367 154818 333376
rect 154026 333160 154082 333169
rect 154026 333095 154082 333104
rect 153934 323912 153990 323921
rect 153934 323847 153990 323856
rect 153842 302696 153898 302705
rect 153842 302631 153898 302640
rect 153856 202162 153884 302631
rect 153948 249762 153976 323847
rect 154040 273222 154068 333095
rect 154776 332926 154804 333367
rect 154764 332920 154816 332926
rect 154578 332888 154634 332897
rect 154764 332862 154816 332868
rect 154578 332823 154580 332832
rect 154632 332823 154634 332832
rect 154580 332794 154632 332800
rect 154868 332722 154896 333911
rect 154946 333704 155002 333713
rect 154946 333639 155002 333648
rect 154960 332790 154988 333639
rect 154948 332784 155000 332790
rect 154948 332726 155000 332732
rect 154856 332716 154908 332722
rect 154856 332658 154908 332664
rect 154762 332616 154818 332625
rect 154762 332551 154818 332560
rect 154776 330546 154804 332551
rect 154946 332072 155002 332081
rect 154946 332007 155002 332016
rect 154854 331528 154910 331537
rect 154960 331498 154988 332007
rect 155038 331800 155094 331809
rect 155038 331735 155094 331744
rect 154854 331463 154910 331472
rect 154948 331492 155000 331498
rect 154868 331430 154896 331463
rect 154948 331434 155000 331440
rect 154856 331424 154908 331430
rect 154856 331366 154908 331372
rect 154948 331356 155000 331362
rect 154948 331298 155000 331304
rect 154960 331265 154988 331298
rect 155052 331294 155080 331735
rect 155040 331288 155092 331294
rect 154946 331256 155002 331265
rect 155040 331230 155092 331236
rect 154946 331191 155002 331200
rect 155038 330984 155094 330993
rect 155038 330919 155094 330928
rect 154764 330540 154816 330546
rect 154764 330482 154816 330488
rect 154854 330440 154910 330449
rect 154854 330375 154910 330384
rect 154868 330002 154896 330375
rect 154946 330168 155002 330177
rect 154946 330103 155002 330112
rect 154960 330070 154988 330103
rect 154948 330064 155000 330070
rect 154948 330006 155000 330012
rect 154856 329996 154908 330002
rect 154856 329938 154908 329944
rect 155052 329934 155080 330919
rect 155130 330712 155186 330721
rect 155130 330647 155186 330656
rect 155040 329928 155092 329934
rect 154578 329896 154634 329905
rect 155040 329870 155092 329876
rect 155144 329866 155172 330647
rect 154578 329831 154634 329840
rect 155132 329860 155184 329866
rect 154592 328778 154620 329831
rect 155132 329802 155184 329808
rect 154854 329624 154910 329633
rect 154854 329559 154910 329568
rect 154580 328772 154632 328778
rect 154580 328714 154632 328720
rect 154868 328642 154896 329559
rect 155130 329352 155186 329361
rect 155130 329287 155186 329296
rect 155038 329080 155094 329089
rect 155038 329015 155094 329024
rect 154946 328808 155002 328817
rect 154946 328743 155002 328752
rect 154960 328710 154988 328743
rect 154948 328704 155000 328710
rect 154948 328646 155000 328652
rect 154856 328636 154908 328642
rect 154856 328578 154908 328584
rect 154580 328568 154632 328574
rect 154578 328536 154580 328545
rect 154632 328536 154634 328545
rect 155052 328506 155080 329015
rect 154578 328471 154634 328480
rect 155040 328500 155092 328506
rect 155040 328442 155092 328448
rect 155038 328264 155094 328273
rect 155038 328199 155094 328208
rect 154670 327992 154726 328001
rect 154670 327927 154726 327936
rect 154580 325848 154632 325854
rect 154578 325816 154580 325825
rect 154632 325816 154634 325825
rect 154578 325751 154634 325760
rect 154578 321736 154634 321745
rect 154578 321671 154634 321680
rect 154592 318102 154620 321671
rect 154684 319462 154712 327927
rect 154854 327720 154910 327729
rect 154854 327655 154910 327664
rect 154764 327344 154816 327350
rect 154764 327286 154816 327292
rect 154776 327185 154804 327286
rect 154868 327214 154896 327655
rect 154946 327448 155002 327457
rect 154946 327383 155002 327392
rect 154960 327282 154988 327383
rect 154948 327276 155000 327282
rect 154948 327218 155000 327224
rect 154856 327208 154908 327214
rect 154762 327176 154818 327185
rect 154856 327150 154908 327156
rect 155052 327146 155080 328199
rect 154762 327111 154818 327120
rect 155040 327140 155092 327146
rect 155040 327082 155092 327088
rect 154854 326904 154910 326913
rect 154854 326839 154910 326848
rect 154762 326360 154818 326369
rect 154762 326295 154818 326304
rect 154776 325786 154804 326295
rect 154868 325990 154896 326839
rect 154946 326632 155002 326641
rect 154946 326567 155002 326576
rect 154856 325984 154908 325990
rect 154856 325926 154908 325932
rect 154960 325922 154988 326567
rect 155038 326088 155094 326097
rect 155038 326023 155094 326032
rect 154948 325916 155000 325922
rect 154948 325858 155000 325864
rect 154764 325780 154816 325786
rect 154764 325722 154816 325728
rect 155052 325718 155080 326023
rect 155040 325712 155092 325718
rect 155040 325654 155092 325660
rect 155038 325544 155094 325553
rect 155038 325479 155094 325488
rect 154762 325272 154818 325281
rect 154762 325207 154818 325216
rect 154776 324426 154804 325207
rect 154854 325000 154910 325009
rect 154854 324935 154910 324944
rect 154868 324494 154896 324935
rect 154946 324728 155002 324737
rect 154946 324663 155002 324672
rect 154960 324630 154988 324663
rect 154948 324624 155000 324630
rect 154948 324566 155000 324572
rect 155052 324562 155080 325479
rect 155040 324556 155092 324562
rect 155040 324498 155092 324504
rect 154856 324488 154908 324494
rect 154856 324430 154908 324436
rect 154946 324456 155002 324465
rect 154764 324420 154816 324426
rect 154946 324391 155002 324400
rect 154764 324362 154816 324368
rect 154960 324358 154988 324391
rect 154948 324352 155000 324358
rect 154948 324294 155000 324300
rect 155038 324184 155094 324193
rect 155038 324119 155094 324128
rect 154946 323640 155002 323649
rect 154946 323575 155002 323584
rect 154854 323368 154910 323377
rect 154854 323303 154910 323312
rect 154868 323066 154896 323303
rect 154960 323270 154988 323575
rect 154948 323264 155000 323270
rect 154948 323206 155000 323212
rect 155052 323202 155080 324119
rect 155040 323196 155092 323202
rect 155040 323138 155092 323144
rect 154948 323128 155000 323134
rect 154946 323096 154948 323105
rect 155000 323096 155002 323105
rect 154856 323060 154908 323066
rect 154946 323031 155002 323040
rect 154856 323002 154908 323008
rect 155038 322824 155094 322833
rect 155038 322759 155094 322768
rect 154762 322552 154818 322561
rect 154762 322487 154818 322496
rect 154776 321638 154804 322487
rect 154854 322280 154910 322289
rect 154854 322215 154910 322224
rect 154868 321842 154896 322215
rect 154946 322008 155002 322017
rect 154946 321943 155002 321952
rect 154856 321836 154908 321842
rect 154856 321778 154908 321784
rect 154960 321706 154988 321943
rect 155052 321774 155080 322759
rect 155040 321768 155092 321774
rect 155040 321710 155092 321716
rect 154948 321700 155000 321706
rect 154948 321642 155000 321648
rect 154764 321632 154816 321638
rect 154764 321574 154816 321580
rect 155038 321464 155094 321473
rect 155038 321399 155094 321408
rect 154762 321192 154818 321201
rect 154762 321127 154818 321136
rect 154776 320346 154804 321127
rect 154946 320920 155002 320929
rect 154946 320855 155002 320864
rect 154854 320648 154910 320657
rect 154854 320583 154910 320592
rect 154868 320414 154896 320583
rect 154960 320482 154988 320855
rect 154948 320476 155000 320482
rect 154948 320418 155000 320424
rect 154856 320408 154908 320414
rect 154856 320350 154908 320356
rect 154946 320376 155002 320385
rect 154764 320340 154816 320346
rect 154946 320311 155002 320320
rect 154764 320282 154816 320288
rect 154960 320278 154988 320311
rect 154948 320272 155000 320278
rect 154948 320214 155000 320220
rect 155052 320210 155080 321399
rect 155040 320204 155092 320210
rect 155040 320146 155092 320152
rect 154854 320104 154910 320113
rect 154854 320039 154910 320048
rect 154762 319832 154818 319841
rect 154762 319767 154818 319776
rect 154672 319456 154724 319462
rect 154672 319398 154724 319404
rect 154776 318986 154804 319767
rect 154868 319054 154896 320039
rect 155038 319560 155094 319569
rect 155038 319495 155094 319504
rect 154946 319288 155002 319297
rect 154946 319223 155002 319232
rect 154856 319048 154908 319054
rect 154856 318990 154908 318996
rect 154764 318980 154816 318986
rect 154764 318922 154816 318928
rect 154960 318918 154988 319223
rect 154948 318912 155000 318918
rect 154948 318854 155000 318860
rect 155052 318850 155080 319495
rect 155040 318844 155092 318850
rect 155040 318786 155092 318792
rect 154670 318744 154726 318753
rect 154670 318679 154726 318688
rect 154580 318096 154632 318102
rect 154580 318038 154632 318044
rect 154684 317490 154712 318679
rect 154762 318472 154818 318481
rect 154762 318407 154818 318416
rect 154776 317558 154804 318407
rect 155038 318200 155094 318209
rect 155038 318135 155094 318144
rect 154854 317928 154910 317937
rect 154854 317863 154910 317872
rect 154868 317762 154896 317863
rect 154856 317756 154908 317762
rect 154856 317698 154908 317704
rect 154948 317688 155000 317694
rect 154946 317656 154948 317665
rect 155000 317656 155002 317665
rect 155052 317626 155080 318135
rect 154946 317591 155002 317600
rect 155040 317620 155092 317626
rect 155040 317562 155092 317568
rect 154764 317552 154816 317558
rect 154764 317494 154816 317500
rect 154672 317484 154724 317490
rect 154672 317426 154724 317432
rect 154762 317384 154818 317393
rect 154762 317319 154818 317328
rect 154578 316840 154634 316849
rect 154578 316775 154634 316784
rect 154592 316402 154620 316775
rect 154580 316396 154632 316402
rect 154580 316338 154632 316344
rect 154776 316266 154804 317319
rect 154854 317112 154910 317121
rect 154854 317047 154910 317056
rect 154868 316334 154896 317047
rect 155038 316568 155094 316577
rect 155038 316503 155094 316512
rect 154856 316328 154908 316334
rect 154856 316270 154908 316276
rect 154946 316296 155002 316305
rect 154764 316260 154816 316266
rect 154946 316231 155002 316240
rect 154764 316202 154816 316208
rect 154960 316130 154988 316231
rect 155052 316198 155080 316503
rect 155040 316192 155092 316198
rect 155040 316134 155092 316140
rect 154948 316124 155000 316130
rect 154948 316066 155000 316072
rect 155038 316024 155094 316033
rect 155038 315959 155094 315968
rect 154854 315752 154910 315761
rect 154854 315687 154910 315696
rect 154762 315480 154818 315489
rect 154762 315415 154818 315424
rect 154776 314770 154804 315415
rect 154868 314838 154896 315687
rect 154946 315208 155002 315217
rect 154946 315143 155002 315152
rect 154856 314832 154908 314838
rect 154856 314774 154908 314780
rect 154764 314764 154816 314770
rect 154764 314706 154816 314712
rect 154960 314702 154988 315143
rect 155052 314906 155080 315959
rect 155040 314900 155092 314906
rect 155040 314842 155092 314848
rect 154948 314696 155000 314702
rect 154762 314664 154818 314673
rect 154948 314638 155000 314644
rect 154762 314599 154818 314608
rect 154578 313848 154634 313857
rect 154578 313783 154634 313792
rect 154592 313546 154620 313783
rect 154580 313540 154632 313546
rect 154580 313482 154632 313488
rect 154776 313342 154804 314599
rect 154854 314392 154910 314401
rect 154854 314327 154910 314336
rect 154868 313410 154896 314327
rect 154948 313608 155000 313614
rect 154946 313576 154948 313585
rect 155000 313576 155002 313585
rect 154946 313511 155002 313520
rect 154948 313472 155000 313478
rect 154948 313414 155000 313420
rect 154856 313404 154908 313410
rect 154856 313346 154908 313352
rect 154764 313336 154816 313342
rect 154960 313313 154988 313414
rect 154764 313278 154816 313284
rect 154946 313304 155002 313313
rect 154946 313239 155002 313248
rect 154854 313032 154910 313041
rect 154854 312967 154910 312976
rect 154762 312760 154818 312769
rect 154762 312695 154818 312704
rect 154578 312488 154634 312497
rect 154578 312423 154634 312432
rect 154592 312118 154620 312423
rect 154580 312112 154632 312118
rect 154580 312054 154632 312060
rect 154776 312050 154804 312695
rect 154764 312044 154816 312050
rect 154764 311986 154816 311992
rect 154868 311982 154896 312967
rect 154946 312216 155002 312225
rect 154946 312151 154948 312160
rect 155000 312151 155002 312160
rect 154948 312122 155000 312128
rect 154856 311976 154908 311982
rect 154578 311944 154634 311953
rect 154856 311918 154908 311924
rect 154578 311879 154580 311888
rect 154632 311879 154634 311888
rect 154580 311850 154632 311856
rect 154762 311672 154818 311681
rect 154762 311607 154818 311616
rect 154672 311228 154724 311234
rect 154672 311170 154724 311176
rect 154578 309768 154634 309777
rect 154578 309703 154634 309712
rect 154592 309262 154620 309703
rect 154580 309256 154632 309262
rect 154580 309198 154632 309204
rect 154578 308136 154634 308145
rect 154578 308071 154634 308080
rect 154592 305590 154620 308071
rect 154580 305584 154632 305590
rect 154580 305526 154632 305532
rect 154578 304056 154634 304065
rect 154578 303991 154634 304000
rect 154592 303822 154620 303991
rect 154580 303816 154632 303822
rect 154580 303758 154632 303764
rect 154684 302546 154712 311170
rect 154776 310622 154804 311607
rect 154854 311400 154910 311409
rect 154854 311335 154910 311344
rect 154868 310826 154896 311335
rect 155038 311128 155094 311137
rect 155038 311063 155094 311072
rect 154946 310856 155002 310865
rect 154856 310820 154908 310826
rect 154946 310791 155002 310800
rect 154856 310762 154908 310768
rect 154960 310758 154988 310791
rect 154948 310752 155000 310758
rect 154948 310694 155000 310700
rect 154856 310684 154908 310690
rect 154856 310626 154908 310632
rect 154764 310616 154816 310622
rect 154868 310593 154896 310626
rect 154764 310558 154816 310564
rect 154854 310584 154910 310593
rect 155052 310554 155080 311063
rect 154854 310519 154910 310528
rect 155040 310548 155092 310554
rect 155040 310490 155092 310496
rect 154854 310312 154910 310321
rect 154854 310247 154910 310256
rect 154762 310040 154818 310049
rect 154762 309975 154818 309984
rect 154776 309398 154804 309975
rect 154868 309466 154896 310247
rect 154946 309496 155002 309505
rect 154856 309460 154908 309466
rect 154946 309431 155002 309440
rect 154856 309402 154908 309408
rect 154764 309392 154816 309398
rect 154764 309334 154816 309340
rect 154960 309330 154988 309431
rect 154948 309324 155000 309330
rect 154948 309266 155000 309272
rect 154946 309224 155002 309233
rect 154946 309159 154948 309168
rect 155000 309159 155002 309168
rect 154948 309130 155000 309136
rect 155038 308952 155094 308961
rect 155038 308887 155094 308896
rect 154762 308680 154818 308689
rect 154762 308615 154818 308624
rect 154776 307970 154804 308615
rect 154854 308408 154910 308417
rect 154854 308343 154910 308352
rect 154764 307964 154816 307970
rect 154764 307906 154816 307912
rect 154868 307834 154896 308343
rect 154948 308032 155000 308038
rect 154948 307974 155000 307980
rect 154960 307873 154988 307974
rect 155052 307902 155080 308887
rect 155040 307896 155092 307902
rect 154946 307864 155002 307873
rect 154856 307828 154908 307834
rect 155040 307838 155092 307844
rect 154946 307799 155002 307808
rect 154856 307770 154908 307776
rect 155038 307592 155094 307601
rect 155038 307527 155094 307536
rect 154762 307320 154818 307329
rect 154762 307255 154818 307264
rect 154776 306406 154804 307255
rect 154946 307048 155002 307057
rect 154946 306983 155002 306992
rect 154854 306776 154910 306785
rect 154854 306711 154910 306720
rect 154868 306542 154896 306711
rect 154960 306610 154988 306983
rect 155052 306678 155080 307527
rect 155040 306672 155092 306678
rect 155040 306614 155092 306620
rect 154948 306604 155000 306610
rect 154948 306546 155000 306552
rect 154856 306536 154908 306542
rect 155040 306536 155092 306542
rect 154856 306478 154908 306484
rect 154946 306504 155002 306513
rect 155040 306478 155092 306484
rect 154946 306439 154948 306448
rect 155000 306439 155002 306448
rect 154948 306410 155000 306416
rect 154764 306400 154816 306406
rect 154764 306342 154816 306348
rect 154856 306400 154908 306406
rect 154908 306348 154988 306374
rect 154856 306346 154988 306348
rect 154856 306342 154908 306346
rect 154854 306232 154910 306241
rect 154854 306167 154910 306176
rect 154762 305960 154818 305969
rect 154762 305895 154818 305904
rect 154776 305114 154804 305895
rect 154868 305182 154896 306167
rect 154960 305522 154988 306346
rect 154948 305516 155000 305522
rect 154948 305458 155000 305464
rect 154946 305416 155002 305425
rect 154946 305351 155002 305360
rect 154856 305176 154908 305182
rect 154856 305118 154908 305124
rect 154764 305108 154816 305114
rect 154764 305050 154816 305056
rect 154960 305046 154988 305351
rect 154948 305040 155000 305046
rect 154948 304982 155000 304988
rect 154854 304872 154910 304881
rect 154854 304807 154910 304816
rect 154762 303784 154818 303793
rect 154868 303754 154896 304807
rect 154946 304600 155002 304609
rect 154946 304535 155002 304544
rect 154960 303890 154988 304535
rect 154948 303884 155000 303890
rect 154948 303826 155000 303832
rect 154762 303719 154818 303728
rect 154856 303748 154908 303754
rect 154776 302938 154804 303719
rect 154856 303690 154908 303696
rect 154946 303512 155002 303521
rect 154946 303447 155002 303456
rect 154854 302968 154910 302977
rect 154764 302932 154816 302938
rect 154854 302903 154910 302912
rect 154764 302874 154816 302880
rect 154592 302518 154712 302546
rect 154592 301442 154620 302518
rect 154672 302456 154724 302462
rect 154670 302424 154672 302433
rect 154724 302424 154726 302433
rect 154670 302359 154726 302368
rect 154868 302326 154896 302903
rect 154960 302530 154988 303447
rect 154948 302524 155000 302530
rect 154948 302466 155000 302472
rect 154856 302320 154908 302326
rect 154856 302262 154908 302268
rect 155052 302234 155080 306478
rect 155144 305250 155172 329287
rect 155132 305244 155184 305250
rect 155132 305186 155184 305192
rect 155130 305144 155186 305153
rect 155130 305079 155186 305088
rect 155144 304298 155172 305079
rect 155132 304292 155184 304298
rect 155132 304234 155184 304240
rect 155130 303240 155186 303249
rect 155130 303175 155186 303184
rect 155144 302394 155172 303175
rect 155132 302388 155184 302394
rect 155132 302330 155184 302336
rect 155052 302206 155172 302234
rect 154854 302152 154910 302161
rect 154854 302087 154910 302096
rect 154762 301880 154818 301889
rect 154762 301815 154818 301824
rect 154670 301608 154726 301617
rect 154670 301543 154726 301552
rect 154120 301436 154172 301442
rect 154120 301378 154172 301384
rect 154580 301436 154632 301442
rect 154580 301378 154632 301384
rect 154132 278730 154160 301378
rect 154578 301336 154634 301345
rect 154578 301271 154634 301280
rect 154592 301102 154620 301271
rect 154580 301096 154632 301102
rect 154580 301038 154632 301044
rect 154684 300898 154712 301543
rect 154776 300966 154804 301815
rect 154868 301034 154896 302087
rect 154856 301028 154908 301034
rect 154856 300970 154908 300976
rect 154764 300960 154816 300966
rect 154764 300902 154816 300908
rect 154672 300892 154724 300898
rect 154672 300834 154724 300840
rect 154854 300520 154910 300529
rect 154854 300455 154910 300464
rect 154762 300248 154818 300257
rect 154762 300183 154818 300192
rect 154670 299976 154726 299985
rect 154670 299911 154726 299920
rect 154684 299742 154712 299911
rect 154672 299736 154724 299742
rect 154578 299704 154634 299713
rect 154672 299678 154724 299684
rect 154578 299639 154580 299648
rect 154632 299639 154634 299648
rect 154580 299610 154632 299616
rect 154776 299606 154804 300183
rect 154764 299600 154816 299606
rect 154764 299542 154816 299548
rect 154868 299538 154896 300455
rect 154856 299532 154908 299538
rect 154856 299474 154908 299480
rect 154762 299432 154818 299441
rect 154762 299367 154818 299376
rect 154578 298888 154634 298897
rect 154578 298823 154634 298832
rect 154592 298246 154620 298823
rect 154670 298344 154726 298353
rect 154670 298279 154726 298288
rect 154580 298240 154632 298246
rect 154580 298182 154632 298188
rect 154578 297528 154634 297537
rect 154578 297463 154634 297472
rect 154592 296886 154620 297463
rect 154684 297430 154712 298279
rect 154776 298178 154804 299367
rect 154946 299160 155002 299169
rect 154946 299095 155002 299104
rect 154854 298616 154910 298625
rect 154854 298551 154910 298560
rect 154868 298314 154896 298551
rect 154960 298382 154988 299095
rect 154948 298376 155000 298382
rect 154948 298318 155000 298324
rect 154856 298308 154908 298314
rect 154856 298250 154908 298256
rect 154764 298172 154816 298178
rect 154764 298114 154816 298120
rect 154946 298072 155002 298081
rect 154946 298007 155002 298016
rect 154762 297800 154818 297809
rect 154762 297735 154818 297744
rect 154672 297424 154724 297430
rect 154672 297366 154724 297372
rect 154580 296880 154632 296886
rect 154580 296822 154632 296828
rect 154776 296818 154804 297735
rect 154764 296812 154816 296818
rect 154764 296754 154816 296760
rect 154960 296750 154988 298007
rect 155038 297256 155094 297265
rect 155038 297191 155094 297200
rect 154948 296744 155000 296750
rect 154854 296712 154910 296721
rect 154948 296686 155000 296692
rect 154854 296647 154910 296656
rect 154762 296168 154818 296177
rect 154762 296103 154818 296112
rect 154670 295896 154726 295905
rect 154670 295831 154726 295840
rect 154580 295656 154632 295662
rect 154578 295624 154580 295633
rect 154632 295624 154634 295633
rect 154578 295559 154634 295568
rect 154684 295458 154712 295831
rect 154776 295526 154804 296103
rect 154868 295594 154896 296647
rect 154946 296440 155002 296449
rect 154946 296375 155002 296384
rect 154856 295588 154908 295594
rect 154856 295530 154908 295536
rect 154764 295520 154816 295526
rect 154764 295462 154816 295468
rect 154672 295452 154724 295458
rect 154672 295394 154724 295400
rect 154960 295390 154988 296375
rect 154948 295384 155000 295390
rect 154948 295326 155000 295332
rect 154762 295080 154818 295089
rect 154762 295015 154818 295024
rect 154670 294808 154726 294817
rect 154670 294743 154726 294752
rect 154578 294264 154634 294273
rect 154684 294234 154712 294743
rect 154578 294199 154634 294208
rect 154672 294228 154724 294234
rect 154592 294166 154620 294199
rect 154672 294170 154724 294176
rect 154580 294160 154632 294166
rect 154580 294102 154632 294108
rect 154776 294098 154804 295015
rect 154854 294536 154910 294545
rect 154854 294471 154910 294480
rect 154868 294302 154896 294471
rect 154856 294296 154908 294302
rect 154856 294238 154908 294244
rect 154764 294092 154816 294098
rect 154764 294034 154816 294040
rect 154580 294024 154632 294030
rect 154578 293992 154580 294001
rect 154632 293992 154634 294001
rect 154578 293927 154634 293936
rect 154578 293720 154634 293729
rect 154578 293655 154634 293664
rect 154592 292738 154620 293655
rect 154670 293448 154726 293457
rect 154670 293383 154726 293392
rect 154580 292732 154632 292738
rect 154580 292674 154632 292680
rect 154684 292670 154712 293383
rect 155052 292754 155080 297191
rect 154868 292726 155080 292754
rect 154672 292664 154724 292670
rect 154578 292632 154634 292641
rect 154672 292606 154724 292612
rect 154578 292567 154580 292576
rect 154632 292567 154634 292576
rect 154868 292574 154896 292726
rect 154948 292664 155000 292670
rect 154948 292606 155000 292612
rect 154580 292538 154632 292544
rect 154684 292546 154896 292574
rect 154684 290494 154712 292546
rect 154672 290488 154724 290494
rect 154672 290430 154724 290436
rect 154960 282198 154988 292606
rect 155144 291854 155172 302206
rect 155236 296682 155264 335310
rect 155328 306474 155356 340138
rect 155420 333266 155448 344986
rect 155498 343224 155554 343233
rect 155498 343159 155554 343168
rect 155512 334626 155540 343159
rect 155604 340202 155632 345335
rect 155682 342680 155738 342689
rect 155682 342615 155738 342624
rect 155592 340196 155644 340202
rect 155592 340138 155644 340144
rect 155696 335374 155724 342615
rect 155684 335368 155736 335374
rect 155590 335336 155646 335345
rect 155684 335310 155736 335316
rect 155590 335271 155646 335280
rect 155500 334620 155552 334626
rect 155500 334562 155552 334568
rect 155408 333260 155460 333266
rect 155408 333202 155460 333208
rect 155604 325694 155632 335271
rect 155866 335064 155922 335073
rect 155866 334999 155922 335008
rect 155774 332344 155830 332353
rect 155774 332279 155830 332288
rect 155420 325666 155632 325694
rect 155420 311234 155448 325666
rect 155498 319016 155554 319025
rect 155498 318951 155554 318960
rect 155408 311228 155460 311234
rect 155408 311170 155460 311176
rect 155316 306468 155368 306474
rect 155316 306410 155368 306416
rect 155512 305658 155540 318951
rect 155590 314936 155646 314945
rect 155590 314871 155646 314880
rect 155604 311166 155632 314871
rect 155682 314120 155738 314129
rect 155682 314055 155738 314064
rect 155592 311160 155644 311166
rect 155592 311102 155644 311108
rect 155696 306542 155724 314055
rect 155684 306536 155736 306542
rect 155684 306478 155736 306484
rect 155590 305688 155646 305697
rect 155500 305652 155552 305658
rect 155590 305623 155646 305632
rect 155500 305594 155552 305600
rect 155316 305516 155368 305522
rect 155316 305458 155368 305464
rect 155328 303618 155356 305458
rect 155408 305244 155460 305250
rect 155408 305186 155460 305192
rect 155316 303612 155368 303618
rect 155316 303554 155368 303560
rect 155314 300792 155370 300801
rect 155314 300727 155370 300736
rect 155224 296676 155276 296682
rect 155224 296618 155276 296624
rect 155222 292904 155278 292913
rect 155222 292839 155278 292848
rect 155132 291848 155184 291854
rect 155132 291790 155184 291796
rect 154948 282192 155000 282198
rect 154948 282134 155000 282140
rect 154120 278724 154172 278730
rect 154120 278666 154172 278672
rect 154028 273216 154080 273222
rect 154028 273158 154080 273164
rect 153936 249756 153988 249762
rect 153936 249698 153988 249704
rect 153844 202156 153896 202162
rect 153844 202098 153896 202104
rect 155236 172514 155264 292839
rect 155328 292670 155356 300727
rect 155420 297226 155448 305186
rect 155498 304328 155554 304337
rect 155498 304263 155554 304272
rect 155512 303686 155540 304263
rect 155500 303680 155552 303686
rect 155500 303622 155552 303628
rect 155604 302234 155632 305623
rect 155684 305584 155736 305590
rect 155684 305526 155736 305532
rect 155512 302206 155632 302234
rect 155512 298790 155540 302206
rect 155590 301064 155646 301073
rect 155590 300999 155646 301008
rect 155500 298784 155552 298790
rect 155500 298726 155552 298732
rect 155408 297220 155460 297226
rect 155408 297162 155460 297168
rect 155498 296984 155554 296993
rect 155498 296919 155554 296928
rect 155406 295352 155462 295361
rect 155406 295287 155462 295296
rect 155316 292664 155368 292670
rect 155316 292606 155368 292612
rect 155314 292360 155370 292369
rect 155314 292295 155370 292304
rect 155224 172508 155276 172514
rect 155224 172450 155276 172456
rect 155328 171086 155356 292295
rect 155420 179382 155448 295287
rect 155512 182170 155540 296919
rect 155604 193186 155632 300999
rect 155696 209778 155724 305526
rect 155788 270502 155816 332279
rect 155880 277370 155908 334999
rect 155868 277364 155920 277370
rect 155868 277306 155920 277312
rect 155776 270496 155828 270502
rect 155776 270438 155828 270444
rect 155684 209772 155736 209778
rect 155684 209714 155736 209720
rect 155592 193180 155644 193186
rect 155592 193122 155644 193128
rect 155500 182164 155552 182170
rect 155500 182106 155552 182112
rect 155408 179376 155460 179382
rect 155408 179318 155460 179324
rect 155316 171080 155368 171086
rect 155316 171022 155368 171028
rect 155224 158024 155276 158030
rect 155224 157966 155276 157972
rect 154028 133680 154080 133686
rect 154028 133622 154080 133628
rect 153844 133544 153896 133550
rect 153844 133486 153896 133492
rect 153200 51740 153252 51746
rect 153200 51682 153252 51688
rect 152554 49192 152610 49201
rect 152554 49127 152610 49136
rect 152464 47524 152516 47530
rect 152464 47466 152516 47472
rect 151268 46776 151320 46782
rect 151268 46718 151320 46724
rect 153856 46714 153884 133486
rect 153936 133204 153988 133210
rect 153936 133146 153988 133152
rect 153948 48929 153976 133146
rect 154040 50454 154068 133622
rect 154120 133612 154172 133618
rect 154120 133554 154172 133560
rect 154132 51814 154160 133554
rect 154212 133476 154264 133482
rect 154212 133418 154264 133424
rect 154224 51950 154252 133418
rect 154948 130416 155000 130422
rect 154948 130358 155000 130364
rect 154960 129985 154988 130358
rect 154946 129976 155002 129985
rect 154946 129911 155002 129920
rect 154946 128072 155002 128081
rect 154946 128007 155002 128016
rect 154960 127634 154988 128007
rect 154948 127628 155000 127634
rect 154948 127570 155000 127576
rect 154946 126168 155002 126177
rect 154946 126103 155002 126112
rect 154960 125662 154988 126103
rect 154948 125656 155000 125662
rect 154948 125598 155000 125604
rect 154486 124264 154542 124273
rect 154486 124199 154542 124208
rect 154500 124166 154528 124199
rect 154488 124160 154540 124166
rect 154488 124102 154540 124108
rect 154946 122360 155002 122369
rect 154946 122295 155002 122304
rect 154960 121514 154988 122295
rect 154948 121508 155000 121514
rect 154948 121450 155000 121456
rect 154578 120456 154634 120465
rect 154578 120391 154634 120400
rect 154592 120154 154620 120391
rect 154580 120148 154632 120154
rect 154580 120090 154632 120096
rect 154578 118552 154634 118561
rect 154578 118487 154634 118496
rect 154592 117366 154620 118487
rect 154580 117360 154632 117366
rect 154580 117302 154632 117308
rect 154762 114744 154818 114753
rect 154762 114679 154818 114688
rect 154776 110430 154804 114679
rect 154946 112840 155002 112849
rect 154946 112775 155002 112784
rect 154854 110936 154910 110945
rect 154854 110871 154910 110880
rect 154764 110424 154816 110430
rect 154764 110366 154816 110372
rect 154578 105224 154634 105233
rect 154578 105159 154634 105168
rect 154592 104922 154620 105159
rect 154580 104916 154632 104922
rect 154580 104858 154632 104864
rect 154868 104854 154896 110871
rect 154960 107642 154988 112775
rect 154948 107636 155000 107642
rect 154948 107578 155000 107584
rect 154856 104848 154908 104854
rect 154856 104790 154908 104796
rect 154578 103320 154634 103329
rect 154578 103255 154634 103264
rect 154592 102202 154620 103255
rect 154580 102196 154632 102202
rect 154580 102138 154632 102144
rect 154946 101416 155002 101425
rect 154946 101351 155002 101360
rect 154960 100774 154988 101351
rect 154948 100768 155000 100774
rect 154948 100710 155000 100716
rect 154946 99512 155002 99521
rect 154946 99447 155002 99456
rect 154960 99414 154988 99447
rect 154948 99408 155000 99414
rect 154948 99350 155000 99356
rect 154854 97608 154910 97617
rect 154854 97543 154910 97552
rect 154868 94518 154896 97543
rect 154946 95704 155002 95713
rect 154946 95639 155002 95648
rect 154960 95266 154988 95639
rect 154948 95260 155000 95266
rect 154948 95202 155000 95208
rect 154856 94512 154908 94518
rect 154856 94454 154908 94460
rect 154578 93800 154634 93809
rect 154578 93735 154634 93744
rect 154592 92546 154620 93735
rect 154580 92540 154632 92546
rect 154580 92482 154632 92488
rect 154946 91896 155002 91905
rect 154946 91831 155002 91840
rect 154960 91118 154988 91831
rect 154948 91112 155000 91118
rect 154948 91054 155000 91060
rect 154946 89992 155002 90001
rect 154946 89927 155002 89936
rect 154960 89758 154988 89927
rect 154948 89752 155000 89758
rect 154948 89694 155000 89700
rect 154946 88088 155002 88097
rect 154946 88023 155002 88032
rect 154960 87038 154988 88023
rect 154948 87032 155000 87038
rect 154948 86974 155000 86980
rect 154946 86184 155002 86193
rect 154946 86119 155002 86128
rect 154960 85610 154988 86119
rect 154948 85604 155000 85610
rect 154948 85546 155000 85552
rect 154946 84280 155002 84289
rect 154946 84215 154948 84224
rect 155000 84215 155002 84224
rect 154948 84186 155000 84192
rect 154946 82376 155002 82385
rect 154946 82311 155002 82320
rect 154960 81462 154988 82311
rect 154948 81456 155000 81462
rect 154948 81398 155000 81404
rect 154762 80472 154818 80481
rect 154762 80407 154818 80416
rect 154776 80102 154804 80407
rect 154764 80096 154816 80102
rect 154764 80038 154816 80044
rect 154946 78568 155002 78577
rect 154946 78503 155002 78512
rect 154960 77314 154988 78503
rect 154948 77308 155000 77314
rect 154948 77250 155000 77256
rect 154946 76664 155002 76673
rect 154946 76599 155002 76608
rect 154960 75954 154988 76599
rect 154948 75948 155000 75954
rect 154948 75890 155000 75896
rect 154946 74760 155002 74769
rect 154946 74695 155002 74704
rect 154960 74594 154988 74695
rect 154948 74588 155000 74594
rect 154948 74530 155000 74536
rect 154578 72856 154634 72865
rect 154578 72791 154634 72800
rect 154592 71806 154620 72791
rect 154580 71800 154632 71806
rect 154580 71742 154632 71748
rect 154946 70952 155002 70961
rect 154946 70887 155002 70896
rect 154580 69080 154632 69086
rect 154578 69048 154580 69057
rect 154632 69048 154634 69057
rect 154578 68983 154634 68992
rect 154960 68338 154988 70887
rect 154948 68332 155000 68338
rect 154948 68274 155000 68280
rect 154946 67144 155002 67153
rect 154946 67079 155002 67088
rect 154960 66298 154988 67079
rect 154948 66292 155000 66298
rect 154948 66234 155000 66240
rect 154578 65240 154634 65249
rect 154578 65175 154634 65184
rect 154592 64938 154620 65175
rect 154580 64932 154632 64938
rect 154580 64874 154632 64880
rect 154578 63336 154634 63345
rect 154578 63271 154634 63280
rect 154592 62150 154620 63271
rect 154580 62144 154632 62150
rect 154580 62086 154632 62092
rect 154946 61432 155002 61441
rect 154946 61367 155002 61376
rect 154960 60790 154988 61367
rect 154948 60784 155000 60790
rect 154948 60726 155000 60732
rect 154946 59528 155002 59537
rect 154946 59463 155002 59472
rect 154960 59430 154988 59463
rect 154948 59424 155000 59430
rect 154948 59366 155000 59372
rect 154946 57624 155002 57633
rect 154946 57559 155002 57568
rect 154960 56642 154988 57559
rect 154948 56636 155000 56642
rect 154948 56578 155000 56584
rect 154946 55720 155002 55729
rect 154946 55655 155002 55664
rect 154960 55282 154988 55655
rect 154948 55276 155000 55282
rect 154948 55218 155000 55224
rect 154946 53816 155002 53825
rect 154946 53751 155002 53760
rect 154960 52494 154988 53751
rect 154948 52488 155000 52494
rect 154948 52430 155000 52436
rect 154212 51944 154264 51950
rect 154212 51886 154264 51892
rect 154120 51808 154172 51814
rect 154120 51750 154172 51756
rect 154028 50448 154080 50454
rect 154028 50390 154080 50396
rect 153934 48920 153990 48929
rect 153934 48855 153990 48864
rect 155236 48414 155264 157966
rect 155406 116648 155462 116657
rect 155406 116583 155462 116592
rect 155420 113150 155448 116583
rect 155408 113144 155460 113150
rect 155408 113086 155460 113092
rect 155498 109032 155554 109041
rect 155498 108967 155554 108976
rect 155314 107128 155370 107137
rect 155314 107063 155370 107072
rect 155328 100706 155356 107063
rect 155512 103494 155540 108967
rect 155500 103488 155552 103494
rect 155500 103430 155552 103436
rect 155316 100700 155368 100706
rect 155316 100642 155368 100648
rect 156616 52086 156644 422282
rect 156696 371272 156748 371278
rect 156696 371214 156748 371220
rect 156604 52080 156656 52086
rect 156604 52022 156656 52028
rect 156708 50862 156736 371214
rect 156788 357468 156840 357474
rect 156788 357410 156840 357416
rect 156696 50856 156748 50862
rect 156696 50798 156748 50804
rect 155224 48408 155276 48414
rect 155224 48350 155276 48356
rect 156800 48074 156828 357410
rect 157892 323604 157944 323610
rect 157892 323546 157944 323552
rect 156880 160744 156932 160750
rect 156880 160686 156932 160692
rect 156892 48482 156920 160686
rect 156972 149116 157024 149122
rect 156972 149058 157024 149064
rect 156880 48476 156932 48482
rect 156880 48418 156932 48424
rect 156984 48142 157012 149058
rect 157156 133340 157208 133346
rect 157156 133282 157208 133288
rect 157064 133272 157116 133278
rect 157064 133214 157116 133220
rect 157076 52630 157104 133214
rect 157064 52624 157116 52630
rect 157064 52566 157116 52572
rect 157168 52562 157196 133282
rect 157156 52556 157208 52562
rect 157156 52498 157208 52504
rect 157904 49609 157932 323546
rect 157996 52193 158024 700266
rect 158076 683188 158128 683194
rect 158076 683130 158128 683136
rect 157982 52184 158038 52193
rect 157982 52119 158038 52128
rect 158088 50153 158116 683130
rect 158168 632120 158220 632126
rect 158168 632062 158220 632068
rect 158074 50144 158130 50153
rect 158074 50079 158130 50088
rect 158076 50040 158128 50046
rect 158076 49982 158128 49988
rect 157890 49600 157946 49609
rect 157890 49535 157946 49544
rect 157800 49496 157852 49502
rect 157800 49438 157852 49444
rect 157708 49156 157760 49162
rect 157708 49098 157760 49104
rect 157616 49088 157668 49094
rect 157616 49030 157668 49036
rect 156972 48136 157024 48142
rect 156972 48078 157024 48084
rect 156788 48068 156840 48074
rect 156788 48010 156840 48016
rect 153844 46708 153896 46714
rect 153844 46650 153896 46656
rect 151176 46640 151228 46646
rect 151176 46582 151228 46588
rect 153200 46436 153252 46442
rect 153200 46378 153252 46384
rect 151820 43512 151872 43518
rect 151820 43454 151872 43460
rect 149058 35184 149114 35193
rect 149058 35119 149114 35128
rect 148416 28280 148468 28286
rect 148416 28222 148468 28228
rect 149072 16574 149100 35119
rect 144932 16546 145512 16574
rect 146312 16546 147168 16574
rect 147692 16546 147904 16574
rect 149072 16546 149560 16574
rect 144736 11688 144788 11694
rect 144736 11630 144788 11636
rect 143552 6886 143672 6914
rect 142436 3664 142488 3670
rect 142436 3606 142488 3612
rect 142448 480 142476 3606
rect 143552 480 143580 6886
rect 144748 480 144776 11630
rect 140014 354 140126 480
rect 139596 326 140126 354
rect 140014 -960 140126 326
rect 141210 -960 141322 480
rect 142406 -960 142518 480
rect 143510 -960 143622 480
rect 144706 -960 144818 480
rect 145484 354 145512 16546
rect 147140 480 147168 16546
rect 145902 354 146014 480
rect 145484 326 146014 354
rect 145902 -960 146014 326
rect 147098 -960 147210 480
rect 147876 354 147904 16546
rect 149532 480 149560 16546
rect 150624 3868 150676 3874
rect 150624 3810 150676 3816
rect 150636 480 150664 3810
rect 151832 480 151860 43454
rect 151912 26988 151964 26994
rect 151912 26930 151964 26936
rect 151924 16574 151952 26930
rect 153212 16574 153240 46378
rect 155960 45008 156012 45014
rect 155960 44950 156012 44956
rect 154580 36712 154632 36718
rect 154580 36654 154632 36660
rect 154592 16574 154620 36654
rect 155972 16574 156000 44950
rect 157340 43580 157392 43586
rect 157340 43522 157392 43528
rect 157352 16574 157380 43522
rect 157628 24614 157656 49030
rect 157616 24608 157668 24614
rect 157616 24550 157668 24556
rect 157720 23934 157748 49098
rect 157812 24818 157840 49438
rect 157984 49428 158036 49434
rect 157984 49370 158036 49376
rect 157800 24812 157852 24818
rect 157800 24754 157852 24760
rect 157708 23928 157760 23934
rect 157708 23870 157760 23876
rect 151924 16546 153056 16574
rect 153212 16546 153792 16574
rect 154592 16546 155448 16574
rect 155972 16546 156184 16574
rect 157352 16546 157840 16574
rect 153028 480 153056 16546
rect 148294 354 148406 480
rect 147876 326 148406 354
rect 148294 -960 148406 326
rect 149490 -960 149602 480
rect 150594 -960 150706 480
rect 151790 -960 151902 480
rect 152986 -960 153098 480
rect 153764 354 153792 16546
rect 155420 480 155448 16546
rect 154182 354 154294 480
rect 153764 326 154294 354
rect 154182 -960 154294 326
rect 155378 -960 155490 480
rect 156156 354 156184 16546
rect 157812 480 157840 16546
rect 157996 3466 158024 49370
rect 158088 3534 158116 49982
rect 158180 49910 158208 632062
rect 169772 429894 169800 702406
rect 202800 700330 202828 703520
rect 202788 700324 202840 700330
rect 202788 700266 202840 700272
rect 158444 429888 158496 429894
rect 158444 429830 158496 429836
rect 169760 429888 169812 429894
rect 169760 429830 169812 429836
rect 158260 327752 158312 327758
rect 158260 327694 158312 327700
rect 158168 49904 158220 49910
rect 158168 49846 158220 49852
rect 158168 49632 158220 49638
rect 158168 49574 158220 49580
rect 158180 3602 158208 49574
rect 158272 49065 158300 327694
rect 158352 159384 158404 159390
rect 158352 159326 158404 159332
rect 158364 49230 158392 159326
rect 158456 52698 158484 429830
rect 158732 270014 159436 270042
rect 160264 270014 160416 270042
rect 158732 151814 158760 270014
rect 160388 266422 160416 270014
rect 160480 270014 161092 270042
rect 161676 270014 161920 270042
rect 162412 270014 162748 270042
rect 162872 270014 163576 270042
rect 164252 270014 164404 270042
rect 164528 270014 165232 270042
rect 165632 270014 166060 270042
rect 166552 270014 166888 270042
rect 167012 270014 167716 270042
rect 168484 270014 168544 270042
rect 169036 270014 169372 270042
rect 169864 270014 170200 270042
rect 170692 270014 171028 270042
rect 171152 270014 171856 270042
rect 172532 270014 172684 270042
rect 172808 270014 173512 270042
rect 174004 270014 174340 270042
rect 174832 270014 175168 270042
rect 175292 270014 175996 270042
rect 176764 270014 176824 270042
rect 177316 270014 177652 270042
rect 178144 270014 178480 270042
rect 178972 270014 179308 270042
rect 179432 270014 180136 270042
rect 180812 270014 180964 270042
rect 181088 270014 181792 270042
rect 182192 270014 182620 270042
rect 183112 270014 183448 270042
rect 183572 270014 184276 270042
rect 184952 270014 185104 270042
rect 185228 270014 185932 270042
rect 186424 270014 186760 270042
rect 187252 270014 187588 270042
rect 187712 270014 188416 270042
rect 189092 270014 189244 270042
rect 189368 270014 190072 270042
rect 190564 270014 190900 270042
rect 191392 270014 191728 270042
rect 191852 270014 192556 270042
rect 193232 270014 193384 270042
rect 193508 270014 194212 270042
rect 194704 270014 195040 270042
rect 195532 270014 195868 270042
rect 195992 270014 196696 270042
rect 197372 270014 197524 270042
rect 197648 270014 198352 270042
rect 198752 270014 199180 270042
rect 199672 270014 200008 270042
rect 200132 270014 200836 270042
rect 201512 270014 201664 270042
rect 201788 270014 202492 270042
rect 202984 270014 203320 270042
rect 203812 270014 204148 270042
rect 204272 270014 204976 270042
rect 205652 270014 205804 270042
rect 205928 270014 206632 270042
rect 207032 270014 207460 270042
rect 207952 270014 208288 270042
rect 208412 270014 209116 270042
rect 209792 270014 209944 270042
rect 210068 270014 210772 270042
rect 211172 270014 211600 270042
rect 211724 270014 212428 270042
rect 212552 270014 213256 270042
rect 213932 270014 214084 270042
rect 214208 270014 214912 270042
rect 215404 270014 215740 270042
rect 216232 270014 216568 270042
rect 160376 266416 160428 266422
rect 160376 266358 160428 266364
rect 160480 258074 160508 270014
rect 161572 266416 161624 266422
rect 161572 266358 161624 266364
rect 161480 262948 161532 262954
rect 161480 262890 161532 262896
rect 160112 258046 160508 258074
rect 158732 151786 159036 151814
rect 159008 131866 159036 151786
rect 160112 131866 160140 258046
rect 161388 133952 161440 133958
rect 161388 133894 161440 133900
rect 161400 131866 161428 133894
rect 159008 131838 159436 131866
rect 160112 131838 160264 131866
rect 161092 131838 161428 131866
rect 161492 131866 161520 262890
rect 161584 132494 161612 266358
rect 161676 133958 161704 270014
rect 162412 262954 162440 270014
rect 162400 262948 162452 262954
rect 162400 262890 162452 262896
rect 162872 151814 162900 270014
rect 162872 151786 163176 151814
rect 161664 133952 161716 133958
rect 161664 133894 161716 133900
rect 161584 132466 162348 132494
rect 162320 131866 162348 132466
rect 163148 131866 163176 151786
rect 164252 131866 164280 270014
rect 164528 151814 164556 270014
rect 164528 151786 164832 151814
rect 164804 131866 164832 151786
rect 165632 131866 165660 270014
rect 166552 258074 166580 270014
rect 165724 258046 166580 258074
rect 165724 151814 165752 258046
rect 167012 151814 167040 270014
rect 168380 262948 168432 262954
rect 168380 262890 168432 262896
rect 165724 151786 166488 151814
rect 167012 151786 167316 151814
rect 166460 131866 166488 151786
rect 167288 131866 167316 151786
rect 168392 137358 168420 262890
rect 168380 137352 168432 137358
rect 168380 137294 168432 137300
rect 168484 131866 168512 270014
rect 169036 262954 169064 270014
rect 169024 262948 169076 262954
rect 169024 262890 169076 262896
rect 169760 262948 169812 262954
rect 169760 262890 169812 262896
rect 169772 137358 169800 262890
rect 169024 137352 169076 137358
rect 169024 137294 169076 137300
rect 169760 137352 169812 137358
rect 169760 137294 169812 137300
rect 169036 131866 169064 137294
rect 169864 131866 169892 270014
rect 170692 262954 170720 270014
rect 170680 262948 170732 262954
rect 170680 262890 170732 262896
rect 171152 151814 171180 270014
rect 171152 151786 171456 151814
rect 170680 137352 170732 137358
rect 170680 137294 170732 137300
rect 170692 131866 170720 137294
rect 171428 131866 171456 151786
rect 172532 131866 172560 270014
rect 172808 151814 172836 270014
rect 173900 262948 173952 262954
rect 173900 262890 173952 262896
rect 172808 151786 173112 151814
rect 173084 131866 173112 151786
rect 173912 139466 173940 262890
rect 173900 139460 173952 139466
rect 173900 139402 173952 139408
rect 174004 131866 174032 270014
rect 174832 262954 174860 270014
rect 174820 262948 174872 262954
rect 174820 262890 174872 262896
rect 175292 151814 175320 270014
rect 176660 262948 176712 262954
rect 176660 262890 176712 262896
rect 175292 151786 175596 151814
rect 174820 139460 174872 139466
rect 174820 139402 174872 139408
rect 174832 131866 174860 139402
rect 175568 131866 175596 151786
rect 176672 137358 176700 262890
rect 176660 137352 176712 137358
rect 176660 137294 176712 137300
rect 176764 131866 176792 270014
rect 177316 262954 177344 270014
rect 177304 262948 177356 262954
rect 177304 262890 177356 262896
rect 178040 262948 178092 262954
rect 178040 262890 178092 262896
rect 178052 140486 178080 262890
rect 178040 140480 178092 140486
rect 178040 140422 178092 140428
rect 177304 137352 177356 137358
rect 177304 137294 177356 137300
rect 177316 131866 177344 137294
rect 178144 131866 178172 270014
rect 178972 262954 179000 270014
rect 178960 262948 179012 262954
rect 178960 262890 179012 262896
rect 179432 151814 179460 270014
rect 179432 151786 179736 151814
rect 178960 140480 179012 140486
rect 178960 140422 179012 140428
rect 178972 131866 179000 140422
rect 179708 131866 179736 151786
rect 180812 131866 180840 270014
rect 181088 151814 181116 270014
rect 181088 151786 181392 151814
rect 181364 131866 181392 151786
rect 182192 131866 182220 270014
rect 183112 258074 183140 270014
rect 182284 258046 183140 258074
rect 182284 151814 182312 258046
rect 183572 151814 183600 270014
rect 182284 151786 183048 151814
rect 183572 151786 183876 151814
rect 183020 131866 183048 151786
rect 183848 131866 183876 151786
rect 184952 131866 184980 270014
rect 185228 151814 185256 270014
rect 186320 262948 186372 262954
rect 186320 262890 186372 262896
rect 185228 151786 185532 151814
rect 185504 131866 185532 151786
rect 186332 140690 186360 262890
rect 186320 140684 186372 140690
rect 186320 140626 186372 140632
rect 186424 131866 186452 270014
rect 187252 262954 187280 270014
rect 187240 262948 187292 262954
rect 187240 262890 187292 262896
rect 187712 151814 187740 270014
rect 187712 151786 188016 151814
rect 187240 140684 187292 140690
rect 187240 140626 187292 140632
rect 187252 131866 187280 140626
rect 187988 131866 188016 151786
rect 189092 131866 189120 270014
rect 189368 151814 189396 270014
rect 190460 262948 190512 262954
rect 190460 262890 190512 262896
rect 189368 151786 189672 151814
rect 189644 131866 189672 151786
rect 190472 137358 190500 262890
rect 190460 137352 190512 137358
rect 190460 137294 190512 137300
rect 190564 131866 190592 270014
rect 191392 262954 191420 270014
rect 191380 262948 191432 262954
rect 191380 262890 191432 262896
rect 191852 151814 191880 270014
rect 191852 151786 192156 151814
rect 191380 137352 191432 137358
rect 191380 137294 191432 137300
rect 191392 131866 191420 137294
rect 192128 131866 192156 151786
rect 193232 131866 193260 270014
rect 193508 151814 193536 270014
rect 194600 261316 194652 261322
rect 194600 261258 194652 261264
rect 193508 151786 193812 151814
rect 193784 131866 193812 151786
rect 194612 140758 194640 261258
rect 194600 140752 194652 140758
rect 194600 140694 194652 140700
rect 194704 131866 194732 270014
rect 195532 261322 195560 270014
rect 195520 261316 195572 261322
rect 195520 261258 195572 261264
rect 195992 151814 196020 270014
rect 195992 151786 196296 151814
rect 195520 140752 195572 140758
rect 195520 140694 195572 140700
rect 195532 131866 195560 140694
rect 196268 131866 196296 151786
rect 197372 131866 197400 270014
rect 197648 151814 197676 270014
rect 197648 151786 197952 151814
rect 197924 131866 197952 151786
rect 198752 131866 198780 270014
rect 199672 258074 199700 270014
rect 198844 258046 199700 258074
rect 198844 151814 198872 258046
rect 200132 151814 200160 270014
rect 198844 151786 199608 151814
rect 200132 151786 200436 151814
rect 199580 131866 199608 151786
rect 200408 131866 200436 151786
rect 201512 131866 201540 270014
rect 201788 151814 201816 270014
rect 202880 261316 202932 261322
rect 202880 261258 202932 261264
rect 201788 151786 202092 151814
rect 202064 131866 202092 151786
rect 202892 137358 202920 261258
rect 202880 137352 202932 137358
rect 202880 137294 202932 137300
rect 202984 131866 203012 270014
rect 203812 261322 203840 270014
rect 203800 261316 203852 261322
rect 203800 261258 203852 261264
rect 204272 151814 204300 270014
rect 204272 151786 204576 151814
rect 203800 137352 203852 137358
rect 203800 137294 203852 137300
rect 203812 131866 203840 137294
rect 204548 131866 204576 151786
rect 205652 131866 205680 270014
rect 205928 151814 205956 270014
rect 205928 151786 206232 151814
rect 206204 131866 206232 151786
rect 207032 131866 207060 270014
rect 207952 258074 207980 270014
rect 207124 258046 207980 258074
rect 207124 151814 207152 258046
rect 208412 151814 208440 270014
rect 207124 151786 207888 151814
rect 208412 151786 208716 151814
rect 207860 131866 207888 151786
rect 208688 131866 208716 151786
rect 209792 131866 209820 270014
rect 210068 151814 210096 270014
rect 210068 151786 210372 151814
rect 210344 131866 210372 151786
rect 211172 131866 211200 270014
rect 211724 258074 211752 270014
rect 211264 258046 211752 258074
rect 211264 151814 211292 258046
rect 212552 151814 212580 270014
rect 211264 151786 212028 151814
rect 212552 151786 212856 151814
rect 212000 131866 212028 151786
rect 212828 131866 212856 151786
rect 213932 131866 213960 270014
rect 214208 151814 214236 270014
rect 215300 260432 215352 260438
rect 215300 260374 215352 260380
rect 214208 151786 214512 151814
rect 214484 131866 214512 151786
rect 215312 139942 215340 260374
rect 215300 139936 215352 139942
rect 215300 139878 215352 139884
rect 215404 131866 215432 270014
rect 216232 260438 216260 270014
rect 216220 260432 216272 260438
rect 216220 260374 216272 260380
rect 216220 139936 216272 139942
rect 216220 139878 216272 139884
rect 216232 131866 216260 139878
rect 161492 131838 161920 131866
rect 162320 131838 162748 131866
rect 163148 131838 163576 131866
rect 164252 131838 164404 131866
rect 164804 131838 165232 131866
rect 165632 131838 166060 131866
rect 166460 131838 166888 131866
rect 167288 131838 167716 131866
rect 168484 131838 168544 131866
rect 169036 131838 169372 131866
rect 169864 131838 170200 131866
rect 170692 131838 171028 131866
rect 171428 131838 171856 131866
rect 172532 131838 172684 131866
rect 173084 131838 173512 131866
rect 174004 131838 174340 131866
rect 174832 131838 175168 131866
rect 175568 131838 175996 131866
rect 176764 131838 176824 131866
rect 177316 131838 177652 131866
rect 178144 131838 178480 131866
rect 178972 131838 179308 131866
rect 179708 131838 180136 131866
rect 180812 131838 180964 131866
rect 181364 131838 181792 131866
rect 182192 131838 182620 131866
rect 183020 131838 183448 131866
rect 183848 131838 184276 131866
rect 184952 131838 185104 131866
rect 185504 131838 185932 131866
rect 186424 131838 186760 131866
rect 187252 131838 187588 131866
rect 187988 131838 188416 131866
rect 189092 131838 189244 131866
rect 189644 131838 190072 131866
rect 190564 131838 190900 131866
rect 191392 131838 191728 131866
rect 192128 131838 192556 131866
rect 193232 131838 193384 131866
rect 193784 131838 194212 131866
rect 194704 131838 195040 131866
rect 195532 131838 195868 131866
rect 196268 131838 196696 131866
rect 197372 131838 197524 131866
rect 197924 131838 198352 131866
rect 198752 131838 199180 131866
rect 199580 131838 200008 131866
rect 200408 131838 200836 131866
rect 201512 131838 201664 131866
rect 202064 131838 202492 131866
rect 202984 131838 203320 131866
rect 203812 131838 204148 131866
rect 204548 131838 204976 131866
rect 205652 131838 205804 131866
rect 206204 131838 206632 131866
rect 207032 131838 207460 131866
rect 207860 131838 208288 131866
rect 208688 131838 209116 131866
rect 209792 131838 209944 131866
rect 210344 131838 210772 131866
rect 211172 131838 211600 131866
rect 212000 131838 212428 131866
rect 212828 131838 213256 131866
rect 213932 131838 214084 131866
rect 214484 131838 214912 131866
rect 215404 131838 215740 131866
rect 216232 131838 216568 131866
rect 216678 52864 216734 52873
rect 216678 52799 216680 52808
rect 216732 52799 216734 52808
rect 216680 52770 216732 52776
rect 216036 52760 216088 52766
rect 216036 52702 216088 52708
rect 175614 52698 175642 52700
rect 175890 52698 175918 52700
rect 177270 52698 177298 52700
rect 158444 52692 158496 52698
rect 158444 52634 158496 52640
rect 175602 52692 175654 52698
rect 175602 52634 175654 52640
rect 175878 52692 175930 52698
rect 175878 52634 175930 52640
rect 177258 52692 177310 52698
rect 177258 52634 177310 52640
rect 176994 52426 177022 52428
rect 200270 52426 200298 52428
rect 216048 52426 216076 52702
rect 159916 52420 159968 52426
rect 159916 52362 159968 52368
rect 176982 52420 177034 52426
rect 176982 52362 177034 52368
rect 200258 52420 200310 52426
rect 200258 52362 200310 52368
rect 216036 52420 216088 52426
rect 216036 52362 216088 52368
rect 159824 52080 159876 52086
rect 159824 52022 159876 52028
rect 159364 51672 159416 51678
rect 159364 51614 159416 51620
rect 159272 51536 159324 51542
rect 159272 51478 159324 51484
rect 159284 50794 159312 51478
rect 159376 51105 159404 51614
rect 159456 51400 159508 51406
rect 159456 51342 159508 51348
rect 159468 51202 159496 51342
rect 159836 51270 159864 52022
rect 159928 52018 159956 52362
rect 216220 52352 216272 52358
rect 216220 52294 216272 52300
rect 189494 52216 189546 52222
rect 189494 52158 189546 52164
rect 214426 52216 214478 52222
rect 214426 52158 214478 52164
rect 189506 52156 189534 52158
rect 214438 52156 214466 52158
rect 215924 52142 216076 52170
rect 182778 52080 182830 52086
rect 159916 52012 159968 52018
rect 159916 51954 159968 51960
rect 160020 52006 160080 52034
rect 182778 52022 182830 52028
rect 184342 52080 184394 52086
rect 184342 52022 184394 52028
rect 188114 52080 188166 52086
rect 188114 52022 188166 52028
rect 190414 52080 190466 52086
rect 190414 52022 190466 52028
rect 192254 52080 192306 52086
rect 192254 52022 192306 52028
rect 208630 52080 208682 52086
rect 208630 52022 208682 52028
rect 182790 52020 182818 52022
rect 184354 52020 184382 52022
rect 188126 52020 188154 52022
rect 190426 52020 190454 52022
rect 192266 52020 192294 52022
rect 208642 52020 208670 52022
rect 159914 51640 159970 51649
rect 159914 51575 159970 51584
rect 159824 51264 159876 51270
rect 159824 51206 159876 51212
rect 159456 51196 159508 51202
rect 159456 51138 159508 51144
rect 159362 51096 159418 51105
rect 159362 51031 159418 51040
rect 159824 50856 159876 50862
rect 159824 50798 159876 50804
rect 159272 50788 159324 50794
rect 159272 50730 159324 50736
rect 159836 50590 159864 50798
rect 159824 50584 159876 50590
rect 159824 50526 159876 50532
rect 159456 50176 159508 50182
rect 159456 50118 159508 50124
rect 158536 49972 158588 49978
rect 158536 49914 158588 49920
rect 158352 49224 158404 49230
rect 158352 49166 158404 49172
rect 158258 49056 158314 49065
rect 158258 48991 158314 49000
rect 158444 48476 158496 48482
rect 158444 48418 158496 48424
rect 158456 21486 158484 48418
rect 158548 24070 158576 49914
rect 158628 49700 158680 49706
rect 158628 49642 158680 49648
rect 158640 24342 158668 49642
rect 159468 49638 159496 50118
rect 159456 49632 159508 49638
rect 159456 49574 159508 49580
rect 159640 48680 159692 48686
rect 159640 48622 159692 48628
rect 159364 47796 159416 47802
rect 159364 47738 159416 47744
rect 158720 45484 158772 45490
rect 158720 45426 158772 45432
rect 158628 24336 158680 24342
rect 158628 24278 158680 24284
rect 158536 24064 158588 24070
rect 158536 24006 158588 24012
rect 158444 21480 158496 21486
rect 158444 21422 158496 21428
rect 158732 15910 158760 45426
rect 158720 15904 158772 15910
rect 158720 15846 158772 15852
rect 159376 4146 159404 47738
rect 159548 47456 159600 47462
rect 159548 47398 159600 47404
rect 159456 46980 159508 46986
rect 159456 46922 159508 46928
rect 159364 4140 159416 4146
rect 159364 4082 159416 4088
rect 159468 3806 159496 46922
rect 159560 21418 159588 47398
rect 159652 24274 159680 48622
rect 159732 48544 159784 48550
rect 159732 48486 159784 48492
rect 159640 24268 159692 24274
rect 159640 24210 159692 24216
rect 159744 24206 159772 48486
rect 159928 46510 159956 51575
rect 159916 46504 159968 46510
rect 159916 46446 159968 46452
rect 160020 45490 160048 52006
rect 160158 51864 160186 52020
rect 160112 51836 160186 51864
rect 160112 49434 160140 51836
rect 160250 51796 160278 52020
rect 160342 51921 160370 52020
rect 160328 51912 160384 51921
rect 160328 51847 160384 51856
rect 160204 51785 160278 51796
rect 160190 51776 160278 51785
rect 160246 51768 160278 51776
rect 160434 51728 160462 52020
rect 160526 51887 160554 52020
rect 160512 51878 160568 51887
rect 160512 51813 160568 51822
rect 160618 51728 160646 52020
rect 160710 51814 160738 52020
rect 160698 51808 160750 51814
rect 160698 51750 160750 51756
rect 160190 51711 160246 51720
rect 160388 51700 160462 51728
rect 160572 51700 160646 51728
rect 160192 51332 160244 51338
rect 160192 51274 160244 51280
rect 160204 51066 160232 51274
rect 160192 51060 160244 51066
rect 160192 51002 160244 51008
rect 160388 50538 160416 51700
rect 160572 51218 160600 51700
rect 160802 51660 160830 52020
rect 160894 51762 160922 52020
rect 160986 51921 161014 52020
rect 160972 51912 161028 51921
rect 161078 51882 161106 52020
rect 160972 51847 161028 51856
rect 161066 51876 161118 51882
rect 161066 51818 161118 51824
rect 161170 51785 161198 52020
rect 161156 51776 161212 51785
rect 160894 51734 161060 51762
rect 160650 51640 160706 51649
rect 160650 51575 160706 51584
rect 160756 51632 160830 51660
rect 160928 51672 160980 51678
rect 160296 50510 160416 50538
rect 160480 51190 160600 51218
rect 160192 49564 160244 49570
rect 160192 49506 160244 49512
rect 160100 49428 160152 49434
rect 160100 49370 160152 49376
rect 160008 45484 160060 45490
rect 160008 45426 160060 45432
rect 160204 44174 160232 49506
rect 160296 47462 160324 50510
rect 160376 50380 160428 50386
rect 160376 50322 160428 50328
rect 160284 47456 160336 47462
rect 160284 47398 160336 47404
rect 160204 44146 160324 44174
rect 159732 24200 159784 24206
rect 159732 24142 159784 24148
rect 159548 21412 159600 21418
rect 159548 21354 159600 21360
rect 160296 14482 160324 44146
rect 160388 18698 160416 50322
rect 160376 18692 160428 18698
rect 160376 18634 160428 18640
rect 160480 18630 160508 51190
rect 160664 51048 160692 51575
rect 160572 51020 160692 51048
rect 160572 50386 160600 51020
rect 160560 50380 160612 50386
rect 160560 50322 160612 50328
rect 160560 49360 160612 49366
rect 160560 49302 160612 49308
rect 160572 22846 160600 49302
rect 160756 46356 160784 51632
rect 160928 51614 160980 51620
rect 160836 49632 160888 49638
rect 160836 49574 160888 49580
rect 160848 47734 160876 49574
rect 160836 47728 160888 47734
rect 160836 47670 160888 47676
rect 160940 47410 160968 51614
rect 161032 49638 161060 51734
rect 161156 51711 161212 51720
rect 161112 51672 161164 51678
rect 161262 51660 161290 52020
rect 161354 51955 161382 52020
rect 161340 51946 161396 51955
rect 161446 51950 161474 52020
rect 161340 51881 161396 51890
rect 161434 51944 161486 51950
rect 161434 51886 161486 51892
rect 161386 51776 161442 51785
rect 161538 51728 161566 52020
rect 161630 51882 161658 52020
rect 161722 51921 161750 52020
rect 161814 51950 161842 52020
rect 161906 51950 161934 52020
rect 161802 51944 161854 51950
rect 161708 51912 161764 51921
rect 161618 51876 161670 51882
rect 161802 51886 161854 51892
rect 161894 51944 161946 51950
rect 161998 51921 162026 52020
rect 161894 51886 161946 51892
rect 161984 51912 162040 51921
rect 161708 51847 161764 51856
rect 161984 51847 162040 51856
rect 161618 51818 161670 51824
rect 162090 51796 162118 52020
rect 162044 51768 162118 51796
rect 161386 51711 161442 51720
rect 161112 51614 161164 51620
rect 161216 51632 161290 51660
rect 161020 49632 161072 49638
rect 161020 49574 161072 49580
rect 161124 49570 161152 51614
rect 161112 49564 161164 49570
rect 161112 49506 161164 49512
rect 161216 48482 161244 51632
rect 161296 51536 161348 51542
rect 161296 51478 161348 51484
rect 161204 48476 161256 48482
rect 161204 48418 161256 48424
rect 160940 47382 161060 47410
rect 160664 46328 160784 46356
rect 160560 22840 160612 22846
rect 160560 22782 160612 22788
rect 160664 22778 160692 46328
rect 160742 46064 160798 46073
rect 160742 45999 160798 46008
rect 160756 24177 160784 45999
rect 160928 43308 160980 43314
rect 160928 43250 160980 43256
rect 160742 24168 160798 24177
rect 160742 24103 160798 24112
rect 160652 22772 160704 22778
rect 160652 22714 160704 22720
rect 160468 18624 160520 18630
rect 160468 18566 160520 18572
rect 160284 14476 160336 14482
rect 160284 14418 160336 14424
rect 160940 5030 160968 43250
rect 161032 11762 161060 47382
rect 161308 43314 161336 51478
rect 161400 49366 161428 51711
rect 161492 51700 161566 51728
rect 161756 51740 161808 51746
rect 161492 50046 161520 51700
rect 161756 51682 161808 51688
rect 161768 51649 161796 51682
rect 161848 51672 161900 51678
rect 161754 51640 161810 51649
rect 161848 51614 161900 51620
rect 161754 51575 161810 51584
rect 161756 51536 161808 51542
rect 161756 51478 161808 51484
rect 161480 50040 161532 50046
rect 161480 49982 161532 49988
rect 161388 49360 161440 49366
rect 161388 49302 161440 49308
rect 161388 49020 161440 49026
rect 161388 48962 161440 48968
rect 161400 48929 161428 48962
rect 161768 48929 161796 51478
rect 161860 50182 161888 51614
rect 161940 51604 161992 51610
rect 161940 51546 161992 51552
rect 161848 50176 161900 50182
rect 161848 50118 161900 50124
rect 161952 49706 161980 51546
rect 161940 49700 161992 49706
rect 161940 49642 161992 49648
rect 161386 48920 161442 48929
rect 161754 48920 161810 48929
rect 161386 48855 161442 48864
rect 161572 48884 161624 48890
rect 161754 48855 161810 48864
rect 161572 48826 161624 48832
rect 161480 48612 161532 48618
rect 161480 48554 161532 48560
rect 161296 43308 161348 43314
rect 161296 43250 161348 43256
rect 161020 11756 161072 11762
rect 161020 11698 161072 11704
rect 161492 9042 161520 48554
rect 161480 9036 161532 9042
rect 161480 8978 161532 8984
rect 161584 7614 161612 48826
rect 162044 48754 162072 51768
rect 162182 51728 162210 52020
rect 162136 51700 162210 51728
rect 162136 48890 162164 51700
rect 162274 51660 162302 52020
rect 162366 51728 162394 52020
rect 162458 51921 162486 52020
rect 162444 51912 162500 51921
rect 162444 51847 162500 51856
rect 162550 51796 162578 52020
rect 162504 51768 162578 51796
rect 162366 51700 162440 51728
rect 162228 51632 162302 51660
rect 162124 48884 162176 48890
rect 162124 48826 162176 48832
rect 161756 48748 161808 48754
rect 161756 48690 161808 48696
rect 162032 48748 162084 48754
rect 162032 48690 162084 48696
rect 161664 48136 161716 48142
rect 161664 48078 161716 48084
rect 161676 13190 161704 48078
rect 161664 13184 161716 13190
rect 161664 13126 161716 13132
rect 161768 13122 161796 48690
rect 162124 48204 162176 48210
rect 162124 48146 162176 48152
rect 161848 46572 161900 46578
rect 161848 46514 161900 46520
rect 161860 15978 161888 46514
rect 161940 46164 161992 46170
rect 161940 46106 161992 46112
rect 161952 17270 161980 46106
rect 162030 45928 162086 45937
rect 162030 45863 162086 45872
rect 162044 19990 162072 45863
rect 162136 22914 162164 48146
rect 162228 46578 162256 51632
rect 162306 51504 162362 51513
rect 162306 51439 162362 51448
rect 162216 46572 162268 46578
rect 162216 46514 162268 46520
rect 162124 22908 162176 22914
rect 162124 22850 162176 22856
rect 162032 19984 162084 19990
rect 162032 19926 162084 19932
rect 161940 17264 161992 17270
rect 161940 17206 161992 17212
rect 161848 15972 161900 15978
rect 161848 15914 161900 15920
rect 161756 13116 161808 13122
rect 161756 13058 161808 13064
rect 161572 7608 161624 7614
rect 161572 7550 161624 7556
rect 160928 5024 160980 5030
rect 160928 4966 160980 4972
rect 162320 4894 162348 51439
rect 162412 48142 162440 51700
rect 162504 48210 162532 51768
rect 162642 51728 162670 52020
rect 162734 51921 162762 52020
rect 162720 51912 162776 51921
rect 162720 51847 162776 51856
rect 162826 51728 162854 52020
rect 162596 51700 162670 51728
rect 162780 51700 162854 51728
rect 162492 48204 162544 48210
rect 162492 48146 162544 48152
rect 162400 48136 162452 48142
rect 162400 48078 162452 48084
rect 162596 46170 162624 51700
rect 162780 51626 162808 51700
rect 162688 51598 162808 51626
rect 162918 51626 162946 52020
rect 163010 51950 163038 52020
rect 162998 51944 163050 51950
rect 162998 51886 163050 51892
rect 162996 51810 163052 51819
rect 162996 51745 163052 51754
rect 163102 51660 163130 52020
rect 163056 51632 163130 51660
rect 162918 51598 162992 51626
rect 162584 46164 162636 46170
rect 162584 46106 162636 46112
rect 162688 45554 162716 51598
rect 162766 51504 162822 51513
rect 162766 51439 162822 51448
rect 162780 48686 162808 51439
rect 162858 51096 162914 51105
rect 162858 51031 162860 51040
rect 162912 51031 162914 51040
rect 162860 51002 162912 51008
rect 162964 48929 162992 51598
rect 162950 48920 163006 48929
rect 162950 48855 163006 48864
rect 162768 48680 162820 48686
rect 162768 48622 162820 48628
rect 163056 48550 163084 51632
rect 163194 51592 163222 52020
rect 163148 51564 163222 51592
rect 163148 48793 163176 51564
rect 163286 51524 163314 52020
rect 163378 51882 163406 52020
rect 163470 51921 163498 52020
rect 163456 51912 163512 51921
rect 163366 51876 163418 51882
rect 163456 51847 163512 51856
rect 163366 51818 163418 51824
rect 163562 51814 163590 52020
rect 163654 51819 163682 52020
rect 163746 51950 163774 52020
rect 163734 51944 163786 51950
rect 163734 51886 163786 51892
rect 163550 51808 163602 51814
rect 163550 51750 163602 51756
rect 163640 51810 163696 51819
rect 163412 51740 163464 51746
rect 163640 51745 163696 51754
rect 163838 51728 163866 52020
rect 163930 51921 163958 52020
rect 164022 51950 164050 52020
rect 164010 51944 164062 51950
rect 163916 51912 163972 51921
rect 164114 51921 164142 52020
rect 164206 51950 164234 52020
rect 164194 51944 164246 51950
rect 164010 51886 164062 51892
rect 164100 51912 164156 51921
rect 163916 51847 163972 51856
rect 164194 51886 164246 51892
rect 164298 51882 164326 52020
rect 164390 51950 164418 52020
rect 164378 51944 164430 51950
rect 164482 51921 164510 52020
rect 164574 51950 164602 52020
rect 164562 51944 164614 51950
rect 164378 51886 164430 51892
rect 164468 51912 164524 51921
rect 164100 51847 164156 51856
rect 164286 51876 164338 51882
rect 164562 51886 164614 51892
rect 164468 51847 164524 51856
rect 164286 51818 164338 51824
rect 164516 51808 164568 51814
rect 163412 51682 163464 51688
rect 163792 51700 163866 51728
rect 164054 51776 164110 51785
rect 164666 51796 164694 52020
rect 164758 51921 164786 52020
rect 164744 51912 164800 51921
rect 164850 51882 164878 52020
rect 164942 51950 164970 52020
rect 165034 51950 165062 52020
rect 165126 51950 165154 52020
rect 164930 51944 164982 51950
rect 164930 51886 164982 51892
rect 165022 51944 165074 51950
rect 165022 51886 165074 51892
rect 165114 51944 165166 51950
rect 165114 51886 165166 51892
rect 164744 51847 164800 51856
rect 164838 51876 164890 51882
rect 164838 51818 164890 51824
rect 164976 51808 165028 51814
rect 164666 51768 164740 51796
rect 164516 51750 164568 51756
rect 164712 51762 164740 51768
rect 164882 51776 164938 51785
rect 164054 51711 164110 51720
rect 164424 51740 164476 51746
rect 163286 51496 163360 51524
rect 163332 48793 163360 51496
rect 163134 48784 163190 48793
rect 163318 48784 163374 48793
rect 163134 48719 163190 48728
rect 163228 48748 163280 48754
rect 163318 48719 163374 48728
rect 163228 48690 163280 48696
rect 163136 48680 163188 48686
rect 163136 48622 163188 48628
rect 163044 48544 163096 48550
rect 163044 48486 163096 48492
rect 162860 48204 162912 48210
rect 162860 48146 162912 48152
rect 162596 45526 162716 45554
rect 162596 24138 162624 45526
rect 162584 24132 162636 24138
rect 162584 24074 162636 24080
rect 162872 21622 162900 48146
rect 163148 48090 163176 48622
rect 163056 48062 163176 48090
rect 162952 45212 163004 45218
rect 162952 45154 163004 45160
rect 162860 21616 162912 21622
rect 162860 21558 162912 21564
rect 162492 6384 162544 6390
rect 162492 6326 162544 6332
rect 162308 4888 162360 4894
rect 162308 4830 162360 4836
rect 160100 4820 160152 4826
rect 160100 4762 160152 4768
rect 159456 3800 159508 3806
rect 159456 3742 159508 3748
rect 158168 3596 158220 3602
rect 158168 3538 158220 3544
rect 158076 3528 158128 3534
rect 158076 3470 158128 3476
rect 157984 3460 158036 3466
rect 157984 3402 158036 3408
rect 158904 3460 158956 3466
rect 158904 3402 158956 3408
rect 158916 480 158944 3402
rect 160112 480 160140 4762
rect 161296 3528 161348 3534
rect 161296 3470 161348 3476
rect 161308 480 161336 3470
rect 162504 480 162532 6326
rect 162964 6186 162992 45154
rect 163056 7682 163084 48062
rect 163240 47546 163268 48690
rect 163148 47518 163268 47546
rect 163148 8974 163176 47518
rect 163228 47456 163280 47462
rect 163228 47398 163280 47404
rect 163240 11830 163268 47398
rect 163424 46986 163452 51682
rect 163502 51640 163558 51649
rect 163792 51626 163820 51700
rect 163502 51575 163558 51584
rect 163700 51598 163820 51626
rect 163516 48634 163544 51575
rect 163596 51536 163648 51542
rect 163596 51478 163648 51484
rect 163608 48754 163636 51478
rect 163700 48754 163728 51598
rect 163964 51536 164016 51542
rect 163964 51478 164016 51484
rect 163596 48748 163648 48754
rect 163596 48690 163648 48696
rect 163688 48748 163740 48754
rect 163688 48690 163740 48696
rect 163516 48606 163728 48634
rect 163596 48476 163648 48482
rect 163596 48418 163648 48424
rect 163412 46980 163464 46986
rect 163412 46922 163464 46928
rect 163410 46880 163466 46889
rect 163410 46815 163466 46824
rect 163320 42900 163372 42906
rect 163320 42842 163372 42848
rect 163332 17338 163360 42842
rect 163424 21554 163452 46815
rect 163608 24410 163636 48418
rect 163596 24404 163648 24410
rect 163596 24346 163648 24352
rect 163412 21548 163464 21554
rect 163412 21490 163464 21496
rect 163320 17332 163372 17338
rect 163320 17274 163372 17280
rect 163228 11824 163280 11830
rect 163228 11766 163280 11772
rect 163136 8968 163188 8974
rect 163136 8910 163188 8916
rect 163044 7676 163096 7682
rect 163044 7618 163096 7624
rect 163700 6914 163728 48606
rect 163976 42906 164004 51478
rect 164068 45218 164096 51711
rect 164424 51682 164476 51688
rect 164148 51672 164200 51678
rect 164148 51614 164200 51620
rect 164160 47462 164188 51614
rect 164240 51604 164292 51610
rect 164240 51546 164292 51552
rect 164252 48210 164280 51546
rect 164436 48657 164464 51682
rect 164422 48648 164478 48657
rect 164422 48583 164478 48592
rect 164528 48482 164556 51750
rect 164712 51734 164786 51762
rect 164608 51672 164660 51678
rect 164608 51614 164660 51620
rect 164516 48476 164568 48482
rect 164516 48418 164568 48424
rect 164424 48340 164476 48346
rect 164424 48282 164476 48288
rect 164240 48204 164292 48210
rect 164240 48146 164292 48152
rect 164148 47456 164200 47462
rect 164148 47398 164200 47404
rect 164056 45212 164108 45218
rect 164056 45154 164108 45160
rect 163964 42900 164016 42906
rect 163964 42842 164016 42848
rect 164436 7818 164464 48282
rect 164620 48192 164648 51614
rect 164758 51524 164786 51734
rect 164976 51750 165028 51756
rect 164882 51711 164938 51720
rect 164758 51496 164832 51524
rect 164698 51368 164754 51377
rect 164698 51303 164754 51312
rect 164528 48164 164648 48192
rect 164528 13258 164556 48164
rect 164712 48090 164740 51303
rect 164804 48482 164832 51496
rect 164792 48476 164844 48482
rect 164792 48418 164844 48424
rect 164792 48204 164844 48210
rect 164792 48146 164844 48152
rect 164620 48062 164740 48090
rect 164620 17406 164648 48062
rect 164700 47932 164752 47938
rect 164700 47874 164752 47880
rect 164712 18834 164740 47874
rect 164700 18828 164752 18834
rect 164700 18770 164752 18776
rect 164804 18766 164832 48146
rect 164896 20058 164924 51711
rect 164988 48346 165016 51750
rect 165068 51740 165120 51746
rect 165068 51682 165120 51688
rect 165080 51649 165108 51682
rect 165218 51660 165246 52020
rect 165310 51785 165338 52020
rect 165402 51955 165430 52020
rect 165388 51946 165444 51955
rect 165494 51950 165522 52020
rect 165586 51955 165614 52020
rect 165388 51881 165444 51890
rect 165482 51944 165534 51950
rect 165482 51886 165534 51892
rect 165572 51946 165628 51955
rect 165678 51950 165706 52020
rect 165770 51950 165798 52020
rect 165862 51955 165890 52020
rect 165572 51881 165628 51890
rect 165666 51944 165718 51950
rect 165666 51886 165718 51892
rect 165758 51944 165810 51950
rect 165758 51886 165810 51892
rect 165848 51946 165904 51955
rect 165954 51950 165982 52020
rect 166046 51950 166074 52020
rect 165848 51881 165904 51890
rect 165942 51944 165994 51950
rect 165942 51886 165994 51892
rect 166034 51944 166086 51950
rect 166138 51921 166166 52020
rect 166230 51950 166258 52020
rect 166322 51950 166350 52020
rect 166218 51944 166270 51950
rect 166034 51886 166086 51892
rect 166124 51912 166180 51921
rect 166218 51886 166270 51892
rect 166310 51944 166362 51950
rect 166310 51886 166362 51892
rect 166414 51882 166442 52020
rect 166124 51847 166180 51856
rect 166402 51876 166454 51882
rect 166402 51818 166454 51824
rect 166506 51814 166534 52020
rect 166598 51882 166626 52020
rect 166690 51955 166718 52020
rect 166676 51946 166732 51955
rect 166586 51876 166638 51882
rect 166676 51881 166732 51890
rect 166586 51818 166638 51824
rect 165528 51808 165580 51814
rect 165296 51776 165352 51785
rect 165528 51750 165580 51756
rect 166494 51808 166546 51814
rect 166782 51785 166810 52020
rect 166494 51750 166546 51756
rect 166768 51776 166824 51785
rect 165296 51711 165352 51720
rect 165066 51640 165122 51649
rect 165218 51632 165384 51660
rect 165066 51575 165122 51584
rect 165068 51536 165120 51542
rect 165068 51478 165120 51484
rect 165250 51504 165306 51513
rect 164976 48340 165028 48346
rect 164976 48282 165028 48288
rect 165080 48226 165108 51478
rect 165250 51439 165306 51448
rect 165158 51368 165214 51377
rect 165158 51303 165214 51312
rect 164988 48198 165108 48226
rect 164988 24478 165016 48198
rect 165068 48136 165120 48142
rect 165068 48078 165120 48084
rect 164976 24472 165028 24478
rect 164976 24414 165028 24420
rect 164884 20052 164936 20058
rect 164884 19994 164936 20000
rect 164792 18760 164844 18766
rect 164792 18702 164844 18708
rect 164608 17400 164660 17406
rect 164608 17342 164660 17348
rect 164516 13252 164568 13258
rect 164516 13194 164568 13200
rect 164424 7812 164476 7818
rect 164424 7754 164476 7760
rect 163608 6886 163728 6914
rect 162952 6180 163004 6186
rect 162952 6122 163004 6128
rect 163608 4962 163636 6886
rect 165080 6254 165108 48078
rect 165172 42794 165200 51303
rect 165264 48618 165292 51439
rect 165252 48612 165304 48618
rect 165252 48554 165304 48560
rect 165252 48476 165304 48482
rect 165252 48418 165304 48424
rect 165264 47580 165292 48418
rect 165356 48142 165384 51632
rect 165434 51640 165490 51649
rect 165434 51575 165490 51584
rect 165344 48136 165396 48142
rect 165344 48078 165396 48084
rect 165448 47938 165476 51575
rect 165540 49094 165568 51750
rect 165896 51740 165948 51746
rect 165896 51682 165948 51688
rect 165988 51740 166040 51746
rect 165988 51682 166040 51688
rect 166172 51740 166224 51746
rect 166172 51682 166224 51688
rect 166264 51740 166316 51746
rect 166768 51711 166824 51720
rect 166264 51682 166316 51688
rect 165712 51672 165764 51678
rect 165712 51614 165764 51620
rect 165620 51468 165672 51474
rect 165620 51410 165672 51416
rect 165528 49088 165580 49094
rect 165528 49030 165580 49036
rect 165632 48210 165660 51410
rect 165724 49473 165752 51614
rect 165802 51368 165858 51377
rect 165802 51303 165858 51312
rect 165710 49464 165766 49473
rect 165710 49399 165766 49408
rect 165816 49162 165844 51303
rect 165908 49473 165936 51682
rect 165894 49464 165950 49473
rect 165894 49399 165950 49408
rect 165804 49156 165856 49162
rect 165804 49098 165856 49104
rect 165620 48204 165672 48210
rect 165620 48146 165672 48152
rect 165436 47932 165488 47938
rect 165436 47874 165488 47880
rect 165264 47552 165476 47580
rect 165172 42766 165292 42794
rect 165264 24546 165292 42766
rect 165252 24540 165304 24546
rect 165252 24482 165304 24488
rect 165448 7750 165476 47552
rect 166000 42794 166028 51682
rect 166080 51604 166132 51610
rect 166080 51546 166132 51552
rect 165816 42766 166028 42794
rect 165816 11898 165844 42766
rect 165988 42628 166040 42634
rect 165988 42570 166040 42576
rect 165896 42492 165948 42498
rect 165896 42434 165948 42440
rect 165908 14618 165936 42434
rect 165896 14612 165948 14618
rect 165896 14554 165948 14560
rect 166000 14550 166028 42570
rect 166092 20126 166120 51546
rect 166184 21690 166212 51682
rect 166276 42634 166304 51682
rect 166356 51672 166408 51678
rect 166874 51660 166902 52020
rect 166966 51887 166994 52020
rect 166952 51878 167008 51887
rect 167058 51882 167086 52020
rect 167150 51950 167178 52020
rect 167138 51944 167190 51950
rect 167138 51886 167190 51892
rect 167242 51882 167270 52020
rect 167334 51950 167362 52020
rect 167426 51950 167454 52020
rect 167322 51944 167374 51950
rect 167322 51886 167374 51892
rect 167414 51944 167466 51950
rect 167414 51886 167466 51892
rect 167518 51882 167546 52020
rect 167610 51955 167638 52020
rect 167596 51946 167652 51955
rect 166952 51813 167008 51822
rect 167046 51876 167098 51882
rect 167046 51818 167098 51824
rect 167230 51876 167282 51882
rect 167230 51818 167282 51824
rect 167506 51876 167558 51882
rect 167596 51881 167652 51890
rect 167506 51818 167558 51824
rect 167414 51808 167466 51814
rect 167274 51776 167330 51785
rect 167000 51740 167052 51746
rect 167000 51682 167052 51688
rect 167184 51740 167236 51746
rect 167274 51711 167330 51720
rect 167412 51776 167414 51785
rect 167466 51776 167468 51785
rect 167702 51762 167730 52020
rect 167794 51955 167822 52020
rect 167780 51946 167836 51955
rect 167886 51950 167914 52020
rect 167780 51881 167836 51890
rect 167874 51944 167926 51950
rect 167874 51886 167926 51892
rect 167978 51887 168006 52020
rect 168070 51950 168098 52020
rect 168162 51950 168190 52020
rect 168058 51944 168110 51950
rect 167964 51878 168020 51887
rect 168058 51886 168110 51892
rect 168150 51944 168202 51950
rect 168150 51886 168202 51892
rect 168254 51882 168282 52020
rect 167964 51813 168020 51822
rect 168242 51876 168294 51882
rect 168242 51818 168294 51824
rect 167412 51711 167468 51720
rect 167564 51734 167730 51762
rect 168012 51740 168064 51746
rect 167184 51682 167236 51688
rect 166356 51614 166408 51620
rect 166722 51640 166778 51649
rect 166368 46170 166396 51614
rect 166722 51575 166778 51584
rect 166828 51632 166902 51660
rect 166630 51504 166686 51513
rect 166448 51468 166500 51474
rect 166630 51439 166686 51448
rect 166448 51410 166500 51416
rect 166356 46164 166408 46170
rect 166356 46106 166408 46112
rect 166460 42794 166488 51410
rect 166368 42766 166488 42794
rect 166264 42628 166316 42634
rect 166264 42570 166316 42576
rect 166264 41676 166316 41682
rect 166264 41618 166316 41624
rect 166276 22982 166304 41618
rect 166264 22976 166316 22982
rect 166264 22918 166316 22924
rect 166172 21684 166224 21690
rect 166172 21626 166224 21632
rect 166080 20120 166132 20126
rect 166080 20062 166132 20068
rect 165988 14544 166040 14550
rect 165988 14486 166040 14492
rect 165804 11892 165856 11898
rect 165804 11834 165856 11840
rect 166080 11824 166132 11830
rect 166080 11766 166132 11772
rect 165436 7744 165488 7750
rect 165436 7686 165488 7692
rect 165068 6248 165120 6254
rect 163686 6216 163742 6225
rect 165068 6190 165120 6196
rect 163686 6151 163742 6160
rect 163596 4956 163648 4962
rect 163596 4898 163648 4904
rect 163700 480 163728 6151
rect 164884 3596 164936 3602
rect 164884 3538 164936 3544
rect 164896 480 164924 3538
rect 166092 480 166120 11766
rect 166368 7886 166396 42766
rect 166644 41682 166672 51439
rect 166736 47598 166764 51575
rect 166724 47592 166776 47598
rect 166724 47534 166776 47540
rect 166722 47424 166778 47433
rect 166722 47359 166778 47368
rect 166632 41676 166684 41682
rect 166632 41618 166684 41624
rect 166736 41414 166764 47359
rect 166828 42498 166856 51632
rect 166908 51536 166960 51542
rect 166908 51478 166960 51484
rect 166920 51270 166948 51478
rect 166908 51264 166960 51270
rect 166908 51206 166960 51212
rect 167012 49502 167040 51682
rect 167092 51672 167144 51678
rect 167092 51614 167144 51620
rect 167000 49496 167052 49502
rect 167000 49438 167052 49444
rect 167104 47433 167132 51614
rect 167090 47424 167146 47433
rect 167090 47359 167146 47368
rect 167000 47320 167052 47326
rect 167000 47262 167052 47268
rect 166908 46164 166960 46170
rect 166908 46106 166960 46112
rect 166816 42492 166868 42498
rect 166816 42434 166868 42440
rect 166460 41386 166764 41414
rect 166460 10334 166488 41386
rect 166920 24682 166948 46106
rect 167012 41414 167040 47262
rect 167196 46209 167224 51682
rect 167288 47705 167316 51711
rect 167368 51672 167420 51678
rect 167368 51614 167420 51620
rect 167460 51672 167512 51678
rect 167460 51614 167512 51620
rect 167274 47696 167330 47705
rect 167274 47631 167330 47640
rect 167276 47592 167328 47598
rect 167380 47569 167408 51614
rect 167472 49230 167500 51614
rect 167460 49224 167512 49230
rect 167460 49166 167512 49172
rect 167276 47534 167328 47540
rect 167366 47560 167422 47569
rect 167182 46200 167238 46209
rect 167182 46135 167238 46144
rect 167012 41386 167224 41414
rect 166908 24676 166960 24682
rect 166908 24618 166960 24624
rect 167196 10470 167224 41386
rect 167288 11966 167316 47534
rect 167366 47495 167422 47504
rect 167460 47456 167512 47462
rect 167460 47398 167512 47404
rect 167368 46844 167420 46850
rect 167368 46786 167420 46792
rect 167380 16182 167408 46786
rect 167368 16176 167420 16182
rect 167368 16118 167420 16124
rect 167472 16114 167500 47398
rect 167460 16108 167512 16114
rect 167460 16050 167512 16056
rect 167564 16046 167592 51734
rect 168346 51728 168374 52020
rect 168012 51682 168064 51688
rect 168300 51700 168374 51728
rect 168438 51728 168466 52020
rect 168530 51796 168558 52020
rect 168622 51955 168650 52020
rect 168608 51946 168664 51955
rect 168608 51881 168664 51890
rect 168714 51814 168742 52020
rect 168806 51921 168834 52020
rect 168792 51912 168848 51921
rect 168898 51882 168926 52020
rect 168792 51847 168848 51856
rect 168886 51876 168938 51882
rect 168886 51818 168938 51824
rect 168702 51808 168754 51814
rect 168530 51768 168604 51796
rect 168438 51700 168512 51728
rect 167734 51640 167790 51649
rect 167656 51598 167734 51626
rect 167656 47598 167684 51598
rect 167734 51575 167790 51584
rect 167828 51604 167880 51610
rect 167828 51546 167880 51552
rect 167734 51504 167790 51513
rect 167734 51439 167790 51448
rect 167644 47592 167696 47598
rect 167644 47534 167696 47540
rect 167748 47462 167776 51439
rect 167736 47456 167788 47462
rect 167736 47398 167788 47404
rect 167840 47326 167868 51546
rect 167828 47320 167880 47326
rect 167828 47262 167880 47268
rect 168024 46866 168052 51682
rect 168104 51672 168156 51678
rect 168104 51614 168156 51620
rect 167656 46838 168052 46866
rect 168116 46850 168144 51614
rect 168196 51604 168248 51610
rect 168196 51546 168248 51552
rect 168104 46844 168156 46850
rect 167656 20194 167684 46838
rect 168104 46786 168156 46792
rect 168208 45898 168236 51546
rect 168300 47666 168328 51700
rect 168380 51604 168432 51610
rect 168380 51546 168432 51552
rect 168288 47660 168340 47666
rect 168288 47602 168340 47608
rect 168392 46374 168420 51546
rect 168484 49978 168512 51700
rect 168472 49972 168524 49978
rect 168472 49914 168524 49920
rect 168472 49224 168524 49230
rect 168472 49166 168524 49172
rect 168380 46368 168432 46374
rect 168380 46310 168432 46316
rect 168484 46186 168512 49166
rect 168576 48113 168604 51768
rect 168990 51785 169018 52020
rect 168702 51750 168754 51756
rect 168976 51776 169032 51785
rect 168840 51740 168892 51746
rect 168976 51711 169032 51720
rect 168840 51682 168892 51688
rect 168748 51672 168800 51678
rect 168654 51640 168710 51649
rect 168748 51614 168800 51620
rect 168654 51575 168710 51584
rect 168562 48104 168618 48113
rect 168562 48039 168618 48048
rect 168564 46980 168616 46986
rect 168564 46922 168616 46928
rect 168300 46158 168512 46186
rect 167736 45892 167788 45898
rect 167736 45834 167788 45840
rect 168196 45892 168248 45898
rect 168196 45834 168248 45840
rect 167644 20188 167696 20194
rect 167644 20130 167696 20136
rect 167552 16040 167604 16046
rect 167552 15982 167604 15988
rect 167276 11960 167328 11966
rect 167276 11902 167328 11908
rect 167184 10464 167236 10470
rect 167184 10406 167236 10412
rect 166448 10328 166500 10334
rect 166448 10270 166500 10276
rect 166356 7880 166408 7886
rect 166356 7822 166408 7828
rect 167748 6322 167776 45834
rect 167826 45792 167882 45801
rect 167826 45727 167882 45736
rect 167840 10402 167868 45727
rect 168300 24750 168328 46158
rect 168380 45076 168432 45082
rect 168380 45018 168432 45024
rect 168288 24744 168340 24750
rect 168288 24686 168340 24692
rect 167828 10396 167880 10402
rect 167828 10338 167880 10344
rect 167736 6316 167788 6322
rect 167736 6258 167788 6264
rect 167182 4856 167238 4865
rect 167182 4791 167238 4800
rect 167196 480 167224 4791
rect 168392 3466 168420 45018
rect 168576 10538 168604 46922
rect 168668 13326 168696 51575
rect 168760 51513 168788 51614
rect 168746 51504 168802 51513
rect 168746 51439 168802 51448
rect 168852 48940 168880 51682
rect 169082 51660 169110 52020
rect 169174 51950 169202 52020
rect 169162 51944 169214 51950
rect 169162 51886 169214 51892
rect 169266 51796 169294 52020
rect 169358 51950 169386 52020
rect 169346 51944 169398 51950
rect 169346 51886 169398 51892
rect 168760 48912 168880 48940
rect 169036 51632 169110 51660
rect 169220 51768 169294 51796
rect 168760 14686 168788 48912
rect 169036 48872 169064 51632
rect 168852 48844 169064 48872
rect 168852 16250 168880 48844
rect 169024 48748 169076 48754
rect 169024 48690 169076 48696
rect 168932 46028 168984 46034
rect 168932 45970 168984 45976
rect 168944 20262 168972 45970
rect 169036 24002 169064 48690
rect 169116 47932 169168 47938
rect 169116 47874 169168 47880
rect 169024 23996 169076 24002
rect 169024 23938 169076 23944
rect 169128 21758 169156 47874
rect 169220 46986 169248 51768
rect 169300 51672 169352 51678
rect 169450 51660 169478 52020
rect 169542 51762 169570 52020
rect 169634 51950 169662 52020
rect 169726 51955 169754 52020
rect 169622 51944 169674 51950
rect 169622 51886 169674 51892
rect 169712 51946 169768 51955
rect 169712 51881 169768 51890
rect 169818 51762 169846 52020
rect 169910 51882 169938 52020
rect 169898 51876 169950 51882
rect 169898 51818 169950 51824
rect 169542 51734 169708 51762
rect 169818 51734 169892 51762
rect 169576 51672 169628 51678
rect 169450 51632 169524 51660
rect 169300 51614 169352 51620
rect 169208 46980 169260 46986
rect 169208 46922 169260 46928
rect 169312 45554 169340 51614
rect 169496 48754 169524 51632
rect 169576 51614 169628 51620
rect 169484 48748 169536 48754
rect 169484 48690 169536 48696
rect 169588 46034 169616 51614
rect 169680 50368 169708 51734
rect 169864 51626 169892 51734
rect 169864 51598 169938 51626
rect 169758 51504 169814 51513
rect 169910 51490 169938 51598
rect 170002 51592 170030 52020
rect 170094 51785 170122 52020
rect 170186 51921 170214 52020
rect 170172 51912 170228 51921
rect 170172 51847 170228 51856
rect 170080 51776 170136 51785
rect 170278 51728 170306 52020
rect 170370 51882 170398 52020
rect 170358 51876 170410 51882
rect 170358 51818 170410 51824
rect 170462 51728 170490 52020
rect 170554 51762 170582 52020
rect 170646 51921 170674 52020
rect 170738 51950 170766 52020
rect 170726 51944 170778 51950
rect 170632 51912 170688 51921
rect 170726 51886 170778 51892
rect 170632 51847 170688 51856
rect 170830 51796 170858 52020
rect 170922 51882 170950 52020
rect 171014 51882 171042 52020
rect 170910 51876 170962 51882
rect 170910 51818 170962 51824
rect 171002 51876 171054 51882
rect 171002 51818 171054 51824
rect 170784 51785 170858 51796
rect 170770 51776 170858 51785
rect 170554 51746 170628 51762
rect 170554 51740 170640 51746
rect 170554 51734 170588 51740
rect 170080 51711 170136 51720
rect 170232 51700 170306 51728
rect 170370 51700 170490 51728
rect 170128 51672 170180 51678
rect 170126 51640 170128 51649
rect 170180 51640 170182 51649
rect 170002 51564 170076 51592
rect 170126 51575 170182 51584
rect 169758 51439 169814 51448
rect 169864 51462 169938 51490
rect 169772 51406 169800 51439
rect 169760 51400 169812 51406
rect 169760 51342 169812 51348
rect 169680 50340 169800 50368
rect 169666 50280 169722 50289
rect 169666 50215 169722 50224
rect 169680 47802 169708 50215
rect 169772 47938 169800 50340
rect 169760 47932 169812 47938
rect 169760 47874 169812 47880
rect 169668 47796 169720 47802
rect 169668 47738 169720 47744
rect 169760 46164 169812 46170
rect 169760 46106 169812 46112
rect 169576 46028 169628 46034
rect 169576 45970 169628 45976
rect 169220 45526 169340 45554
rect 169116 21752 169168 21758
rect 169116 21694 169168 21700
rect 168932 20256 168984 20262
rect 168932 20198 168984 20204
rect 168840 16244 168892 16250
rect 168840 16186 168892 16192
rect 168748 14680 168800 14686
rect 168748 14622 168800 14628
rect 168656 13320 168708 13326
rect 168656 13262 168708 13268
rect 168564 10532 168616 10538
rect 168564 10474 168616 10480
rect 169220 9110 169248 45526
rect 169772 36582 169800 46106
rect 169760 36576 169812 36582
rect 169760 36518 169812 36524
rect 169760 33788 169812 33794
rect 169760 33730 169812 33736
rect 169772 16574 169800 33730
rect 169864 20534 169892 51462
rect 169942 51368 169998 51377
rect 169942 51303 169998 51312
rect 169956 36650 169984 51303
rect 170048 46170 170076 51564
rect 170128 51536 170180 51542
rect 170128 51478 170180 51484
rect 170140 51105 170168 51478
rect 170126 51096 170182 51105
rect 170126 51031 170182 51040
rect 170036 46164 170088 46170
rect 170036 46106 170088 46112
rect 170128 46096 170180 46102
rect 170128 46038 170180 46044
rect 170036 46028 170088 46034
rect 170036 45970 170088 45976
rect 170048 40050 170076 45970
rect 170036 40044 170088 40050
rect 170036 39986 170088 39992
rect 170140 39914 170168 46038
rect 170232 39982 170260 51700
rect 170370 51626 170398 51700
rect 170826 51768 170858 51776
rect 171106 51728 171134 52020
rect 170770 51711 170826 51720
rect 170588 51682 170640 51688
rect 171060 51700 171134 51728
rect 170864 51672 170916 51678
rect 170586 51640 170642 51649
rect 170370 51598 170444 51626
rect 170312 51536 170364 51542
rect 170312 51478 170364 51484
rect 170324 48793 170352 51478
rect 170310 48784 170366 48793
rect 170310 48719 170366 48728
rect 170310 48648 170366 48657
rect 170310 48583 170366 48592
rect 170324 41410 170352 48583
rect 170312 41404 170364 41410
rect 170312 41346 170364 41352
rect 170416 41138 170444 51598
rect 170496 51604 170548 51610
rect 170586 51575 170642 51584
rect 170784 51620 170864 51626
rect 170784 51614 170916 51620
rect 170784 51598 170904 51614
rect 170496 51546 170548 51552
rect 170508 42090 170536 51546
rect 170496 42084 170548 42090
rect 170496 42026 170548 42032
rect 170600 42022 170628 51575
rect 170680 51536 170732 51542
rect 170680 51478 170732 51484
rect 170692 46034 170720 51478
rect 170784 50289 170812 51598
rect 170956 51536 171008 51542
rect 170862 51504 170918 51513
rect 170956 51478 171008 51484
rect 170862 51439 170918 51448
rect 170770 50280 170826 50289
rect 170770 50215 170826 50224
rect 170876 48314 170904 51439
rect 170968 50930 170996 51478
rect 170956 50924 171008 50930
rect 170956 50866 171008 50872
rect 171060 50833 171088 51700
rect 171198 51660 171226 52020
rect 171290 51921 171318 52020
rect 171276 51912 171332 51921
rect 171276 51847 171332 51856
rect 171152 51632 171226 51660
rect 171046 50824 171102 50833
rect 171046 50759 171102 50768
rect 170876 48286 170996 48314
rect 170968 46102 170996 48286
rect 170956 46096 171008 46102
rect 170956 46038 171008 46044
rect 171152 46034 171180 51632
rect 171382 51592 171410 52020
rect 171474 51660 171502 52020
rect 171566 51762 171594 52020
rect 171658 51921 171686 52020
rect 171644 51912 171700 51921
rect 171644 51847 171700 51856
rect 171750 51762 171778 52020
rect 171566 51734 171640 51762
rect 171474 51632 171548 51660
rect 171612 51649 171640 51734
rect 171704 51734 171778 51762
rect 171336 51564 171410 51592
rect 171230 51504 171286 51513
rect 171230 51439 171286 51448
rect 171244 50182 171272 51439
rect 171232 50176 171284 50182
rect 171232 50118 171284 50124
rect 171336 48314 171364 51564
rect 171414 51368 171470 51377
rect 171414 51303 171470 51312
rect 171520 51320 171548 51632
rect 171598 51640 171654 51649
rect 171598 51575 171654 51584
rect 171244 48286 171364 48314
rect 170680 46028 170732 46034
rect 170680 45970 170732 45976
rect 171140 46028 171192 46034
rect 171140 45970 171192 45976
rect 171140 44192 171192 44198
rect 171140 44134 171192 44140
rect 170588 42016 170640 42022
rect 170588 41958 170640 41964
rect 170404 41132 170456 41138
rect 170404 41074 170456 41080
rect 170220 39976 170272 39982
rect 170220 39918 170272 39924
rect 170128 39908 170180 39914
rect 170128 39850 170180 39856
rect 169944 36644 169996 36650
rect 169944 36586 169996 36592
rect 169852 20528 169904 20534
rect 169852 20470 169904 20476
rect 171152 16574 171180 44134
rect 171244 39846 171272 48286
rect 171324 46368 171376 46374
rect 171324 46310 171376 46316
rect 171232 39840 171284 39846
rect 171232 39782 171284 39788
rect 171336 39778 171364 46310
rect 171324 39772 171376 39778
rect 171324 39714 171376 39720
rect 171428 39710 171456 51303
rect 171520 51292 171640 51320
rect 171506 51232 171562 51241
rect 171506 51167 171562 51176
rect 171520 46374 171548 51167
rect 171508 46368 171560 46374
rect 171508 46310 171560 46316
rect 171508 46164 171560 46170
rect 171508 46106 171560 46112
rect 171520 41274 171548 46106
rect 171612 41342 171640 51292
rect 171704 46170 171732 51734
rect 171842 51660 171870 52020
rect 171934 51762 171962 52020
rect 172026 51950 172054 52020
rect 172014 51944 172066 51950
rect 172014 51886 172066 51892
rect 172118 51887 172146 52020
rect 172104 51878 172160 51887
rect 172104 51813 172160 51822
rect 172210 51762 172238 52020
rect 172302 51882 172330 52020
rect 172290 51876 172342 51882
rect 172290 51818 172342 51824
rect 172394 51762 172422 52020
rect 171934 51734 172100 51762
rect 172210 51734 172284 51762
rect 171796 51632 171870 51660
rect 171968 51672 172020 51678
rect 171796 50862 171824 51632
rect 171968 51614 172020 51620
rect 171876 51468 171928 51474
rect 171876 51410 171928 51416
rect 171888 51134 171916 51410
rect 171876 51128 171928 51134
rect 171876 51070 171928 51076
rect 171784 50856 171836 50862
rect 171784 50798 171836 50804
rect 171876 50176 171928 50182
rect 171876 50118 171928 50124
rect 171692 46164 171744 46170
rect 171692 46106 171744 46112
rect 171692 46028 171744 46034
rect 171692 45970 171744 45976
rect 171704 41954 171732 45970
rect 171692 41948 171744 41954
rect 171692 41890 171744 41896
rect 171888 41414 171916 50118
rect 171980 49230 172008 51614
rect 171968 49224 172020 49230
rect 171968 49166 172020 49172
rect 172072 48550 172100 51734
rect 172152 51672 172204 51678
rect 172152 51614 172204 51620
rect 172164 49502 172192 51614
rect 172256 50930 172284 51734
rect 172348 51734 172422 51762
rect 172348 51513 172376 51734
rect 172486 51660 172514 52020
rect 172578 51762 172606 52020
rect 172670 51887 172698 52020
rect 172656 51878 172712 51887
rect 172656 51813 172712 51822
rect 172762 51762 172790 52020
rect 172578 51734 172652 51762
rect 172440 51632 172514 51660
rect 172334 51504 172390 51513
rect 172334 51439 172390 51448
rect 172334 51368 172390 51377
rect 172334 51303 172390 51312
rect 172244 50924 172296 50930
rect 172244 50866 172296 50872
rect 172348 50386 172376 51303
rect 172336 50380 172388 50386
rect 172336 50322 172388 50328
rect 172152 49496 172204 49502
rect 172440 49473 172468 51632
rect 172518 51504 172574 51513
rect 172518 51439 172574 51448
rect 172152 49438 172204 49444
rect 172426 49464 172482 49473
rect 172426 49399 172482 49408
rect 172532 49366 172560 51439
rect 172520 49360 172572 49366
rect 172520 49302 172572 49308
rect 172150 48920 172206 48929
rect 172150 48855 172206 48864
rect 172060 48544 172112 48550
rect 172060 48486 172112 48492
rect 171704 41386 171916 41414
rect 171600 41336 171652 41342
rect 171600 41278 171652 41284
rect 171508 41268 171560 41274
rect 171508 41210 171560 41216
rect 171704 41070 171732 41386
rect 172164 41206 172192 48855
rect 172520 41472 172572 41478
rect 172520 41414 172572 41420
rect 172152 41200 172204 41206
rect 172152 41142 172204 41148
rect 171692 41064 171744 41070
rect 171692 41006 171744 41012
rect 171416 39704 171468 39710
rect 171416 39646 171468 39652
rect 172532 38622 172560 41414
rect 172520 38616 172572 38622
rect 172520 38558 172572 38564
rect 172624 38554 172652 51734
rect 172716 51734 172790 51762
rect 172716 49298 172744 51734
rect 172854 51660 172882 52020
rect 172946 51814 172974 52020
rect 173038 51814 173066 52020
rect 173130 51921 173158 52020
rect 173116 51912 173172 51921
rect 173116 51847 173172 51856
rect 172934 51808 172986 51814
rect 172934 51750 172986 51756
rect 173026 51808 173078 51814
rect 173026 51750 173078 51756
rect 173222 51762 173250 52020
rect 173314 51882 173342 52020
rect 173302 51876 173354 51882
rect 173302 51818 173354 51824
rect 173406 51814 173434 52020
rect 173394 51808 173446 51814
rect 173222 51734 173296 51762
rect 173394 51750 173446 51756
rect 172980 51672 173032 51678
rect 172854 51632 172928 51660
rect 172794 51504 172850 51513
rect 172794 51439 172850 51448
rect 172704 49292 172756 49298
rect 172704 49234 172756 49240
rect 172808 49094 172836 51439
rect 172900 50561 172928 51632
rect 172980 51614 173032 51620
rect 173072 51672 173124 51678
rect 173072 51614 173124 51620
rect 173164 51672 173216 51678
rect 173164 51614 173216 51620
rect 172886 50552 172942 50561
rect 172886 50487 172942 50496
rect 172796 49088 172848 49094
rect 172796 49030 172848 49036
rect 172992 46918 173020 51614
rect 173084 51377 173112 51614
rect 173070 51368 173126 51377
rect 173070 51303 173126 51312
rect 173176 49570 173204 51614
rect 173164 49564 173216 49570
rect 173164 49506 173216 49512
rect 173268 48958 173296 51734
rect 173348 51672 173400 51678
rect 173498 51660 173526 52020
rect 173590 51814 173618 52020
rect 173578 51808 173630 51814
rect 173578 51750 173630 51756
rect 173682 51762 173710 52020
rect 173774 51921 173802 52020
rect 173760 51912 173816 51921
rect 173760 51847 173816 51856
rect 173866 51785 173894 52020
rect 173958 51921 173986 52020
rect 173944 51912 174000 51921
rect 173944 51847 174000 51856
rect 173852 51776 173908 51785
rect 173682 51734 173756 51762
rect 173624 51672 173676 51678
rect 173498 51632 173572 51660
rect 173348 51614 173400 51620
rect 173256 48952 173308 48958
rect 173256 48894 173308 48900
rect 173256 47592 173308 47598
rect 173162 47560 173218 47569
rect 173256 47534 173308 47540
rect 173162 47495 173218 47504
rect 172980 46912 173032 46918
rect 172980 46854 173032 46860
rect 172612 38548 172664 38554
rect 172612 38490 172664 38496
rect 169772 16546 170352 16574
rect 171152 16546 172008 16574
rect 169208 9104 169260 9110
rect 169208 9046 169260 9052
rect 168472 4140 168524 4146
rect 168472 4082 168524 4088
rect 168380 3460 168432 3466
rect 168380 3402 168432 3408
rect 168484 2122 168512 4082
rect 169576 3460 169628 3466
rect 169576 3402 169628 3408
rect 168392 2094 168512 2122
rect 168392 480 168420 2094
rect 169588 480 169616 3402
rect 156574 354 156686 480
rect 156156 326 156686 354
rect 156574 -960 156686 326
rect 157770 -960 157882 480
rect 158874 -960 158986 480
rect 160070 -960 160182 480
rect 161266 -960 161378 480
rect 162462 -960 162574 480
rect 163658 -960 163770 480
rect 164854 -960 164966 480
rect 166050 -960 166162 480
rect 167154 -960 167266 480
rect 168350 -960 168462 480
rect 169546 -960 169658 480
rect 170324 354 170352 16546
rect 171980 480 172008 16546
rect 173176 4146 173204 47495
rect 173164 4140 173216 4146
rect 173164 4082 173216 4088
rect 173268 3874 173296 47534
rect 173360 41478 173388 51614
rect 173440 51400 173492 51406
rect 173440 51342 173492 51348
rect 173452 51066 173480 51342
rect 173440 51060 173492 51066
rect 173440 51002 173492 51008
rect 173544 46850 173572 51632
rect 173624 51614 173676 51620
rect 173728 51626 173756 51734
rect 173852 51711 173908 51720
rect 173636 48482 173664 51614
rect 173728 51598 173848 51626
rect 173820 51513 173848 51598
rect 174050 51592 174078 52020
rect 174142 51660 174170 52020
rect 174234 51785 174262 52020
rect 174220 51776 174276 51785
rect 174220 51711 174276 51720
rect 174326 51728 174354 52020
rect 174418 51921 174446 52020
rect 174404 51912 174460 51921
rect 174404 51847 174460 51856
rect 174510 51796 174538 52020
rect 174464 51785 174538 51796
rect 174450 51776 174538 51785
rect 174326 51700 174400 51728
rect 174506 51768 174538 51776
rect 174602 51796 174630 52020
rect 174694 51950 174722 52020
rect 174682 51944 174734 51950
rect 174682 51886 174734 51892
rect 174602 51785 174676 51796
rect 174602 51776 174690 51785
rect 174602 51768 174634 51776
rect 174450 51711 174506 51720
rect 174786 51728 174814 52020
rect 174878 51921 174906 52020
rect 174864 51912 174920 51921
rect 174864 51847 174920 51856
rect 174970 51796 174998 52020
rect 174634 51711 174690 51720
rect 174142 51632 174308 51660
rect 174050 51564 174124 51592
rect 173806 51504 173862 51513
rect 174096 51490 174124 51564
rect 174096 51462 174170 51490
rect 173806 51439 173862 51448
rect 174142 51456 174170 51462
rect 174142 51428 174216 51456
rect 174188 51377 174216 51428
rect 174174 51368 174230 51377
rect 173716 51332 173768 51338
rect 174174 51303 174230 51312
rect 173716 51274 173768 51280
rect 173728 50998 173756 51274
rect 173716 50992 173768 50998
rect 173716 50934 173768 50940
rect 174280 50182 174308 51632
rect 174372 50833 174400 51700
rect 174740 51700 174814 51728
rect 174924 51768 174998 51796
rect 174358 50824 174414 50833
rect 174358 50759 174414 50768
rect 174268 50176 174320 50182
rect 174268 50118 174320 50124
rect 173990 50008 174046 50017
rect 173990 49943 174046 49952
rect 174266 50008 174322 50017
rect 174266 49943 174322 49952
rect 173808 49224 173860 49230
rect 173808 49166 173860 49172
rect 173624 48476 173676 48482
rect 173624 48418 173676 48424
rect 173532 46844 173584 46850
rect 173532 46786 173584 46792
rect 173820 41886 173848 49166
rect 174004 48249 174032 49943
rect 173990 48240 174046 48249
rect 173990 48175 174046 48184
rect 174280 48113 174308 49943
rect 174740 48142 174768 51700
rect 174924 51066 174952 51768
rect 175062 51728 175090 52020
rect 175016 51700 175090 51728
rect 175016 51134 175044 51700
rect 175154 51660 175182 52020
rect 175108 51632 175182 51660
rect 175108 51270 175136 51632
rect 175246 51592 175274 52020
rect 175338 51660 175366 52020
rect 175430 51762 175458 52020
rect 175522 51898 175550 52020
rect 175706 51950 175734 52020
rect 175694 51944 175746 51950
rect 175522 51870 175596 51898
rect 175798 51932 175826 52020
rect 175798 51904 175872 51932
rect 175694 51886 175746 51892
rect 175430 51734 175504 51762
rect 175338 51632 175412 51660
rect 175200 51564 175274 51592
rect 175096 51264 175148 51270
rect 175096 51206 175148 51212
rect 175004 51128 175056 51134
rect 175004 51070 175056 51076
rect 174912 51060 174964 51066
rect 174912 51002 174964 51008
rect 175200 48210 175228 51564
rect 175278 51096 175334 51105
rect 175278 51031 175334 51040
rect 175292 50998 175320 51031
rect 175280 50992 175332 50998
rect 175280 50934 175332 50940
rect 175384 49638 175412 51632
rect 175372 49632 175424 49638
rect 175372 49574 175424 49580
rect 175188 48204 175240 48210
rect 175188 48146 175240 48152
rect 174728 48136 174780 48142
rect 174266 48104 174322 48113
rect 174728 48078 174780 48084
rect 174266 48039 174322 48048
rect 175476 47394 175504 51734
rect 175568 50794 175596 51870
rect 175646 51776 175702 51785
rect 175646 51711 175702 51720
rect 175740 51740 175792 51746
rect 175660 51610 175688 51711
rect 175740 51682 175792 51688
rect 175752 51610 175780 51682
rect 175648 51604 175700 51610
rect 175648 51546 175700 51552
rect 175740 51604 175792 51610
rect 175740 51546 175792 51552
rect 175844 51490 175872 51904
rect 175982 51864 176010 52020
rect 176074 51882 176102 52020
rect 176166 51955 176194 52020
rect 176152 51946 176208 51955
rect 175648 51468 175700 51474
rect 175648 51410 175700 51416
rect 175752 51462 175872 51490
rect 175936 51836 176010 51864
rect 176062 51876 176114 51882
rect 176152 51881 176208 51890
rect 175556 50788 175608 50794
rect 175556 50730 175608 50736
rect 175660 50046 175688 51410
rect 175752 51406 175780 51462
rect 175740 51400 175792 51406
rect 175740 51342 175792 51348
rect 175936 50726 175964 51836
rect 176062 51818 176114 51824
rect 176258 51796 176286 52020
rect 176106 51776 176162 51785
rect 176106 51711 176162 51720
rect 176212 51768 176286 51796
rect 176016 51604 176068 51610
rect 176016 51546 176068 51552
rect 175924 50720 175976 50726
rect 175924 50662 175976 50668
rect 176028 50250 176056 51546
rect 176120 51542 176148 51711
rect 176108 51536 176160 51542
rect 176108 51478 176160 51484
rect 176016 50244 176068 50250
rect 176016 50186 176068 50192
rect 175648 50040 175700 50046
rect 175648 49982 175700 49988
rect 176212 49026 176240 51768
rect 176350 51728 176378 52020
rect 176442 51762 176470 52020
rect 176534 51950 176562 52020
rect 176522 51944 176574 51950
rect 176522 51886 176574 51892
rect 176626 51814 176654 52020
rect 176614 51808 176666 51814
rect 176442 51734 176516 51762
rect 176614 51750 176666 51756
rect 176718 51762 176746 52020
rect 176810 51950 176838 52020
rect 176798 51944 176850 51950
rect 176798 51886 176850 51892
rect 176718 51734 176792 51762
rect 176304 51700 176378 51728
rect 176304 50114 176332 51700
rect 176384 51604 176436 51610
rect 176384 51546 176436 51552
rect 176396 51202 176424 51546
rect 176384 51196 176436 51202
rect 176384 51138 176436 51144
rect 176488 50153 176516 51734
rect 176568 51672 176620 51678
rect 176568 51614 176620 51620
rect 176580 50318 176608 51614
rect 176568 50312 176620 50318
rect 176568 50254 176620 50260
rect 176474 50144 176530 50153
rect 176292 50108 176344 50114
rect 176474 50079 176530 50088
rect 176292 50050 176344 50056
rect 176764 49910 176792 51734
rect 176902 51728 176930 52020
rect 177086 51814 177114 52020
rect 177074 51808 177126 51814
rect 177074 51750 177126 51756
rect 177178 51728 177206 52020
rect 177362 51796 177390 52020
rect 177316 51768 177390 51796
rect 176902 51700 176976 51728
rect 177178 51700 177252 51728
rect 176752 49904 176804 49910
rect 176752 49846 176804 49852
rect 176948 49450 176976 51700
rect 177120 51604 177172 51610
rect 177120 51546 177172 51552
rect 177026 49600 177082 49609
rect 177026 49535 177028 49544
rect 177080 49535 177082 49544
rect 177028 49506 177080 49512
rect 176856 49422 176976 49450
rect 176200 49020 176252 49026
rect 176200 48962 176252 48968
rect 176856 48006 176884 49422
rect 176936 49360 176988 49366
rect 176936 49302 176988 49308
rect 176948 48657 176976 49302
rect 177132 49065 177160 51546
rect 177118 49056 177174 49065
rect 177118 48991 177174 49000
rect 177120 48884 177172 48890
rect 177120 48826 177172 48832
rect 176934 48648 176990 48657
rect 176934 48583 176990 48592
rect 176844 48000 176896 48006
rect 176844 47942 176896 47948
rect 176660 47456 176712 47462
rect 176660 47398 176712 47404
rect 175464 47388 175516 47394
rect 175464 47330 175516 47336
rect 175280 46368 175332 46374
rect 175280 46310 175332 46316
rect 174542 46200 174598 46209
rect 174542 46135 174598 46144
rect 173808 41880 173860 41886
rect 173808 41822 173860 41828
rect 173348 41472 173400 41478
rect 173348 41414 173400 41420
rect 173256 3868 173308 3874
rect 173256 3810 173308 3816
rect 174556 3602 174584 46135
rect 174820 43920 174872 43926
rect 174820 43862 174872 43868
rect 174636 43852 174688 43858
rect 174636 43794 174688 43800
rect 174544 3596 174596 3602
rect 174544 3538 174596 3544
rect 174648 3534 174676 43794
rect 174832 43518 174860 43862
rect 174820 43512 174872 43518
rect 174820 43454 174872 43460
rect 175292 16574 175320 46310
rect 175292 16546 175504 16574
rect 173164 3528 173216 3534
rect 173164 3470 173216 3476
rect 174636 3528 174688 3534
rect 174636 3470 174688 3476
rect 173176 480 173204 3470
rect 174268 3460 174320 3466
rect 174268 3402 174320 3408
rect 174280 480 174308 3402
rect 175476 480 175504 16546
rect 176672 11762 176700 47398
rect 177132 45082 177160 48826
rect 177224 46714 177252 51700
rect 177316 49337 177344 51768
rect 177454 51728 177482 52020
rect 177546 51955 177574 52020
rect 177532 51946 177588 51955
rect 177532 51881 177588 51890
rect 177638 51796 177666 52020
rect 177408 51700 177482 51728
rect 177592 51768 177666 51796
rect 177302 49328 177358 49337
rect 177302 49263 177358 49272
rect 177304 48748 177356 48754
rect 177304 48690 177356 48696
rect 177212 46708 177264 46714
rect 177212 46650 177264 46656
rect 177120 45076 177172 45082
rect 177120 45018 177172 45024
rect 176752 43512 176804 43518
rect 176752 43454 176804 43460
rect 176660 11756 176712 11762
rect 176660 11698 176712 11704
rect 176764 6914 176792 43454
rect 176672 6886 176792 6914
rect 176672 480 176700 6886
rect 177316 3398 177344 48690
rect 177408 46646 177436 51700
rect 177592 48521 177620 51768
rect 177730 51728 177758 52020
rect 177684 51700 177758 51728
rect 177684 49201 177712 51700
rect 177822 51660 177850 52020
rect 177914 51728 177942 52020
rect 178006 51921 178034 52020
rect 177992 51912 178048 51921
rect 177992 51847 178048 51856
rect 178098 51796 178126 52020
rect 178052 51768 178126 51796
rect 177914 51700 177988 51728
rect 177776 51632 177850 51660
rect 177776 51513 177804 51632
rect 177762 51504 177818 51513
rect 177762 51439 177818 51448
rect 177960 50522 177988 51700
rect 178052 50590 178080 51768
rect 178190 51728 178218 52020
rect 178144 51700 178218 51728
rect 178040 50584 178092 50590
rect 178040 50526 178092 50532
rect 177948 50516 178000 50522
rect 177948 50458 178000 50464
rect 177764 50448 177816 50454
rect 177764 50390 177816 50396
rect 177776 50153 177804 50390
rect 177762 50144 177818 50153
rect 177762 50079 177818 50088
rect 178144 50046 178172 51700
rect 178282 51660 178310 52020
rect 178374 51950 178402 52020
rect 178362 51944 178414 51950
rect 178362 51886 178414 51892
rect 178466 51728 178494 52020
rect 178236 51632 178310 51660
rect 178420 51700 178494 51728
rect 178558 51728 178586 52020
rect 178650 51921 178678 52020
rect 178636 51912 178692 51921
rect 178636 51847 178692 51856
rect 178742 51762 178770 52020
rect 178834 51882 178862 52020
rect 178926 51921 178954 52020
rect 179018 51950 179046 52020
rect 179110 51950 179138 52020
rect 179006 51944 179058 51950
rect 178912 51912 178968 51921
rect 178822 51876 178874 51882
rect 179006 51886 179058 51892
rect 179098 51944 179150 51950
rect 179098 51886 179150 51892
rect 178912 51847 178968 51856
rect 178822 51818 178874 51824
rect 178696 51734 178770 51762
rect 178958 51776 179014 51785
rect 178558 51700 178632 51728
rect 178132 50040 178184 50046
rect 177762 50008 177818 50017
rect 178132 49982 178184 49988
rect 177762 49943 177818 49952
rect 177670 49192 177726 49201
rect 177670 49127 177726 49136
rect 177672 48544 177724 48550
rect 177578 48512 177634 48521
rect 177672 48486 177724 48492
rect 177578 48447 177634 48456
rect 177488 47184 177540 47190
rect 177488 47126 177540 47132
rect 177396 46640 177448 46646
rect 177396 46582 177448 46588
rect 177500 46288 177528 47126
rect 177580 46980 177632 46986
rect 177580 46922 177632 46928
rect 177408 46260 177528 46288
rect 177408 3942 177436 46260
rect 177488 46164 177540 46170
rect 177488 46106 177540 46112
rect 177396 3936 177448 3942
rect 177396 3878 177448 3884
rect 177500 3738 177528 46106
rect 177592 20670 177620 46922
rect 177684 24857 177712 48486
rect 177776 47530 177804 49943
rect 177854 49328 177910 49337
rect 177854 49263 177910 49272
rect 177948 49292 178000 49298
rect 177868 49094 177896 49263
rect 177948 49234 178000 49240
rect 177960 49201 177988 49234
rect 177946 49192 178002 49201
rect 177946 49127 178002 49136
rect 177856 49088 177908 49094
rect 177856 49030 177908 49036
rect 177948 48952 178000 48958
rect 177946 48920 177948 48929
rect 178000 48920 178002 48929
rect 177946 48855 178002 48864
rect 178236 48074 178264 51632
rect 178420 50810 178448 51700
rect 178500 51604 178552 51610
rect 178500 51546 178552 51552
rect 178328 50782 178448 50810
rect 178328 48385 178356 50782
rect 178408 50584 178460 50590
rect 178408 50526 178460 50532
rect 178314 48376 178370 48385
rect 178314 48311 178370 48320
rect 178420 48278 178448 50526
rect 178512 49434 178540 51546
rect 178500 49428 178552 49434
rect 178500 49370 178552 49376
rect 178408 48272 178460 48278
rect 178408 48214 178460 48220
rect 178224 48068 178276 48074
rect 178224 48010 178276 48016
rect 177764 47524 177816 47530
rect 177764 47466 177816 47472
rect 177764 47252 177816 47258
rect 177764 47194 177816 47200
rect 177776 46170 177804 47194
rect 178604 46782 178632 51700
rect 178696 48686 178724 51734
rect 179202 51762 179230 52020
rect 179294 51882 179322 52020
rect 179386 51950 179414 52020
rect 179374 51944 179426 51950
rect 179374 51886 179426 51892
rect 179478 51882 179506 52020
rect 179570 51882 179598 52020
rect 179662 51921 179690 52020
rect 179648 51912 179704 51921
rect 179282 51876 179334 51882
rect 179282 51818 179334 51824
rect 179466 51876 179518 51882
rect 179466 51818 179518 51824
rect 179558 51876 179610 51882
rect 179648 51847 179704 51856
rect 179558 51818 179610 51824
rect 179754 51796 179782 52020
rect 179708 51768 179782 51796
rect 178958 51711 179014 51720
rect 179052 51740 179104 51746
rect 178866 51504 178922 51513
rect 178972 51474 179000 51711
rect 179202 51734 179322 51762
rect 179052 51682 179104 51688
rect 178866 51439 178922 51448
rect 178960 51468 179012 51474
rect 178776 51196 178828 51202
rect 178776 51138 178828 51144
rect 178788 51105 178816 51138
rect 178774 51096 178830 51105
rect 178774 51031 178830 51040
rect 178880 50182 178908 51439
rect 178960 51410 179012 51416
rect 178960 51332 179012 51338
rect 178960 51274 179012 51280
rect 178868 50176 178920 50182
rect 178868 50118 178920 50124
rect 178684 48680 178736 48686
rect 178684 48622 178736 48628
rect 178868 47320 178920 47326
rect 178868 47262 178920 47268
rect 178684 47116 178736 47122
rect 178684 47058 178736 47064
rect 178592 46776 178644 46782
rect 178592 46718 178644 46724
rect 177764 46164 177816 46170
rect 177764 46106 177816 46112
rect 178040 44940 178092 44946
rect 178040 44882 178092 44888
rect 177670 24848 177726 24857
rect 177670 24783 177726 24792
rect 177580 20664 177632 20670
rect 177580 20606 177632 20612
rect 178052 16574 178080 44882
rect 178052 16546 178632 16574
rect 177856 11756 177908 11762
rect 177856 11698 177908 11704
rect 177488 3732 177540 3738
rect 177488 3674 177540 3680
rect 177304 3392 177356 3398
rect 177304 3334 177356 3340
rect 177868 480 177896 11698
rect 170742 354 170854 480
rect 170324 326 170854 354
rect 170742 -960 170854 326
rect 171938 -960 172050 480
rect 173134 -960 173246 480
rect 174238 -960 174350 480
rect 175434 -960 175546 480
rect 176630 -960 176742 480
rect 177826 -960 177938 480
rect 178604 354 178632 16546
rect 178696 3330 178724 47058
rect 178776 47048 178828 47054
rect 178776 46990 178828 46996
rect 178788 3670 178816 46990
rect 178776 3664 178828 3670
rect 178776 3606 178828 3612
rect 178880 3466 178908 47262
rect 178972 12034 179000 51274
rect 179064 50658 179092 51682
rect 179294 51660 179322 51734
rect 179604 51740 179656 51746
rect 179604 51682 179656 51688
rect 179420 51672 179472 51678
rect 179294 51632 179368 51660
rect 179142 51232 179198 51241
rect 179142 51167 179144 51176
rect 179196 51167 179198 51176
rect 179144 51138 179196 51144
rect 179236 50788 179288 50794
rect 179236 50730 179288 50736
rect 179052 50652 179104 50658
rect 179052 50594 179104 50600
rect 179248 50386 179276 50730
rect 179236 50380 179288 50386
rect 179236 50322 179288 50328
rect 179340 48822 179368 51632
rect 179420 51614 179472 51620
rect 179432 48958 179460 51614
rect 179512 51604 179564 51610
rect 179512 51546 179564 51552
rect 179524 50590 179552 51546
rect 179512 50584 179564 50590
rect 179512 50526 179564 50532
rect 179512 50448 179564 50454
rect 179512 50390 179564 50396
rect 179420 48952 179472 48958
rect 179420 48894 179472 48900
rect 179328 48816 179380 48822
rect 179328 48758 179380 48764
rect 179052 48680 179104 48686
rect 179052 48622 179104 48628
rect 178960 12028 179012 12034
rect 178960 11970 179012 11976
rect 179064 11830 179092 48622
rect 179144 48408 179196 48414
rect 179144 48350 179196 48356
rect 179156 25498 179184 48350
rect 179524 48346 179552 50390
rect 179616 49162 179644 51682
rect 179604 49156 179656 49162
rect 179604 49098 179656 49104
rect 179604 49020 179656 49026
rect 179604 48962 179656 48968
rect 179236 48340 179288 48346
rect 179236 48282 179288 48288
rect 179512 48340 179564 48346
rect 179512 48282 179564 48288
rect 179248 25566 179276 48282
rect 179616 48090 179644 48962
rect 179432 48062 179644 48090
rect 179708 48090 179736 51768
rect 179846 51728 179874 52020
rect 179800 51700 179874 51728
rect 179800 50810 179828 51700
rect 179938 51592 179966 52020
rect 180030 51882 180058 52020
rect 180122 51950 180150 52020
rect 180214 51950 180242 52020
rect 180110 51944 180162 51950
rect 180110 51886 180162 51892
rect 180202 51944 180254 51950
rect 180202 51886 180254 51892
rect 180018 51876 180070 51882
rect 180018 51818 180070 51824
rect 180306 51728 180334 52020
rect 180398 51921 180426 52020
rect 180490 51950 180518 52020
rect 180478 51944 180530 51950
rect 180384 51912 180440 51921
rect 180478 51886 180530 51892
rect 180582 51882 180610 52020
rect 180384 51847 180440 51856
rect 180570 51876 180622 51882
rect 180570 51818 180622 51824
rect 180674 51814 180702 52020
rect 180432 51808 180484 51814
rect 180432 51750 180484 51756
rect 180662 51808 180714 51814
rect 180662 51750 180714 51756
rect 180260 51700 180334 51728
rect 179938 51564 180012 51592
rect 179800 50782 179920 50810
rect 179788 50652 179840 50658
rect 179788 50594 179840 50600
rect 179800 49094 179828 50594
rect 179892 50454 179920 50782
rect 179880 50448 179932 50454
rect 179880 50390 179932 50396
rect 179880 49156 179932 49162
rect 179880 49098 179932 49104
rect 179788 49088 179840 49094
rect 179788 49030 179840 49036
rect 179788 48952 179840 48958
rect 179788 48894 179840 48900
rect 179800 48550 179828 48894
rect 179788 48544 179840 48550
rect 179788 48486 179840 48492
rect 179708 48062 179828 48090
rect 179432 29646 179460 48062
rect 179604 48000 179656 48006
rect 179604 47942 179656 47948
rect 179420 29640 179472 29646
rect 179420 29582 179472 29588
rect 179236 25560 179288 25566
rect 179236 25502 179288 25508
rect 179144 25492 179196 25498
rect 179144 25434 179196 25440
rect 179420 22772 179472 22778
rect 179420 22714 179472 22720
rect 179432 16574 179460 22714
rect 179616 17474 179644 47942
rect 179696 47932 179748 47938
rect 179696 47874 179748 47880
rect 179708 25634 179736 47874
rect 179800 25702 179828 48062
rect 179892 25770 179920 49098
rect 179984 48414 180012 51564
rect 180260 51490 180288 51700
rect 180214 51462 180288 51490
rect 180340 51536 180392 51542
rect 180340 51478 180392 51484
rect 180214 51456 180242 51462
rect 180168 51428 180242 51456
rect 180064 51400 180116 51406
rect 180064 51342 180116 51348
rect 179972 48408 180024 48414
rect 179972 48350 180024 48356
rect 179970 47968 180026 47977
rect 180076 47938 180104 51342
rect 180168 47977 180196 51428
rect 180248 51128 180300 51134
rect 180248 51070 180300 51076
rect 180154 47968 180210 47977
rect 179970 47903 180026 47912
rect 180064 47932 180116 47938
rect 179880 25764 179932 25770
rect 179880 25706 179932 25712
rect 179788 25696 179840 25702
rect 179788 25638 179840 25644
rect 179696 25628 179748 25634
rect 179696 25570 179748 25576
rect 179984 25430 180012 47903
rect 180154 47903 180210 47912
rect 180064 47874 180116 47880
rect 180260 46238 180288 51070
rect 180352 46986 180380 51478
rect 180444 47977 180472 51750
rect 180524 51740 180576 51746
rect 180524 51682 180576 51688
rect 180536 50658 180564 51682
rect 180616 51672 180668 51678
rect 180766 51660 180794 52020
rect 180858 51814 180886 52020
rect 180846 51808 180898 51814
rect 180846 51750 180898 51756
rect 180950 51660 180978 52020
rect 181042 51955 181070 52020
rect 181028 51946 181084 51955
rect 181134 51950 181162 52020
rect 181226 51950 181254 52020
rect 181318 51955 181346 52020
rect 181028 51881 181084 51890
rect 181122 51944 181174 51950
rect 181122 51886 181174 51892
rect 181214 51944 181266 51950
rect 181214 51886 181266 51892
rect 181304 51946 181360 51955
rect 181304 51881 181360 51890
rect 181260 51808 181312 51814
rect 180616 51614 180668 51620
rect 180720 51632 180794 51660
rect 180904 51632 180978 51660
rect 181088 51768 181260 51796
rect 180524 50652 180576 50658
rect 180524 50594 180576 50600
rect 180524 48408 180576 48414
rect 180524 48350 180576 48356
rect 180430 47968 180486 47977
rect 180430 47903 180486 47912
rect 180340 46980 180392 46986
rect 180340 46922 180392 46928
rect 180248 46232 180300 46238
rect 180248 46174 180300 46180
rect 180536 44198 180564 48350
rect 180628 48006 180656 51614
rect 180616 48000 180668 48006
rect 180616 47942 180668 47948
rect 180524 44192 180576 44198
rect 180524 44134 180576 44140
rect 180720 41414 180748 51632
rect 180800 51468 180852 51474
rect 180800 51410 180852 51416
rect 180812 51134 180840 51410
rect 180904 51338 180932 51632
rect 181088 51490 181116 51768
rect 181260 51750 181312 51756
rect 181168 51672 181220 51678
rect 181220 51632 181300 51660
rect 181168 51614 181220 51620
rect 180996 51462 181116 51490
rect 181168 51536 181220 51542
rect 181168 51478 181220 51484
rect 180892 51332 180944 51338
rect 180892 51274 180944 51280
rect 180800 51128 180852 51134
rect 180800 51070 180852 51076
rect 180890 48512 180946 48521
rect 180890 48447 180946 48456
rect 180800 48068 180852 48074
rect 180800 48010 180852 48016
rect 180260 41386 180748 41414
rect 179972 25424 180024 25430
rect 179972 25366 180024 25372
rect 180260 17542 180288 41386
rect 180248 17536 180300 17542
rect 180248 17478 180300 17484
rect 179604 17468 179656 17474
rect 179604 17410 179656 17416
rect 180812 16574 180840 48010
rect 180904 47190 180932 48447
rect 180892 47184 180944 47190
rect 180892 47126 180944 47132
rect 180996 44174 181024 51462
rect 181076 51400 181128 51406
rect 181076 51342 181128 51348
rect 181088 44849 181116 51342
rect 181180 47977 181208 51478
rect 181272 48385 181300 51632
rect 181410 51626 181438 52020
rect 181502 51728 181530 52020
rect 181594 51882 181622 52020
rect 181582 51876 181634 51882
rect 181582 51818 181634 51824
rect 181686 51762 181714 52020
rect 181640 51746 181714 51762
rect 181628 51740 181714 51746
rect 181502 51700 181576 51728
rect 181364 51598 181438 51626
rect 181258 48376 181314 48385
rect 181258 48311 181314 48320
rect 181166 47968 181222 47977
rect 181166 47903 181222 47912
rect 181260 47184 181312 47190
rect 181260 47126 181312 47132
rect 181074 44840 181130 44849
rect 181074 44775 181130 44784
rect 180904 44146 181024 44174
rect 180904 43450 180932 44146
rect 180892 43444 180944 43450
rect 180892 43386 180944 43392
rect 181272 41414 181300 47126
rect 181364 44174 181392 51598
rect 181444 51536 181496 51542
rect 181444 51478 181496 51484
rect 181456 47190 181484 51478
rect 181548 47258 181576 51700
rect 181680 51734 181714 51740
rect 181628 51682 181680 51688
rect 181778 51660 181806 52020
rect 181870 51814 181898 52020
rect 181858 51808 181910 51814
rect 181858 51750 181910 51756
rect 181732 51632 181806 51660
rect 181732 51626 181760 51632
rect 181640 51598 181760 51626
rect 181536 47252 181588 47258
rect 181536 47194 181588 47200
rect 181444 47184 181496 47190
rect 181444 47126 181496 47132
rect 181640 44878 181668 51598
rect 181720 51536 181772 51542
rect 181962 51524 181990 52020
rect 182054 51762 182082 52020
rect 182146 51882 182174 52020
rect 182238 51950 182266 52020
rect 182330 51950 182358 52020
rect 182422 51955 182450 52020
rect 182226 51944 182278 51950
rect 182226 51886 182278 51892
rect 182318 51944 182370 51950
rect 182318 51886 182370 51892
rect 182408 51946 182464 51955
rect 182514 51950 182542 52020
rect 182606 51950 182634 52020
rect 182698 51950 182726 52020
rect 182882 51950 182910 52020
rect 182974 51955 183002 52020
rect 182134 51876 182186 51882
rect 182408 51881 182464 51890
rect 182502 51944 182554 51950
rect 182502 51886 182554 51892
rect 182594 51944 182646 51950
rect 182594 51886 182646 51892
rect 182686 51944 182738 51950
rect 182686 51886 182738 51892
rect 182870 51944 182922 51950
rect 182870 51886 182922 51892
rect 182960 51946 183016 51955
rect 182960 51881 183016 51890
rect 182134 51818 182186 51824
rect 182364 51808 182416 51814
rect 182054 51734 182128 51762
rect 182364 51750 182416 51756
rect 182100 51626 182128 51734
rect 182272 51672 182324 51678
rect 182100 51598 182220 51626
rect 182272 51614 182324 51620
rect 181720 51478 181772 51484
rect 181916 51496 181990 51524
rect 182088 51536 182140 51542
rect 181628 44872 181680 44878
rect 181628 44814 181680 44820
rect 181364 44146 181576 44174
rect 181272 41386 181392 41414
rect 181364 37942 181392 41386
rect 181352 37936 181404 37942
rect 181352 37878 181404 37884
rect 181548 26926 181576 44146
rect 181732 35222 181760 51478
rect 181812 49836 181864 49842
rect 181812 49778 181864 49784
rect 181824 47462 181852 49778
rect 181812 47456 181864 47462
rect 181812 47398 181864 47404
rect 181916 47054 181944 51496
rect 182088 51478 182140 51484
rect 181996 49904 182048 49910
rect 181996 49846 182048 49852
rect 181904 47048 181956 47054
rect 181904 46990 181956 46996
rect 182008 45014 182036 49846
rect 182100 46306 182128 51478
rect 182192 49910 182220 51598
rect 182180 49904 182232 49910
rect 182180 49846 182232 49852
rect 182180 49768 182232 49774
rect 182180 49710 182232 49716
rect 182192 47569 182220 49710
rect 182284 48793 182312 51614
rect 182376 49065 182404 51750
rect 182548 51740 182600 51746
rect 182548 51682 182600 51688
rect 182454 49736 182510 49745
rect 182454 49671 182510 49680
rect 182362 49056 182418 49065
rect 182362 48991 182418 49000
rect 182364 48952 182416 48958
rect 182364 48894 182416 48900
rect 182270 48784 182326 48793
rect 182270 48719 182326 48728
rect 182178 47560 182234 47569
rect 182178 47495 182234 47504
rect 182376 46374 182404 48894
rect 182364 46368 182416 46374
rect 182364 46310 182416 46316
rect 182088 46300 182140 46306
rect 182088 46242 182140 46248
rect 181996 45008 182048 45014
rect 181996 44950 182048 44956
rect 182468 36718 182496 49671
rect 182560 48521 182588 51682
rect 182732 51672 182784 51678
rect 182732 51614 182784 51620
rect 183066 51626 183094 52020
rect 183158 51950 183186 52020
rect 183250 51950 183278 52020
rect 183342 51950 183370 52020
rect 183146 51944 183198 51950
rect 183146 51886 183198 51892
rect 183238 51944 183290 51950
rect 183238 51886 183290 51892
rect 183330 51944 183382 51950
rect 183330 51886 183382 51892
rect 183284 51808 183336 51814
rect 183284 51750 183336 51756
rect 183192 51740 183244 51746
rect 183192 51682 183244 51688
rect 182640 51604 182692 51610
rect 182640 51546 182692 51552
rect 182546 48512 182602 48521
rect 182546 48447 182602 48456
rect 182652 47598 182680 51546
rect 182744 51490 182772 51614
rect 182916 51604 182968 51610
rect 183066 51598 183140 51626
rect 182916 51546 182968 51552
rect 182744 51462 182864 51490
rect 182732 51400 182784 51406
rect 182732 51342 182784 51348
rect 182640 47592 182692 47598
rect 182640 47534 182692 47540
rect 182456 36712 182508 36718
rect 182456 36654 182508 36660
rect 181720 35216 181772 35222
rect 181720 35158 181772 35164
rect 181536 26920 181588 26926
rect 181536 26862 181588 26868
rect 179432 16546 180288 16574
rect 180812 16546 181024 16574
rect 179052 11824 179104 11830
rect 179052 11766 179104 11772
rect 178868 3460 178920 3466
rect 178868 3402 178920 3408
rect 178684 3324 178736 3330
rect 178684 3266 178736 3272
rect 180260 480 180288 16546
rect 179022 354 179134 480
rect 178604 326 179134 354
rect 179022 -960 179134 326
rect 180218 -960 180330 480
rect 180996 354 181024 16546
rect 182364 11484 182416 11490
rect 182364 11426 182416 11432
rect 181414 354 181526 480
rect 180996 326 181526 354
rect 182376 354 182404 11426
rect 182744 4826 182772 51342
rect 182836 43926 182864 51462
rect 182928 46442 182956 51546
rect 183008 51536 183060 51542
rect 183008 51478 183060 51484
rect 182916 46436 182968 46442
rect 182916 46378 182968 46384
rect 182916 46300 182968 46306
rect 182916 46242 182968 46248
rect 182824 43920 182876 43926
rect 182824 43862 182876 43868
rect 182928 6390 182956 46242
rect 183020 26994 183048 51478
rect 183112 45082 183140 51598
rect 183100 45076 183152 45082
rect 183100 45018 183152 45024
rect 183204 43790 183232 51682
rect 183296 47122 183324 51750
rect 183434 51626 183462 52020
rect 183526 51796 183554 52020
rect 183618 51921 183646 52020
rect 183710 51950 183738 52020
rect 183698 51944 183750 51950
rect 183604 51912 183660 51921
rect 183698 51886 183750 51892
rect 183604 51847 183660 51856
rect 183652 51808 183704 51814
rect 183526 51768 183600 51796
rect 183388 51598 183462 51626
rect 183388 48754 183416 51598
rect 183572 51490 183600 51768
rect 183652 51750 183704 51756
rect 183480 51462 183600 51490
rect 183376 48748 183428 48754
rect 183376 48690 183428 48696
rect 183284 47116 183336 47122
rect 183284 47058 183336 47064
rect 183480 46306 183508 51462
rect 183664 49688 183692 51750
rect 183802 51728 183830 52020
rect 183894 51950 183922 52020
rect 183986 51950 184014 52020
rect 184078 51950 184106 52020
rect 183882 51944 183934 51950
rect 183882 51886 183934 51892
rect 183974 51944 184026 51950
rect 183974 51886 184026 51892
rect 184066 51944 184118 51950
rect 184170 51921 184198 52020
rect 184262 51950 184290 52020
rect 184250 51944 184302 51950
rect 184066 51886 184118 51892
rect 184156 51912 184212 51921
rect 184446 51898 184474 52020
rect 184250 51886 184302 51892
rect 184400 51882 184474 51898
rect 184156 51847 184212 51856
rect 184388 51876 184474 51882
rect 184440 51870 184474 51876
rect 184388 51818 184440 51824
rect 184204 51808 184256 51814
rect 184204 51750 184256 51756
rect 183572 49660 183692 49688
rect 183756 51700 183830 51728
rect 184020 51740 184072 51746
rect 183572 47104 183600 49660
rect 183756 48686 183784 51700
rect 184020 51682 184072 51688
rect 184112 51740 184164 51746
rect 184112 51682 184164 51688
rect 183928 51672 183980 51678
rect 183928 51614 183980 51620
rect 183836 50448 183888 50454
rect 183836 50390 183888 50396
rect 183744 48680 183796 48686
rect 183744 48622 183796 48628
rect 183848 48074 183876 50390
rect 183940 49745 183968 51614
rect 184032 49774 184060 51682
rect 184020 49768 184072 49774
rect 183926 49736 183982 49745
rect 184020 49710 184072 49716
rect 183926 49671 183982 49680
rect 184124 49450 184152 51682
rect 183940 49422 184152 49450
rect 183940 48890 183968 49422
rect 184216 49008 184244 51750
rect 184388 51740 184440 51746
rect 184538 51728 184566 52020
rect 184630 51921 184658 52020
rect 184616 51912 184672 51921
rect 184616 51847 184672 51856
rect 184722 51796 184750 52020
rect 184676 51768 184750 51796
rect 184538 51700 184612 51728
rect 184388 51682 184440 51688
rect 184296 51672 184348 51678
rect 184296 51614 184348 51620
rect 184032 48980 184244 49008
rect 183928 48884 183980 48890
rect 183928 48826 183980 48832
rect 184032 48414 184060 48980
rect 184308 48770 184336 51614
rect 184124 48742 184336 48770
rect 184020 48408 184072 48414
rect 184020 48350 184072 48356
rect 183836 48068 183888 48074
rect 183836 48010 183888 48016
rect 183572 47076 183692 47104
rect 183560 46980 183612 46986
rect 183560 46922 183612 46928
rect 183468 46300 183520 46306
rect 183468 46242 183520 46248
rect 183192 43784 183244 43790
rect 183192 43726 183244 43732
rect 183008 26988 183060 26994
rect 183008 26930 183060 26936
rect 183572 16574 183600 46922
rect 183664 46209 183692 47076
rect 183650 46200 183706 46209
rect 183650 46135 183706 46144
rect 184124 43722 184152 48742
rect 184204 48544 184256 48550
rect 184204 48486 184256 48492
rect 184112 43716 184164 43722
rect 184112 43658 184164 43664
rect 183572 16546 183784 16574
rect 182916 6384 182968 6390
rect 182916 6326 182968 6332
rect 182732 4820 182784 4826
rect 182732 4762 182784 4768
rect 183756 480 183784 16546
rect 184216 11490 184244 48486
rect 184400 47326 184428 51682
rect 184584 48958 184612 51700
rect 184676 49842 184704 51768
rect 184814 51626 184842 52020
rect 184906 51950 184934 52020
rect 184894 51944 184946 51950
rect 184894 51886 184946 51892
rect 184998 51762 185026 52020
rect 185090 51814 185118 52020
rect 185182 51950 185210 52020
rect 185274 51950 185302 52020
rect 185366 51950 185394 52020
rect 185458 51950 185486 52020
rect 185170 51944 185222 51950
rect 185170 51886 185222 51892
rect 185262 51944 185314 51950
rect 185262 51886 185314 51892
rect 185354 51944 185406 51950
rect 185354 51886 185406 51892
rect 185446 51944 185498 51950
rect 185446 51886 185498 51892
rect 184768 51598 184842 51626
rect 184952 51734 185026 51762
rect 185078 51808 185130 51814
rect 185078 51750 185130 51756
rect 185550 51762 185578 52020
rect 185642 51921 185670 52020
rect 185628 51912 185684 51921
rect 185628 51847 185684 51856
rect 185216 51740 185268 51746
rect 184664 49836 184716 49842
rect 184664 49778 184716 49784
rect 184572 48952 184624 48958
rect 184572 48894 184624 48900
rect 184478 48784 184534 48793
rect 184768 48770 184796 51598
rect 184848 51536 184900 51542
rect 184848 51478 184900 51484
rect 184478 48719 184534 48728
rect 184676 48742 184796 48770
rect 184388 47320 184440 47326
rect 184388 47262 184440 47268
rect 184388 47184 184440 47190
rect 184388 47126 184440 47132
rect 184400 22778 184428 47126
rect 184492 33794 184520 48719
rect 184570 48512 184626 48521
rect 184570 48447 184626 48456
rect 184584 43518 184612 48447
rect 184676 44946 184704 48742
rect 184754 48376 184810 48385
rect 184754 48311 184810 48320
rect 184664 44940 184716 44946
rect 184664 44882 184716 44888
rect 184572 43512 184624 43518
rect 184572 43454 184624 43460
rect 184768 41414 184796 48311
rect 184860 47190 184888 51478
rect 184952 50454 184980 51734
rect 185216 51682 185268 51688
rect 185308 51740 185360 51746
rect 185308 51682 185360 51688
rect 185400 51740 185452 51746
rect 185550 51734 185624 51762
rect 185400 51682 185452 51688
rect 185032 51672 185084 51678
rect 185032 51614 185084 51620
rect 185124 51672 185176 51678
rect 185124 51614 185176 51620
rect 184940 50448 184992 50454
rect 184940 50390 184992 50396
rect 184940 50176 184992 50182
rect 184940 50118 184992 50124
rect 184848 47184 184900 47190
rect 184848 47126 184900 47132
rect 184952 46986 184980 50118
rect 185044 48550 185072 51614
rect 185032 48544 185084 48550
rect 185032 48486 185084 48492
rect 184940 46980 184992 46986
rect 184940 46922 184992 46928
rect 184768 41386 184888 41414
rect 184480 33788 184532 33794
rect 184480 33730 184532 33736
rect 184388 22772 184440 22778
rect 184388 22714 184440 22720
rect 184204 11484 184256 11490
rect 184204 11426 184256 11432
rect 184860 3330 184888 41386
rect 185136 5574 185164 51614
rect 185228 46510 185256 51682
rect 185216 46504 185268 46510
rect 185216 46446 185268 46452
rect 185216 46368 185268 46374
rect 185216 46310 185268 46316
rect 185228 12442 185256 46310
rect 185320 46238 185348 51682
rect 185308 46232 185360 46238
rect 185308 46174 185360 46180
rect 185308 46096 185360 46102
rect 185308 46038 185360 46044
rect 185320 22778 185348 46038
rect 185412 25702 185440 51682
rect 185596 51678 185624 51734
rect 185584 51672 185636 51678
rect 185584 51614 185636 51620
rect 185734 51592 185762 52020
rect 185826 51882 185854 52020
rect 185918 51950 185946 52020
rect 185906 51944 185958 51950
rect 185906 51886 185958 51892
rect 185814 51876 185866 51882
rect 185814 51818 185866 51824
rect 186010 51660 186038 52020
rect 186102 51882 186130 52020
rect 186090 51876 186142 51882
rect 186090 51818 186142 51824
rect 186194 51762 186222 52020
rect 186286 51950 186314 52020
rect 186274 51944 186326 51950
rect 186274 51886 186326 51892
rect 186378 51882 186406 52020
rect 186366 51876 186418 51882
rect 186366 51818 186418 51824
rect 186470 51762 186498 52020
rect 186562 51950 186590 52020
rect 186550 51944 186602 51950
rect 186550 51886 186602 51892
rect 186654 51762 186682 52020
rect 185688 51564 185762 51592
rect 185964 51632 186038 51660
rect 186148 51734 186222 51762
rect 186424 51734 186498 51762
rect 186608 51734 186682 51762
rect 185584 51536 185636 51542
rect 185584 51478 185636 51484
rect 185596 50182 185624 51478
rect 185584 50176 185636 50182
rect 185584 50118 185636 50124
rect 185688 48314 185716 51564
rect 185768 51468 185820 51474
rect 185768 51410 185820 51416
rect 185596 48286 185716 48314
rect 185596 45286 185624 48286
rect 185780 46374 185808 51410
rect 185860 51400 185912 51406
rect 185860 51342 185912 51348
rect 185872 46986 185900 51342
rect 185860 46980 185912 46986
rect 185860 46922 185912 46928
rect 185860 46504 185912 46510
rect 185860 46446 185912 46452
rect 185768 46368 185820 46374
rect 185768 46310 185820 46316
rect 185768 46232 185820 46238
rect 185768 46174 185820 46180
rect 185584 45280 185636 45286
rect 185584 45222 185636 45228
rect 185400 25696 185452 25702
rect 185400 25638 185452 25644
rect 185308 22772 185360 22778
rect 185308 22714 185360 22720
rect 185216 12436 185268 12442
rect 185216 12378 185268 12384
rect 185124 5568 185176 5574
rect 185124 5510 185176 5516
rect 184940 3596 184992 3602
rect 184940 3538 184992 3544
rect 184848 3324 184900 3330
rect 184848 3266 184900 3272
rect 184952 480 184980 3538
rect 185780 3482 185808 46174
rect 185872 3602 185900 46446
rect 185964 46102 185992 51632
rect 186044 51536 186096 51542
rect 186044 51478 186096 51484
rect 186056 48521 186084 51478
rect 186042 48512 186098 48521
rect 186042 48447 186098 48456
rect 186148 48385 186176 51734
rect 186228 51672 186280 51678
rect 186228 51614 186280 51620
rect 186240 48890 186268 51614
rect 186320 51604 186372 51610
rect 186320 51546 186372 51552
rect 186228 48884 186280 48890
rect 186228 48826 186280 48832
rect 186134 48376 186190 48385
rect 186134 48311 186190 48320
rect 186044 46980 186096 46986
rect 186044 46922 186096 46928
rect 185952 46096 186004 46102
rect 185952 46038 186004 46044
rect 186056 42838 186084 46922
rect 186044 42832 186096 42838
rect 186044 42774 186096 42780
rect 186332 3874 186360 51546
rect 186424 3942 186452 51734
rect 186504 51672 186556 51678
rect 186504 51614 186556 51620
rect 186516 50232 186544 51614
rect 186608 51542 186636 51734
rect 186746 51660 186774 52020
rect 186838 51882 186866 52020
rect 186826 51876 186878 51882
rect 186826 51818 186878 51824
rect 186930 51762 186958 52020
rect 187022 51921 187050 52020
rect 187008 51912 187064 51921
rect 187008 51847 187064 51856
rect 187114 51762 187142 52020
rect 186700 51632 186774 51660
rect 186884 51734 186958 51762
rect 187068 51734 187142 51762
rect 187206 51762 187234 52020
rect 187298 51882 187326 52020
rect 187390 51882 187418 52020
rect 187482 51950 187510 52020
rect 187470 51944 187522 51950
rect 187470 51886 187522 51892
rect 187286 51876 187338 51882
rect 187286 51818 187338 51824
rect 187378 51876 187430 51882
rect 187378 51818 187430 51824
rect 187574 51762 187602 52020
rect 187206 51734 187280 51762
rect 186596 51536 186648 51542
rect 186596 51478 186648 51484
rect 186516 50204 186636 50232
rect 186502 50144 186558 50153
rect 186502 50079 186558 50088
rect 186412 3936 186464 3942
rect 186412 3878 186464 3884
rect 186320 3868 186372 3874
rect 186320 3810 186372 3816
rect 186516 3806 186544 50079
rect 186608 46306 186636 50204
rect 186700 48686 186728 51632
rect 186780 51536 186832 51542
rect 186780 51478 186832 51484
rect 186792 49434 186820 51478
rect 186780 49428 186832 49434
rect 186780 49370 186832 49376
rect 186780 49292 186832 49298
rect 186780 49234 186832 49240
rect 186688 48680 186740 48686
rect 186688 48622 186740 48628
rect 186792 46442 186820 49234
rect 186780 46436 186832 46442
rect 186780 46378 186832 46384
rect 186596 46300 186648 46306
rect 186596 46242 186648 46248
rect 186884 46186 186912 51734
rect 186964 51672 187016 51678
rect 186964 51614 187016 51620
rect 186976 49298 187004 51614
rect 186964 49292 187016 49298
rect 186964 49234 187016 49240
rect 186964 49156 187016 49162
rect 186964 49098 187016 49104
rect 186976 46986 187004 49098
rect 186964 46980 187016 46986
rect 186964 46922 187016 46928
rect 186608 46158 186912 46186
rect 186608 10334 186636 46158
rect 187068 41414 187096 51734
rect 187148 51672 187200 51678
rect 187148 51614 187200 51620
rect 187160 49162 187188 51614
rect 187148 49156 187200 49162
rect 187148 49098 187200 49104
rect 187146 49056 187202 49065
rect 187146 48991 187202 49000
rect 187160 48385 187188 48991
rect 187252 48521 187280 51734
rect 187344 51734 187602 51762
rect 187344 49026 187372 51734
rect 187424 51672 187476 51678
rect 187424 51614 187476 51620
rect 187516 51672 187568 51678
rect 187666 51660 187694 52020
rect 187758 51762 187786 52020
rect 187850 51950 187878 52020
rect 187838 51944 187890 51950
rect 187838 51886 187890 51892
rect 187758 51734 187832 51762
rect 187516 51614 187568 51620
rect 187620 51632 187694 51660
rect 187332 49020 187384 49026
rect 187332 48962 187384 48968
rect 187332 48884 187384 48890
rect 187332 48826 187384 48832
rect 187238 48512 187294 48521
rect 187238 48447 187294 48456
rect 187146 48376 187202 48385
rect 187146 48311 187202 48320
rect 187344 41414 187372 48826
rect 187436 48385 187464 51614
rect 187528 48657 187556 51614
rect 187620 48793 187648 51632
rect 187700 51536 187752 51542
rect 187700 51478 187752 51484
rect 187712 49706 187740 51478
rect 187700 49700 187752 49706
rect 187700 49642 187752 49648
rect 187700 49428 187752 49434
rect 187700 49370 187752 49376
rect 187606 48784 187662 48793
rect 187606 48719 187662 48728
rect 187712 48668 187740 49370
rect 187514 48648 187570 48657
rect 187514 48583 187570 48592
rect 187620 48640 187740 48668
rect 187422 48376 187478 48385
rect 187422 48311 187478 48320
rect 187620 44130 187648 48640
rect 187608 44124 187660 44130
rect 187608 44066 187660 44072
rect 186700 41386 187096 41414
rect 187160 41386 187372 41414
rect 186700 19990 186728 41386
rect 186780 25696 186832 25702
rect 186780 25638 186832 25644
rect 186688 19984 186740 19990
rect 186688 19926 186740 19932
rect 186792 16574 186820 25638
rect 186792 16546 186912 16574
rect 186596 10328 186648 10334
rect 186596 10270 186648 10276
rect 186504 3800 186556 3806
rect 186504 3742 186556 3748
rect 185860 3596 185912 3602
rect 185860 3538 185912 3544
rect 185780 3454 186176 3482
rect 186148 480 186176 3454
rect 182518 354 182630 480
rect 182376 326 182630 354
rect 181414 -960 181526 326
rect 182518 -960 182630 326
rect 183714 -960 183826 480
rect 184910 -960 185022 480
rect 186106 -960 186218 480
rect 186884 354 186912 16546
rect 187160 10402 187188 41386
rect 187148 10396 187200 10402
rect 187148 10338 187200 10344
rect 187804 6866 187832 51734
rect 187942 51660 187970 52020
rect 188034 51932 188062 52020
rect 188034 51904 188154 51932
rect 188126 51762 188154 51904
rect 188218 51882 188246 52020
rect 188310 51882 188338 52020
rect 188206 51876 188258 51882
rect 188206 51818 188258 51824
rect 188298 51876 188350 51882
rect 188298 51818 188350 51824
rect 188402 51762 188430 52020
rect 188494 51882 188522 52020
rect 188482 51876 188534 51882
rect 188482 51818 188534 51824
rect 188126 51734 188200 51762
rect 187942 51632 188108 51660
rect 187976 51536 188028 51542
rect 187896 51496 187976 51524
rect 187792 6860 187844 6866
rect 187792 6802 187844 6808
rect 187896 6798 187924 51496
rect 187976 51478 188028 51484
rect 187976 51400 188028 51406
rect 187976 51342 188028 51348
rect 187884 6792 187936 6798
rect 187884 6734 187936 6740
rect 187988 6662 188016 51342
rect 188080 50250 188108 51632
rect 188068 50244 188120 50250
rect 188068 50186 188120 50192
rect 188068 49700 188120 49706
rect 188068 49642 188120 49648
rect 188080 49094 188108 49642
rect 188068 49088 188120 49094
rect 188068 49030 188120 49036
rect 188068 46232 188120 46238
rect 188068 46174 188120 46180
rect 187976 6656 188028 6662
rect 187976 6598 188028 6604
rect 188080 6458 188108 46174
rect 188172 9450 188200 51734
rect 188264 51734 188430 51762
rect 188264 32434 188292 51734
rect 188344 51672 188396 51678
rect 188586 51626 188614 52020
rect 188678 51814 188706 52020
rect 188666 51808 188718 51814
rect 188666 51750 188718 51756
rect 188770 51660 188798 52020
rect 188862 51921 188890 52020
rect 188848 51912 188904 51921
rect 188954 51882 188982 52020
rect 188848 51847 188904 51856
rect 188942 51876 188994 51882
rect 188942 51818 188994 51824
rect 189046 51762 189074 52020
rect 188344 51614 188396 51620
rect 188356 50318 188384 51614
rect 188540 51598 188614 51626
rect 188724 51632 188798 51660
rect 189000 51734 189074 51762
rect 188436 51332 188488 51338
rect 188436 51274 188488 51280
rect 188344 50312 188396 50318
rect 188344 50254 188396 50260
rect 188448 46714 188476 51274
rect 188436 46708 188488 46714
rect 188436 46650 188488 46656
rect 188540 46594 188568 51598
rect 188724 50658 188752 51632
rect 188896 51468 188948 51474
rect 188896 51410 188948 51416
rect 188908 51134 188936 51410
rect 188896 51128 188948 51134
rect 188896 51070 188948 51076
rect 188712 50652 188764 50658
rect 188712 50594 188764 50600
rect 188896 50652 188948 50658
rect 188896 50594 188948 50600
rect 188712 50448 188764 50454
rect 188712 50390 188764 50396
rect 188620 48680 188672 48686
rect 188620 48622 188672 48628
rect 188448 46566 188568 46594
rect 188448 45014 188476 46566
rect 188528 46300 188580 46306
rect 188528 46242 188580 46248
rect 188436 45008 188488 45014
rect 188436 44950 188488 44956
rect 188252 32428 188304 32434
rect 188252 32370 188304 32376
rect 188160 9444 188212 9450
rect 188160 9386 188212 9392
rect 188540 6914 188568 46242
rect 188448 6886 188568 6914
rect 188068 6452 188120 6458
rect 188068 6394 188120 6400
rect 188448 3398 188476 6886
rect 188528 5568 188580 5574
rect 188528 5510 188580 5516
rect 188436 3392 188488 3398
rect 188436 3334 188488 3340
rect 188540 480 188568 5510
rect 188632 3738 188660 48622
rect 188724 46238 188752 50390
rect 188804 50244 188856 50250
rect 188804 50186 188856 50192
rect 188712 46232 188764 46238
rect 188712 46174 188764 46180
rect 188620 3732 188672 3738
rect 188620 3674 188672 3680
rect 188816 3670 188844 50186
rect 188908 48657 188936 50594
rect 188894 48648 188950 48657
rect 188894 48583 188950 48592
rect 189000 48385 189028 51734
rect 189138 51660 189166 52020
rect 189230 51950 189258 52020
rect 189218 51944 189270 51950
rect 189218 51886 189270 51892
rect 189092 51632 189166 51660
rect 189322 51660 189350 52020
rect 189414 51864 189442 52020
rect 189598 51882 189626 52020
rect 189586 51876 189638 51882
rect 189414 51836 189534 51864
rect 189506 51762 189534 51836
rect 189586 51818 189638 51824
rect 189690 51762 189718 52020
rect 189782 51882 189810 52020
rect 189770 51876 189822 51882
rect 189770 51818 189822 51824
rect 189874 51762 189902 52020
rect 189506 51734 189580 51762
rect 189448 51672 189500 51678
rect 189322 51632 189396 51660
rect 188986 48376 189042 48385
rect 188986 48311 189042 48320
rect 188804 3664 188856 3670
rect 188804 3606 188856 3612
rect 189092 3602 189120 51632
rect 189172 51536 189224 51542
rect 189172 51478 189224 51484
rect 189264 51536 189316 51542
rect 189264 51478 189316 51484
rect 189184 50658 189212 51478
rect 189172 50652 189224 50658
rect 189172 50594 189224 50600
rect 189276 50017 189304 51478
rect 189262 50008 189318 50017
rect 189262 49943 189318 49952
rect 189368 47462 189396 51632
rect 189448 51614 189500 51620
rect 189356 47456 189408 47462
rect 189356 47398 189408 47404
rect 189460 47326 189488 51614
rect 189448 47320 189500 47326
rect 189448 47262 189500 47268
rect 189552 46646 189580 51734
rect 189644 51734 189718 51762
rect 189828 51734 189902 51762
rect 189540 46640 189592 46646
rect 189540 46582 189592 46588
rect 189644 46186 189672 51734
rect 189724 51672 189776 51678
rect 189724 51614 189776 51620
rect 189736 48385 189764 51614
rect 189722 48376 189778 48385
rect 189722 48311 189778 48320
rect 189828 47274 189856 51734
rect 189966 51660 189994 52020
rect 189920 51632 189994 51660
rect 190058 51660 190086 52020
rect 190150 51950 190178 52020
rect 190242 51950 190270 52020
rect 190138 51944 190190 51950
rect 190138 51886 190190 51892
rect 190230 51944 190282 51950
rect 190334 51932 190362 52020
rect 190334 51904 190408 51932
rect 190230 51886 190282 51892
rect 190380 51864 190408 51904
rect 190334 51836 190408 51864
rect 190184 51808 190236 51814
rect 190184 51750 190236 51756
rect 190058 51632 190132 51660
rect 189920 48006 189948 51632
rect 190104 51074 190132 51632
rect 190012 51046 190132 51074
rect 189908 48000 189960 48006
rect 189908 47942 189960 47948
rect 189828 47246 189948 47274
rect 189184 46158 189672 46186
rect 189184 9382 189212 46158
rect 189264 46096 189316 46102
rect 189264 46038 189316 46044
rect 189276 15910 189304 46038
rect 189814 45520 189870 45529
rect 189814 45455 189870 45464
rect 189724 45280 189776 45286
rect 189724 45222 189776 45228
rect 189264 15904 189316 15910
rect 189264 15846 189316 15852
rect 189172 9376 189224 9382
rect 189172 9318 189224 9324
rect 189736 4146 189764 45222
rect 189724 4140 189776 4146
rect 189724 4082 189776 4088
rect 189080 3596 189132 3602
rect 189080 3538 189132 3544
rect 189828 3534 189856 45455
rect 189920 43586 189948 47246
rect 190012 46102 190040 51046
rect 190196 50182 190224 51750
rect 190334 51660 190362 51836
rect 190518 51762 190546 52020
rect 190288 51632 190362 51660
rect 190472 51734 190546 51762
rect 190184 50176 190236 50182
rect 190184 50118 190236 50124
rect 190184 47320 190236 47326
rect 190184 47262 190236 47268
rect 190092 46980 190144 46986
rect 190092 46922 190144 46928
rect 190000 46096 190052 46102
rect 190000 46038 190052 46044
rect 190104 45914 190132 46922
rect 190012 45886 190132 45914
rect 189908 43580 189960 43586
rect 189908 43522 189960 43528
rect 189908 42832 189960 42838
rect 189908 42774 189960 42780
rect 189816 3528 189868 3534
rect 189816 3470 189868 3476
rect 189724 3324 189776 3330
rect 189724 3266 189776 3272
rect 189736 480 189764 3266
rect 189920 3194 189948 42774
rect 190012 4078 190040 45886
rect 190090 44432 190146 44441
rect 190090 44367 190146 44376
rect 190000 4072 190052 4078
rect 190000 4014 190052 4020
rect 190104 3262 190132 44367
rect 190196 43654 190224 47262
rect 190288 44946 190316 51632
rect 190368 51536 190420 51542
rect 190368 51478 190420 51484
rect 190380 50658 190408 51478
rect 190368 50652 190420 50658
rect 190368 50594 190420 50600
rect 190368 50176 190420 50182
rect 190368 50118 190420 50124
rect 190380 47938 190408 50118
rect 190368 47932 190420 47938
rect 190368 47874 190420 47880
rect 190472 47870 190500 51734
rect 190610 51660 190638 52020
rect 190702 51762 190730 52020
rect 190794 51882 190822 52020
rect 190886 51882 190914 52020
rect 190782 51876 190834 51882
rect 190782 51818 190834 51824
rect 190874 51876 190926 51882
rect 190874 51818 190926 51824
rect 190978 51762 191006 52020
rect 190702 51734 190776 51762
rect 190610 51632 190684 51660
rect 190552 51536 190604 51542
rect 190552 51478 190604 51484
rect 190460 47864 190512 47870
rect 190460 47806 190512 47812
rect 190368 47456 190420 47462
rect 190368 47398 190420 47404
rect 190276 44940 190328 44946
rect 190276 44882 190328 44888
rect 190380 43722 190408 47398
rect 190460 46368 190512 46374
rect 190460 46310 190512 46316
rect 190368 43716 190420 43722
rect 190368 43658 190420 43664
rect 190184 43648 190236 43654
rect 190184 43590 190236 43596
rect 190472 41414 190500 46310
rect 190564 46186 190592 51478
rect 190656 50386 190684 51632
rect 190644 50380 190696 50386
rect 190644 50322 190696 50328
rect 190644 48068 190696 48074
rect 190644 48010 190696 48016
rect 190656 46458 190684 48010
rect 190748 47682 190776 51734
rect 190932 51734 191006 51762
rect 190828 51468 190880 51474
rect 190828 51410 190880 51416
rect 190840 48074 190868 51410
rect 190932 48074 190960 51734
rect 191070 51660 191098 52020
rect 191162 51762 191190 52020
rect 191254 51882 191282 52020
rect 191346 51950 191374 52020
rect 191334 51944 191386 51950
rect 191334 51886 191386 51892
rect 191242 51876 191294 51882
rect 191242 51818 191294 51824
rect 191438 51762 191466 52020
rect 191162 51734 191236 51762
rect 191024 51632 191098 51660
rect 190828 48068 190880 48074
rect 190828 48010 190880 48016
rect 190920 48068 190972 48074
rect 190920 48010 190972 48016
rect 190748 47654 190960 47682
rect 190656 46430 190868 46458
rect 190736 46300 190788 46306
rect 190736 46242 190788 46248
rect 190564 46158 190684 46186
rect 190472 41386 190592 41414
rect 190564 4049 190592 41386
rect 190656 20602 190684 46158
rect 190644 20596 190696 20602
rect 190644 20538 190696 20544
rect 190550 4040 190606 4049
rect 190550 3975 190606 3984
rect 190748 3913 190776 46242
rect 190840 21690 190868 46430
rect 190932 44878 190960 47654
rect 191024 46578 191052 51632
rect 191104 51536 191156 51542
rect 191104 51478 191156 51484
rect 191012 46572 191064 46578
rect 191012 46514 191064 46520
rect 191012 46436 191064 46442
rect 191012 46378 191064 46384
rect 191024 46050 191052 46378
rect 191116 46186 191144 51478
rect 191208 46374 191236 51734
rect 191300 51734 191466 51762
rect 191530 51762 191558 52020
rect 191622 51950 191650 52020
rect 191610 51944 191662 51950
rect 191610 51886 191662 51892
rect 191714 51882 191742 52020
rect 191702 51876 191754 51882
rect 191702 51818 191754 51824
rect 191806 51814 191834 52020
rect 191898 51814 191926 52020
rect 191990 51814 192018 52020
rect 192082 51950 192110 52020
rect 192070 51944 192122 51950
rect 192070 51886 192122 51892
rect 192174 51864 192202 52020
rect 192174 51836 192248 51864
rect 191794 51808 191846 51814
rect 191530 51734 191604 51762
rect 191794 51750 191846 51756
rect 191886 51808 191938 51814
rect 191886 51750 191938 51756
rect 191978 51808 192030 51814
rect 191978 51750 192030 51756
rect 191196 46368 191248 46374
rect 191196 46310 191248 46316
rect 191300 46306 191328 51734
rect 191576 51490 191604 51734
rect 192116 51740 192168 51746
rect 192116 51682 192168 51688
rect 191748 51604 191800 51610
rect 191748 51546 191800 51552
rect 191840 51604 191892 51610
rect 191840 51546 191892 51552
rect 192024 51604 192076 51610
rect 192024 51546 192076 51552
rect 191380 51468 191432 51474
rect 191380 51410 191432 51416
rect 191484 51462 191604 51490
rect 191656 51536 191708 51542
rect 191656 51478 191708 51484
rect 191392 50017 191420 51410
rect 191378 50008 191434 50017
rect 191378 49943 191434 49952
rect 191484 49881 191512 51462
rect 191564 51400 191616 51406
rect 191564 51342 191616 51348
rect 191470 49872 191526 49881
rect 191470 49807 191526 49816
rect 191380 48068 191432 48074
rect 191380 48010 191432 48016
rect 191288 46300 191340 46306
rect 191288 46242 191340 46248
rect 191116 46158 191328 46186
rect 191024 46022 191236 46050
rect 190920 44872 190972 44878
rect 190920 44814 190972 44820
rect 191104 44124 191156 44130
rect 191104 44066 191156 44072
rect 190828 21684 190880 21690
rect 190828 21626 190880 21632
rect 190828 4140 190880 4146
rect 190828 4082 190880 4088
rect 190734 3904 190790 3913
rect 190734 3839 190790 3848
rect 190092 3256 190144 3262
rect 190092 3198 190144 3204
rect 189908 3188 189960 3194
rect 189908 3130 189960 3136
rect 190840 480 190868 4082
rect 191116 3398 191144 44066
rect 191208 4010 191236 46022
rect 191300 41414 191328 46158
rect 191392 43518 191420 48010
rect 191576 47598 191604 51342
rect 191668 50017 191696 51478
rect 191760 50153 191788 51546
rect 191746 50144 191802 50153
rect 191746 50079 191802 50088
rect 191654 50008 191710 50017
rect 191654 49943 191710 49952
rect 191564 47592 191616 47598
rect 191564 47534 191616 47540
rect 191380 43512 191432 43518
rect 191380 43454 191432 43460
rect 191300 41386 191512 41414
rect 191196 4004 191248 4010
rect 191196 3946 191248 3952
rect 191484 3466 191512 41386
rect 191852 6730 191880 51546
rect 191932 51468 191984 51474
rect 191932 51410 191984 51416
rect 191944 47734 191972 51410
rect 191932 47728 191984 47734
rect 191932 47670 191984 47676
rect 192036 47666 192064 51546
rect 192024 47660 192076 47666
rect 192024 47602 192076 47608
rect 192024 43036 192076 43042
rect 192024 42978 192076 42984
rect 192036 13138 192064 42978
rect 192128 13326 192156 51682
rect 192220 19242 192248 51836
rect 192358 51762 192386 52020
rect 192312 51734 192386 51762
rect 192312 43042 192340 51734
rect 192450 51660 192478 52020
rect 192542 51955 192570 52020
rect 192528 51946 192584 51955
rect 192634 51950 192662 52020
rect 192528 51881 192584 51890
rect 192622 51944 192674 51950
rect 192622 51886 192674 51892
rect 192576 51808 192628 51814
rect 192726 51762 192754 52020
rect 192576 51750 192628 51756
rect 192404 51632 192478 51660
rect 192300 43036 192352 43042
rect 192300 42978 192352 42984
rect 192300 42900 192352 42906
rect 192300 42842 192352 42848
rect 192208 19236 192260 19242
rect 192208 19178 192260 19184
rect 192312 19106 192340 42842
rect 192404 19174 192432 51632
rect 192484 46232 192536 46238
rect 192484 46174 192536 46180
rect 192496 28626 192524 46174
rect 192588 41414 192616 51750
rect 192680 51734 192754 51762
rect 192680 42906 192708 51734
rect 192818 51660 192846 52020
rect 192910 51921 192938 52020
rect 192896 51912 192952 51921
rect 192896 51847 192952 51856
rect 192772 51632 192846 51660
rect 193002 51660 193030 52020
rect 193094 51762 193122 52020
rect 193186 51882 193214 52020
rect 193174 51876 193226 51882
rect 193174 51818 193226 51824
rect 193278 51762 193306 52020
rect 193370 51921 193398 52020
rect 193356 51912 193412 51921
rect 193462 51882 193490 52020
rect 193554 51955 193582 52020
rect 193540 51946 193596 51955
rect 193356 51847 193412 51856
rect 193450 51876 193502 51882
rect 193540 51881 193596 51890
rect 193450 51818 193502 51824
rect 193094 51734 193168 51762
rect 193278 51734 193352 51762
rect 193002 51632 193076 51660
rect 192772 46238 192800 51632
rect 192944 51536 192996 51542
rect 192944 51478 192996 51484
rect 192956 48793 192984 51478
rect 192942 48784 192998 48793
rect 192942 48719 192998 48728
rect 193048 48521 193076 51632
rect 193140 48657 193168 51734
rect 193126 48648 193182 48657
rect 193126 48583 193182 48592
rect 193034 48512 193090 48521
rect 193034 48447 193090 48456
rect 193220 47524 193272 47530
rect 193220 47466 193272 47472
rect 192760 46232 192812 46238
rect 192760 46174 192812 46180
rect 192668 42900 192720 42906
rect 192668 42842 192720 42848
rect 192588 41386 192800 41414
rect 192484 28620 192536 28626
rect 192484 28562 192536 28568
rect 192392 19168 192444 19174
rect 192392 19110 192444 19116
rect 192300 19100 192352 19106
rect 192300 19042 192352 19048
rect 192116 13320 192168 13326
rect 192116 13262 192168 13268
rect 192036 13110 192156 13138
rect 192024 12436 192076 12442
rect 192024 12378 192076 12384
rect 191840 6724 191892 6730
rect 191840 6666 191892 6672
rect 191472 3460 191524 3466
rect 191472 3402 191524 3408
rect 191104 3392 191156 3398
rect 191104 3334 191156 3340
rect 192036 480 192064 12378
rect 192128 11694 192156 13110
rect 192116 11688 192168 11694
rect 192116 11630 192168 11636
rect 192772 10606 192800 41386
rect 192760 10600 192812 10606
rect 192760 10542 192812 10548
rect 193232 4146 193260 47466
rect 193324 46102 193352 51734
rect 193646 51592 193674 52020
rect 193738 51660 193766 52020
rect 193830 51728 193858 52020
rect 193922 51921 193950 52020
rect 194014 51950 194042 52020
rect 194106 51950 194134 52020
rect 194198 51950 194226 52020
rect 194290 51950 194318 52020
rect 194002 51944 194054 51950
rect 193908 51912 193964 51921
rect 194002 51886 194054 51892
rect 194094 51944 194146 51950
rect 194094 51886 194146 51892
rect 194186 51944 194238 51950
rect 194186 51886 194238 51892
rect 194278 51944 194330 51950
rect 194278 51886 194330 51892
rect 194382 51882 194410 52020
rect 194474 51882 194502 52020
rect 193908 51847 193964 51856
rect 194370 51876 194422 51882
rect 194370 51818 194422 51824
rect 194462 51876 194514 51882
rect 194462 51818 194514 51824
rect 194048 51740 194100 51746
rect 193830 51700 193996 51728
rect 193738 51632 193812 51660
rect 193646 51564 193720 51592
rect 193404 50176 193456 50182
rect 193404 50118 193456 50124
rect 193312 46096 193364 46102
rect 193312 46038 193364 46044
rect 193312 45960 193364 45966
rect 193312 45902 193364 45908
rect 193324 6594 193352 45902
rect 193416 41414 193444 50118
rect 193692 49434 193720 51564
rect 193680 49428 193732 49434
rect 193680 49370 193732 49376
rect 193680 47456 193732 47462
rect 193586 47424 193642 47433
rect 193680 47398 193732 47404
rect 193586 47359 193642 47368
rect 193416 41386 193536 41414
rect 193508 18970 193536 41386
rect 193600 19038 193628 47359
rect 193692 23390 193720 47398
rect 193784 27266 193812 51632
rect 193968 50182 193996 51700
rect 194048 51682 194100 51688
rect 194140 51740 194192 51746
rect 194140 51682 194192 51688
rect 194244 51734 194410 51762
rect 193956 50176 194008 50182
rect 193956 50118 194008 50124
rect 193862 50008 193918 50017
rect 193862 49943 193918 49952
rect 193876 47530 193904 49943
rect 193864 47524 193916 47530
rect 193864 47466 193916 47472
rect 194060 47410 194088 51682
rect 193876 47382 194088 47410
rect 193876 35494 193904 47382
rect 193956 46096 194008 46102
rect 193956 46038 194008 46044
rect 193968 40866 193996 46038
rect 194152 45966 194180 51682
rect 194244 50153 194272 51734
rect 194382 51728 194410 51734
rect 194566 51728 194594 52020
rect 194382 51700 194594 51728
rect 194658 51728 194686 52020
rect 194750 51950 194778 52020
rect 194738 51944 194790 51950
rect 194842 51921 194870 52020
rect 194934 51950 194962 52020
rect 194922 51944 194974 51950
rect 194738 51886 194790 51892
rect 194828 51912 194884 51921
rect 194922 51886 194974 51892
rect 194828 51847 194884 51856
rect 194784 51808 194836 51814
rect 194784 51750 194836 51756
rect 195026 51762 195054 52020
rect 195118 51921 195146 52020
rect 195210 51950 195238 52020
rect 195302 51950 195330 52020
rect 195394 51950 195422 52020
rect 195486 51955 195514 52020
rect 195198 51944 195250 51950
rect 195104 51912 195160 51921
rect 195198 51886 195250 51892
rect 195290 51944 195342 51950
rect 195290 51886 195342 51892
rect 195382 51944 195434 51950
rect 195382 51886 195434 51892
rect 195472 51946 195528 51955
rect 195578 51950 195606 52020
rect 195472 51881 195528 51890
rect 195566 51944 195618 51950
rect 195566 51886 195618 51892
rect 195670 51882 195698 52020
rect 195104 51847 195160 51856
rect 195658 51876 195710 51882
rect 195658 51818 195710 51824
rect 195762 51796 195790 52020
rect 195854 51955 195882 52020
rect 195840 51946 195896 51955
rect 195840 51881 195896 51890
rect 195762 51768 195836 51796
rect 194658 51700 194732 51728
rect 194324 51604 194376 51610
rect 194324 51546 194376 51552
rect 194416 51604 194468 51610
rect 194416 51546 194468 51552
rect 194230 50144 194286 50153
rect 194230 50079 194286 50088
rect 194336 47433 194364 51546
rect 194428 47569 194456 51546
rect 194600 51536 194652 51542
rect 194600 51478 194652 51484
rect 194508 51400 194560 51406
rect 194508 51342 194560 51348
rect 194414 47560 194470 47569
rect 194414 47495 194470 47504
rect 194322 47424 194378 47433
rect 194322 47359 194378 47368
rect 194140 45960 194192 45966
rect 194140 45902 194192 45908
rect 193956 40860 194008 40866
rect 193956 40802 194008 40808
rect 193864 35488 193916 35494
rect 193864 35430 193916 35436
rect 193772 27260 193824 27266
rect 193772 27202 193824 27208
rect 193680 23384 193732 23390
rect 193680 23326 193732 23332
rect 193680 22772 193732 22778
rect 193680 22714 193732 22720
rect 193588 19032 193640 19038
rect 193588 18974 193640 18980
rect 193496 18964 193548 18970
rect 193496 18906 193548 18912
rect 193692 16574 193720 22714
rect 193692 16546 194456 16574
rect 193312 6588 193364 6594
rect 193312 6530 193364 6536
rect 193220 4140 193272 4146
rect 193220 4082 193272 4088
rect 193220 3188 193272 3194
rect 193220 3130 193272 3136
rect 193232 480 193260 3130
rect 194428 480 194456 16546
rect 194520 10538 194548 51342
rect 194612 47462 194640 51478
rect 194704 51074 194732 51700
rect 194796 51406 194824 51750
rect 195026 51734 195192 51762
rect 195060 51672 195112 51678
rect 195060 51614 195112 51620
rect 194784 51400 194836 51406
rect 194784 51342 194836 51348
rect 194704 51046 195008 51074
rect 194690 47560 194746 47569
rect 194690 47495 194746 47504
rect 194600 47456 194652 47462
rect 194600 47398 194652 47404
rect 194508 10532 194560 10538
rect 194508 10474 194560 10480
rect 194600 10396 194652 10402
rect 194600 10338 194652 10344
rect 194612 490 194640 10338
rect 194704 6526 194732 47495
rect 194784 47456 194836 47462
rect 194784 47398 194836 47404
rect 194874 47424 194930 47433
rect 194796 8022 194824 47398
rect 194874 47359 194930 47368
rect 194888 17202 194916 47359
rect 194980 18902 195008 51046
rect 195072 24478 195100 51614
rect 195164 28490 195192 51734
rect 195336 51740 195388 51746
rect 195336 51682 195388 51688
rect 195244 51604 195296 51610
rect 195244 51546 195296 51552
rect 195256 28558 195284 51546
rect 195348 29986 195376 51682
rect 195428 51672 195480 51678
rect 195428 51614 195480 51620
rect 195612 51672 195664 51678
rect 195612 51614 195664 51620
rect 195440 31346 195468 51614
rect 195520 51604 195572 51610
rect 195520 51546 195572 51552
rect 195532 47462 195560 51546
rect 195624 47569 195652 51614
rect 195702 49736 195758 49745
rect 195702 49671 195758 49680
rect 195716 47802 195744 49671
rect 195704 47796 195756 47802
rect 195704 47738 195756 47744
rect 195610 47560 195666 47569
rect 195610 47495 195666 47504
rect 195520 47456 195572 47462
rect 195808 47433 195836 51768
rect 195946 51728 195974 52020
rect 196038 51950 196066 52020
rect 196026 51944 196078 51950
rect 196026 51886 196078 51892
rect 196130 51728 196158 52020
rect 196222 51950 196250 52020
rect 196210 51944 196262 51950
rect 196210 51886 196262 51892
rect 195900 51700 195974 51728
rect 196084 51700 196158 51728
rect 196314 51728 196342 52020
rect 196406 51796 196434 52020
rect 196498 51950 196526 52020
rect 196486 51944 196538 51950
rect 196590 51921 196618 52020
rect 196486 51886 196538 51892
rect 196576 51912 196632 51921
rect 196576 51847 196632 51856
rect 196682 51796 196710 52020
rect 196406 51768 196480 51796
rect 196314 51700 196388 51728
rect 195900 47705 195928 51700
rect 195980 51536 196032 51542
rect 195980 51478 196032 51484
rect 195886 47696 195942 47705
rect 195886 47631 195942 47640
rect 195520 47398 195572 47404
rect 195794 47424 195850 47433
rect 195794 47359 195850 47368
rect 195610 47288 195666 47297
rect 195610 47223 195666 47232
rect 195428 31340 195480 31346
rect 195428 31282 195480 31288
rect 195336 29980 195388 29986
rect 195336 29922 195388 29928
rect 195244 28552 195296 28558
rect 195244 28494 195296 28500
rect 195152 28484 195204 28490
rect 195152 28426 195204 28432
rect 195060 24472 195112 24478
rect 195060 24414 195112 24420
rect 194968 18896 195020 18902
rect 194968 18838 195020 18844
rect 194876 17196 194928 17202
rect 194876 17138 194928 17144
rect 194784 8016 194836 8022
rect 194784 7958 194836 7964
rect 194692 6520 194744 6526
rect 194692 6462 194744 6468
rect 195624 5166 195652 47223
rect 195612 5160 195664 5166
rect 195612 5102 195664 5108
rect 195992 5098 196020 51478
rect 196084 48482 196112 51700
rect 196360 50130 196388 51700
rect 196452 50590 196480 51768
rect 196636 51768 196710 51796
rect 196532 51672 196584 51678
rect 196532 51614 196584 51620
rect 196440 50584 196492 50590
rect 196440 50526 196492 50532
rect 196176 50102 196388 50130
rect 196072 48476 196124 48482
rect 196072 48418 196124 48424
rect 196176 48074 196204 50102
rect 196346 49736 196402 49745
rect 196346 49671 196402 49680
rect 196256 48816 196308 48822
rect 196256 48758 196308 48764
rect 196164 48068 196216 48074
rect 196164 48010 196216 48016
rect 196164 47456 196216 47462
rect 196164 47398 196216 47404
rect 196070 21448 196126 21457
rect 196070 21383 196126 21392
rect 196084 6914 196112 21383
rect 196176 15094 196204 47398
rect 196164 15088 196216 15094
rect 196164 15030 196216 15036
rect 196268 14346 196296 48758
rect 196360 18834 196388 49671
rect 196544 48822 196572 51614
rect 196532 48816 196584 48822
rect 196532 48758 196584 48764
rect 196532 48340 196584 48346
rect 196532 48282 196584 48288
rect 196440 48068 196492 48074
rect 196440 48010 196492 48016
rect 196452 23322 196480 48010
rect 196544 25770 196572 48282
rect 196636 31278 196664 51768
rect 196774 51728 196802 52020
rect 196866 51950 196894 52020
rect 196854 51944 196906 51950
rect 196854 51886 196906 51892
rect 196728 51700 196802 51728
rect 196958 51728 196986 52020
rect 197050 51796 197078 52020
rect 197142 51921 197170 52020
rect 197234 51950 197262 52020
rect 197326 51950 197354 52020
rect 197222 51944 197274 51950
rect 197128 51912 197184 51921
rect 197222 51886 197274 51892
rect 197314 51944 197366 51950
rect 197314 51886 197366 51892
rect 197418 51882 197446 52020
rect 197510 51882 197538 52020
rect 197128 51847 197184 51856
rect 197406 51876 197458 51882
rect 197406 51818 197458 51824
rect 197498 51876 197550 51882
rect 197498 51818 197550 51824
rect 197050 51768 197124 51796
rect 196958 51700 197032 51728
rect 196728 51610 196756 51700
rect 196716 51604 196768 51610
rect 196716 51546 196768 51552
rect 196808 51536 196860 51542
rect 196808 51478 196860 51484
rect 196900 51536 196952 51542
rect 196900 51478 196952 51484
rect 196716 51468 196768 51474
rect 196716 51410 196768 51416
rect 196728 33862 196756 51410
rect 196820 38350 196848 51478
rect 196912 45554 196940 51478
rect 197004 48346 197032 51700
rect 196992 48340 197044 48346
rect 196992 48282 197044 48288
rect 197096 47462 197124 51768
rect 197268 51740 197320 51746
rect 197268 51682 197320 51688
rect 197360 51740 197412 51746
rect 197602 51728 197630 52020
rect 197694 51950 197722 52020
rect 197682 51944 197734 51950
rect 197682 51886 197734 51892
rect 197786 51728 197814 52020
rect 197878 51882 197906 52020
rect 197866 51876 197918 51882
rect 197866 51818 197918 51824
rect 197970 51814 197998 52020
rect 198062 51950 198090 52020
rect 198050 51944 198102 51950
rect 198050 51886 198102 51892
rect 197958 51808 198010 51814
rect 198154 51796 198182 52020
rect 197958 51750 198010 51756
rect 198108 51768 198182 51796
rect 197602 51700 197676 51728
rect 197786 51700 197860 51728
rect 197360 51682 197412 51688
rect 197176 51604 197228 51610
rect 197176 51546 197228 51552
rect 197084 47456 197136 47462
rect 197084 47398 197136 47404
rect 196912 45526 197124 45554
rect 197096 43382 197124 45526
rect 197084 43376 197136 43382
rect 197084 43318 197136 43324
rect 196808 38344 196860 38350
rect 196808 38286 196860 38292
rect 196716 33856 196768 33862
rect 196716 33798 196768 33804
rect 196624 31272 196676 31278
rect 196624 31214 196676 31220
rect 196532 25764 196584 25770
rect 196532 25706 196584 25712
rect 196440 23316 196492 23322
rect 196440 23258 196492 23264
rect 196348 18828 196400 18834
rect 196348 18770 196400 18776
rect 197188 14414 197216 51546
rect 197280 48657 197308 51682
rect 197372 48686 197400 51682
rect 197544 51604 197596 51610
rect 197544 51546 197596 51552
rect 197556 50454 197584 51546
rect 197544 50448 197596 50454
rect 197544 50390 197596 50396
rect 197544 48952 197596 48958
rect 197544 48894 197596 48900
rect 197360 48680 197412 48686
rect 197266 48648 197322 48657
rect 197360 48622 197412 48628
rect 197266 48583 197322 48592
rect 197360 46164 197412 46170
rect 197360 46106 197412 46112
rect 197176 14408 197228 14414
rect 197176 14350 197228 14356
rect 196256 14340 196308 14346
rect 196256 14282 196308 14288
rect 197372 7886 197400 46106
rect 197556 45554 197584 48894
rect 197464 45526 197584 45554
rect 197464 7954 197492 45526
rect 197544 43376 197596 43382
rect 197544 43318 197596 43324
rect 197556 9654 197584 43318
rect 197648 15026 197676 51700
rect 197832 51626 197860 51700
rect 198004 51672 198056 51678
rect 197728 51604 197780 51610
rect 197832 51598 197952 51626
rect 198004 51614 198056 51620
rect 197728 51546 197780 51552
rect 197636 15020 197688 15026
rect 197636 14962 197688 14968
rect 197740 14958 197768 51546
rect 197820 51536 197872 51542
rect 197820 51478 197872 51484
rect 197832 23254 197860 51478
rect 197924 27198 197952 51598
rect 198016 48770 198044 51614
rect 198108 48958 198136 51768
rect 198246 51728 198274 52020
rect 198200 51700 198274 51728
rect 198338 51728 198366 52020
rect 198430 51921 198458 52020
rect 198416 51912 198472 51921
rect 198416 51847 198472 51856
rect 198522 51814 198550 52020
rect 198614 51955 198642 52020
rect 198600 51946 198656 51955
rect 198600 51881 198656 51890
rect 198510 51808 198562 51814
rect 198706 51762 198734 52020
rect 198798 51882 198826 52020
rect 198786 51876 198838 51882
rect 198786 51818 198838 51824
rect 198890 51762 198918 52020
rect 198510 51750 198562 51756
rect 198660 51734 198734 51762
rect 198844 51734 198918 51762
rect 198338 51700 198412 51728
rect 198096 48952 198148 48958
rect 198096 48894 198148 48900
rect 198016 48742 198136 48770
rect 198004 48680 198056 48686
rect 198004 48622 198056 48628
rect 198016 29918 198044 48622
rect 198108 39574 198136 48742
rect 198200 40798 198228 51700
rect 198280 51604 198332 51610
rect 198280 51546 198332 51552
rect 198292 48414 198320 51546
rect 198280 48408 198332 48414
rect 198280 48350 198332 48356
rect 198384 46170 198412 51700
rect 198464 51672 198516 51678
rect 198464 51614 198516 51620
rect 198476 48929 198504 51614
rect 198660 51610 198688 51734
rect 198740 51672 198792 51678
rect 198740 51614 198792 51620
rect 198648 51604 198700 51610
rect 198648 51546 198700 51552
rect 198556 51468 198608 51474
rect 198556 51410 198608 51416
rect 198462 48920 198518 48929
rect 198462 48855 198518 48864
rect 198568 48657 198596 51410
rect 198554 48648 198610 48657
rect 198554 48583 198610 48592
rect 198372 46164 198424 46170
rect 198372 46106 198424 46112
rect 198752 45898 198780 51614
rect 198844 47122 198872 51734
rect 198982 51660 199010 52020
rect 199074 51950 199102 52020
rect 199062 51944 199114 51950
rect 199062 51886 199114 51892
rect 199166 51762 199194 52020
rect 198936 51632 199010 51660
rect 199120 51734 199194 51762
rect 199258 51762 199286 52020
rect 199350 51882 199378 52020
rect 199338 51876 199390 51882
rect 199338 51818 199390 51824
rect 199442 51762 199470 52020
rect 199534 51882 199562 52020
rect 199522 51876 199574 51882
rect 199522 51818 199574 51824
rect 199626 51762 199654 52020
rect 199258 51734 199332 51762
rect 199442 51734 199516 51762
rect 198832 47116 198884 47122
rect 198832 47058 198884 47064
rect 198832 46028 198884 46034
rect 198832 45970 198884 45976
rect 198740 45892 198792 45898
rect 198740 45834 198792 45840
rect 198740 45756 198792 45762
rect 198740 45698 198792 45704
rect 198188 40792 198240 40798
rect 198188 40734 198240 40740
rect 198096 39568 198148 39574
rect 198096 39510 198148 39516
rect 198004 29912 198056 29918
rect 198004 29854 198056 29860
rect 197912 27192 197964 27198
rect 197912 27134 197964 27140
rect 197820 23248 197872 23254
rect 197820 23190 197872 23196
rect 197728 14952 197780 14958
rect 197728 14894 197780 14900
rect 197544 9648 197596 9654
rect 197544 9590 197596 9596
rect 197452 7948 197504 7954
rect 197452 7890 197504 7896
rect 197360 7880 197412 7886
rect 197360 7822 197412 7828
rect 196084 6886 196848 6914
rect 195980 5092 196032 5098
rect 195980 5034 196032 5040
rect 187302 354 187414 480
rect 186884 326 187414 354
rect 187302 -960 187414 326
rect 188498 -960 188610 480
rect 189694 -960 189806 480
rect 190798 -960 190910 480
rect 191994 -960 192106 480
rect 193190 -960 193302 480
rect 194386 -960 194498 480
rect 194612 462 195192 490
rect 196820 480 196848 6886
rect 198752 5030 198780 45698
rect 198844 7818 198872 45970
rect 198936 9518 198964 51632
rect 199016 51536 199068 51542
rect 199016 51478 199068 51484
rect 199028 48385 199056 51478
rect 199014 48376 199070 48385
rect 199014 48311 199070 48320
rect 199120 46220 199148 51734
rect 199200 51672 199252 51678
rect 199200 51614 199252 51620
rect 199212 48686 199240 51614
rect 199200 48680 199252 48686
rect 199200 48622 199252 48628
rect 199200 47116 199252 47122
rect 199200 47058 199252 47064
rect 199028 46192 199148 46220
rect 199028 24410 199056 46192
rect 199108 46096 199160 46102
rect 199108 46038 199160 46044
rect 199120 25702 199148 46038
rect 199212 28422 199240 47058
rect 199304 35426 199332 51734
rect 199384 51604 199436 51610
rect 199384 51546 199436 51552
rect 199396 39370 199424 51546
rect 199488 46034 199516 51734
rect 199580 51734 199654 51762
rect 199718 51762 199746 52020
rect 199810 51882 199838 52020
rect 199798 51876 199850 51882
rect 199798 51818 199850 51824
rect 199902 51762 199930 52020
rect 199994 51882 200022 52020
rect 200086 51882 200114 52020
rect 199982 51876 200034 51882
rect 199982 51818 200034 51824
rect 200074 51876 200126 51882
rect 200074 51818 200126 51824
rect 200178 51762 200206 52020
rect 200362 51932 200390 52020
rect 199718 51734 199792 51762
rect 199902 51734 200068 51762
rect 199580 46102 199608 51734
rect 199660 51672 199712 51678
rect 199660 51614 199712 51620
rect 199568 46096 199620 46102
rect 199568 46038 199620 46044
rect 199476 46028 199528 46034
rect 199476 45970 199528 45976
rect 199476 45892 199528 45898
rect 199476 45834 199528 45840
rect 199488 39506 199516 45834
rect 199672 45762 199700 51614
rect 199764 48385 199792 51734
rect 199844 51672 199896 51678
rect 199844 51614 199896 51620
rect 199936 51672 199988 51678
rect 199936 51614 199988 51620
rect 199856 48657 199884 51614
rect 199842 48648 199898 48657
rect 199842 48583 199898 48592
rect 199948 48521 199976 51614
rect 200040 48754 200068 51734
rect 200132 51734 200206 51762
rect 200316 51904 200390 51932
rect 200028 48748 200080 48754
rect 200028 48690 200080 48696
rect 199934 48512 199990 48521
rect 199844 48476 199896 48482
rect 200132 48482 200160 51734
rect 200212 51672 200264 51678
rect 200212 51614 200264 51620
rect 199934 48447 199990 48456
rect 200120 48476 200172 48482
rect 199844 48418 199896 48424
rect 200120 48418 200172 48424
rect 199750 48376 199806 48385
rect 199750 48311 199806 48320
rect 199660 45756 199712 45762
rect 199660 45698 199712 45704
rect 199856 41414 199884 48418
rect 200224 46220 200252 51614
rect 200132 46192 200252 46220
rect 199580 41386 199884 41414
rect 200026 41440 200082 41449
rect 199476 39500 199528 39506
rect 199476 39442 199528 39448
rect 199384 39364 199436 39370
rect 199384 39306 199436 39312
rect 199292 35420 199344 35426
rect 199292 35362 199344 35368
rect 199580 33930 199608 41386
rect 200026 41375 200082 41384
rect 200040 36009 200068 41375
rect 200026 36000 200082 36009
rect 200026 35935 200082 35944
rect 199568 33924 199620 33930
rect 199568 33866 199620 33872
rect 199200 28416 199252 28422
rect 199200 28358 199252 28364
rect 199108 25696 199160 25702
rect 199108 25638 199160 25644
rect 199016 24404 199068 24410
rect 199016 24346 199068 24352
rect 198924 9512 198976 9518
rect 198924 9454 198976 9460
rect 200132 9314 200160 46192
rect 200212 46096 200264 46102
rect 200212 46038 200264 46044
rect 200120 9308 200172 9314
rect 200120 9250 200172 9256
rect 200224 9246 200252 46038
rect 200316 46034 200344 51904
rect 200454 51864 200482 52020
rect 200408 51836 200482 51864
rect 200304 46028 200356 46034
rect 200304 45970 200356 45976
rect 200304 45892 200356 45898
rect 200304 45834 200356 45840
rect 200316 12306 200344 45834
rect 200408 20398 200436 51836
rect 200546 51762 200574 52020
rect 200500 51734 200574 51762
rect 200500 50522 200528 51734
rect 200638 51660 200666 52020
rect 200730 51882 200758 52020
rect 200718 51876 200770 51882
rect 200718 51818 200770 51824
rect 200822 51762 200850 52020
rect 200592 51632 200666 51660
rect 200776 51734 200850 51762
rect 200488 50516 200540 50522
rect 200488 50458 200540 50464
rect 200592 46220 200620 51632
rect 200500 46192 200620 46220
rect 200500 24342 200528 46192
rect 200776 46152 200804 51734
rect 200914 51660 200942 52020
rect 201006 51728 201034 52020
rect 201098 51882 201126 52020
rect 201086 51876 201138 51882
rect 201086 51818 201138 51824
rect 201190 51796 201218 52020
rect 201282 51921 201310 52020
rect 201268 51912 201324 51921
rect 201268 51847 201324 51856
rect 201190 51768 201264 51796
rect 201006 51700 201172 51728
rect 200592 46124 200804 46152
rect 200868 51632 200942 51660
rect 200592 25634 200620 46124
rect 200672 46028 200724 46034
rect 200672 45970 200724 45976
rect 200764 46028 200816 46034
rect 200764 45970 200816 45976
rect 200684 27130 200712 45970
rect 200776 28354 200804 45970
rect 200868 37126 200896 51632
rect 201040 51604 201092 51610
rect 201040 51546 201092 51552
rect 200948 51536 201000 51542
rect 200948 51478 201000 51484
rect 200960 40730 200988 51478
rect 201052 49842 201080 51546
rect 201040 49836 201092 49842
rect 201040 49778 201092 49784
rect 201144 46034 201172 51700
rect 201132 46028 201184 46034
rect 201132 45970 201184 45976
rect 201236 45898 201264 51768
rect 201374 51762 201402 52020
rect 201328 51734 201402 51762
rect 201328 46102 201356 51734
rect 201466 51660 201494 52020
rect 201420 51632 201494 51660
rect 201420 48385 201448 51632
rect 201558 51524 201586 52020
rect 201650 51814 201678 52020
rect 201742 51950 201770 52020
rect 201834 51955 201862 52020
rect 201730 51944 201782 51950
rect 201730 51886 201782 51892
rect 201820 51946 201876 51955
rect 201820 51881 201876 51890
rect 201638 51808 201690 51814
rect 201638 51750 201690 51756
rect 201776 51808 201828 51814
rect 201776 51750 201828 51756
rect 201926 51762 201954 52020
rect 202018 51882 202046 52020
rect 202006 51876 202058 51882
rect 202006 51818 202058 51824
rect 201684 51672 201736 51678
rect 201684 51614 201736 51620
rect 201512 51496 201586 51524
rect 201406 48376 201462 48385
rect 201406 48311 201462 48320
rect 201512 48142 201540 51496
rect 201592 51400 201644 51406
rect 201592 51342 201644 51348
rect 201604 50658 201632 51342
rect 201592 50652 201644 50658
rect 201592 50594 201644 50600
rect 201500 48136 201552 48142
rect 201500 48078 201552 48084
rect 201500 46708 201552 46714
rect 201500 46650 201552 46656
rect 201408 46640 201460 46646
rect 201408 46582 201460 46588
rect 201316 46096 201368 46102
rect 201316 46038 201368 46044
rect 201224 45892 201276 45898
rect 201224 45834 201276 45840
rect 201420 43382 201448 46582
rect 201512 46209 201540 46650
rect 201592 46436 201644 46442
rect 201592 46378 201644 46384
rect 201498 46200 201554 46209
rect 201498 46135 201554 46144
rect 201500 46096 201552 46102
rect 201500 46038 201552 46044
rect 201408 43376 201460 43382
rect 201408 43318 201460 43324
rect 200948 40724 201000 40730
rect 200948 40666 201000 40672
rect 200856 37120 200908 37126
rect 200856 37062 200908 37068
rect 200764 28348 200816 28354
rect 200764 28290 200816 28296
rect 200672 27124 200724 27130
rect 200672 27066 200724 27072
rect 200580 25628 200632 25634
rect 200580 25570 200632 25576
rect 200488 24336 200540 24342
rect 200488 24278 200540 24284
rect 200396 20392 200448 20398
rect 200396 20334 200448 20340
rect 200304 12300 200356 12306
rect 200304 12242 200356 12248
rect 200212 9240 200264 9246
rect 200212 9182 200264 9188
rect 198832 7812 198884 7818
rect 198832 7754 198884 7760
rect 198740 5024 198792 5030
rect 198740 4966 198792 4972
rect 201512 4962 201540 46038
rect 201604 6390 201632 46378
rect 201696 46170 201724 51614
rect 201788 46714 201816 51750
rect 201926 51734 202000 51762
rect 201868 51672 201920 51678
rect 201868 51614 201920 51620
rect 201776 46708 201828 46714
rect 201776 46650 201828 46656
rect 201880 46646 201908 51614
rect 201972 46753 202000 51734
rect 202110 51626 202138 52020
rect 202202 51950 202230 52020
rect 202190 51944 202242 51950
rect 202190 51886 202242 51892
rect 202294 51796 202322 52020
rect 202386 51921 202414 52020
rect 202372 51912 202428 51921
rect 202372 51847 202428 51856
rect 202294 51768 202368 51796
rect 202236 51672 202288 51678
rect 202110 51598 202184 51626
rect 202236 51614 202288 51620
rect 202052 51400 202104 51406
rect 202052 51342 202104 51348
rect 202064 50590 202092 51342
rect 202052 50584 202104 50590
rect 202052 50526 202104 50532
rect 202050 49736 202106 49745
rect 202050 49671 202106 49680
rect 202064 48346 202092 49671
rect 202052 48340 202104 48346
rect 202052 48282 202104 48288
rect 201958 46744 202014 46753
rect 201958 46679 202014 46688
rect 201868 46640 201920 46646
rect 201868 46582 201920 46588
rect 201866 46472 201922 46481
rect 201866 46407 201922 46416
rect 201880 46288 201908 46407
rect 201880 46260 202000 46288
rect 201866 46200 201922 46209
rect 201684 46164 201736 46170
rect 201866 46135 201922 46144
rect 201684 46106 201736 46112
rect 201684 46028 201736 46034
rect 201684 45970 201736 45976
rect 201696 7750 201724 45970
rect 201776 43376 201828 43382
rect 201776 43318 201828 43324
rect 201788 10470 201816 43318
rect 201880 23186 201908 46135
rect 201868 23180 201920 23186
rect 201868 23122 201920 23128
rect 201972 23118 202000 46260
rect 202052 46164 202104 46170
rect 202052 46106 202104 46112
rect 202064 29850 202092 46106
rect 202156 38282 202184 51598
rect 202248 46102 202276 51614
rect 202340 46442 202368 51768
rect 202478 51762 202506 52020
rect 202432 51734 202506 51762
rect 202328 46436 202380 46442
rect 202328 46378 202380 46384
rect 202236 46096 202288 46102
rect 202236 46038 202288 46044
rect 202432 46034 202460 51734
rect 202570 51660 202598 52020
rect 202662 51882 202690 52020
rect 202650 51876 202702 51882
rect 202650 51818 202702 51824
rect 202754 51762 202782 52020
rect 202524 51632 202598 51660
rect 202708 51734 202782 51762
rect 202524 48929 202552 51632
rect 202604 51536 202656 51542
rect 202604 51478 202656 51484
rect 202510 48920 202566 48929
rect 202510 48855 202566 48864
rect 202616 48657 202644 51478
rect 202602 48648 202658 48657
rect 202602 48583 202658 48592
rect 202512 48408 202564 48414
rect 202708 48385 202736 51734
rect 202846 51660 202874 52020
rect 202938 51882 202966 52020
rect 203030 51950 203058 52020
rect 203018 51944 203070 51950
rect 203018 51886 203070 51892
rect 202926 51876 202978 51882
rect 202926 51818 202978 51824
rect 203122 51762 203150 52020
rect 202800 51632 202874 51660
rect 202984 51734 203150 51762
rect 202800 48521 202828 51632
rect 202786 48512 202842 48521
rect 202786 48447 202842 48456
rect 202512 48350 202564 48356
rect 202694 48376 202750 48385
rect 202420 46028 202472 46034
rect 202420 45970 202472 45976
rect 202524 41414 202552 48350
rect 202694 48311 202750 48320
rect 202880 46096 202932 46102
rect 202880 46038 202932 46044
rect 202432 41386 202552 41414
rect 202144 38276 202196 38282
rect 202144 38218 202196 38224
rect 202052 29844 202104 29850
rect 202052 29786 202104 29792
rect 201960 23112 202012 23118
rect 201960 23054 202012 23060
rect 202432 15162 202460 41386
rect 202420 15156 202472 15162
rect 202420 15098 202472 15104
rect 201776 10464 201828 10470
rect 201776 10406 201828 10412
rect 202892 9178 202920 46038
rect 202984 16386 203012 51734
rect 203064 51672 203116 51678
rect 203214 51626 203242 52020
rect 203306 51762 203334 52020
rect 203398 51882 203426 52020
rect 203386 51876 203438 51882
rect 203386 51818 203438 51824
rect 203490 51762 203518 52020
rect 203582 51882 203610 52020
rect 203674 51882 203702 52020
rect 203766 51882 203794 52020
rect 203570 51876 203622 51882
rect 203570 51818 203622 51824
rect 203662 51876 203714 51882
rect 203662 51818 203714 51824
rect 203754 51876 203806 51882
rect 203754 51818 203806 51824
rect 203858 51762 203886 52020
rect 203306 51734 203380 51762
rect 203490 51734 203748 51762
rect 203064 51614 203116 51620
rect 203076 47530 203104 51614
rect 203168 51598 203242 51626
rect 203168 48414 203196 51598
rect 203248 51536 203300 51542
rect 203248 51478 203300 51484
rect 203156 48408 203208 48414
rect 203156 48350 203208 48356
rect 203064 47524 203116 47530
rect 203064 47466 203116 47472
rect 203064 46164 203116 46170
rect 203064 46106 203116 46112
rect 202972 16380 203024 16386
rect 202972 16322 203024 16328
rect 203076 16318 203104 46106
rect 203156 44464 203208 44470
rect 203156 44406 203208 44412
rect 203064 16312 203116 16318
rect 203064 16254 203116 16260
rect 203168 16250 203196 44406
rect 203260 20126 203288 51478
rect 203352 27062 203380 51734
rect 203432 51672 203484 51678
rect 203432 51614 203484 51620
rect 203524 51672 203576 51678
rect 203524 51614 203576 51620
rect 203444 46170 203472 51614
rect 203432 46164 203484 46170
rect 203432 46106 203484 46112
rect 203536 46102 203564 51614
rect 203616 51604 203668 51610
rect 203616 51546 203668 51552
rect 203524 46096 203576 46102
rect 203524 46038 203576 46044
rect 203628 44470 203656 51546
rect 203720 49298 203748 51734
rect 203812 51734 203886 51762
rect 203950 51762 203978 52020
rect 204042 51882 204070 52020
rect 204134 51921 204162 52020
rect 204120 51912 204176 51921
rect 204030 51876 204082 51882
rect 204120 51847 204176 51856
rect 204030 51818 204082 51824
rect 204226 51762 204254 52020
rect 203950 51734 204024 51762
rect 203708 49292 203760 49298
rect 203708 49234 203760 49240
rect 203812 48385 203840 51734
rect 203892 51672 203944 51678
rect 203892 51614 203944 51620
rect 203904 49706 203932 51614
rect 203892 49700 203944 49706
rect 203892 49642 203944 49648
rect 203996 48929 204024 51734
rect 204180 51734 204254 51762
rect 204318 51762 204346 52020
rect 204410 51950 204438 52020
rect 204398 51944 204450 51950
rect 204502 51921 204530 52020
rect 204594 51950 204622 52020
rect 204686 51950 204714 52020
rect 204778 51950 204806 52020
rect 204870 51950 204898 52020
rect 204962 51950 204990 52020
rect 205054 51950 205082 52020
rect 204582 51944 204634 51950
rect 204398 51886 204450 51892
rect 204488 51912 204544 51921
rect 204582 51886 204634 51892
rect 204674 51944 204726 51950
rect 204674 51886 204726 51892
rect 204766 51944 204818 51950
rect 204766 51886 204818 51892
rect 204858 51944 204910 51950
rect 204858 51886 204910 51892
rect 204950 51944 205002 51950
rect 204950 51886 205002 51892
rect 205042 51944 205094 51950
rect 205042 51886 205094 51892
rect 204488 51847 204544 51856
rect 204950 51808 205002 51814
rect 204318 51734 204392 51762
rect 204950 51750 205002 51756
rect 204076 51604 204128 51610
rect 204076 51546 204128 51552
rect 204088 49910 204116 51546
rect 204180 50153 204208 51734
rect 204260 51672 204312 51678
rect 204260 51614 204312 51620
rect 204272 50318 204300 51614
rect 204260 50312 204312 50318
rect 204260 50254 204312 50260
rect 204166 50144 204222 50153
rect 204166 50079 204222 50088
rect 204076 49904 204128 49910
rect 204076 49846 204128 49852
rect 203982 48920 204038 48929
rect 203982 48855 204038 48864
rect 203984 48680 204036 48686
rect 203984 48622 204036 48628
rect 203892 48476 203944 48482
rect 203892 48418 203944 48424
rect 203798 48376 203854 48385
rect 203708 48340 203760 48346
rect 203798 48311 203854 48320
rect 203708 48282 203760 48288
rect 203616 44464 203668 44470
rect 203616 44406 203668 44412
rect 203720 44282 203748 48282
rect 203628 44254 203748 44282
rect 203628 41414 203656 44254
rect 203708 44192 203760 44198
rect 203708 44134 203760 44140
rect 203536 41386 203656 41414
rect 203340 27056 203392 27062
rect 203340 26998 203392 27004
rect 203536 20262 203564 41386
rect 203720 39438 203748 44134
rect 203904 41414 203932 48418
rect 203996 44198 204024 48622
rect 204364 46782 204392 51734
rect 204628 51740 204680 51746
rect 204628 51682 204680 51688
rect 204720 51740 204772 51746
rect 204720 51682 204772 51688
rect 204444 51536 204496 51542
rect 204444 51478 204496 51484
rect 204456 49774 204484 51478
rect 204640 50658 204668 51682
rect 204628 50652 204680 50658
rect 204628 50594 204680 50600
rect 204732 50402 204760 51682
rect 204962 51660 204990 51750
rect 205146 51728 205174 52020
rect 205238 51955 205266 52020
rect 205224 51946 205280 51955
rect 205330 51950 205358 52020
rect 205224 51881 205280 51890
rect 205318 51944 205370 51950
rect 205422 51921 205450 52020
rect 205514 51950 205542 52020
rect 205606 51950 205634 52020
rect 205698 51950 205726 52020
rect 205790 51950 205818 52020
rect 205502 51944 205554 51950
rect 205318 51886 205370 51892
rect 205408 51912 205464 51921
rect 205502 51886 205554 51892
rect 205594 51944 205646 51950
rect 205594 51886 205646 51892
rect 205686 51944 205738 51950
rect 205686 51886 205738 51892
rect 205778 51944 205830 51950
rect 205778 51886 205830 51892
rect 205882 51882 205910 52020
rect 205408 51847 205464 51856
rect 205870 51876 205922 51882
rect 205870 51818 205922 51824
rect 205974 51814 206002 52020
rect 205272 51808 205324 51814
rect 205272 51750 205324 51756
rect 205456 51808 205508 51814
rect 205456 51750 205508 51756
rect 205732 51808 205784 51814
rect 205732 51750 205784 51756
rect 205962 51808 206014 51814
rect 205962 51750 206014 51756
rect 205146 51700 205220 51728
rect 204962 51632 205128 51660
rect 204640 50374 204760 50402
rect 204640 50164 204668 50374
rect 204996 50244 205048 50250
rect 204996 50186 205048 50192
rect 204812 50176 204864 50182
rect 204534 50144 204590 50153
rect 204640 50136 204760 50164
rect 204534 50079 204590 50088
rect 204444 49768 204496 49774
rect 204444 49710 204496 49716
rect 204444 48748 204496 48754
rect 204444 48690 204496 48696
rect 204352 46776 204404 46782
rect 204352 46718 204404 46724
rect 204456 46510 204484 48690
rect 204444 46504 204496 46510
rect 204444 46446 204496 46452
rect 204352 46436 204404 46442
rect 204352 46378 204404 46384
rect 204260 46096 204312 46102
rect 204260 46038 204312 46044
rect 203984 44192 204036 44198
rect 203984 44134 204036 44140
rect 203812 41386 203932 41414
rect 203708 39432 203760 39438
rect 203708 39374 203760 39380
rect 203524 20256 203576 20262
rect 203524 20198 203576 20204
rect 203248 20120 203300 20126
rect 203248 20062 203300 20068
rect 203524 19984 203576 19990
rect 203524 19926 203576 19932
rect 203156 16244 203208 16250
rect 203156 16186 203208 16192
rect 202880 9172 202932 9178
rect 202880 9114 202932 9120
rect 201684 7744 201736 7750
rect 201684 7686 201736 7692
rect 201592 6384 201644 6390
rect 201592 6326 201644 6332
rect 201500 4956 201552 4962
rect 201500 4898 201552 4904
rect 201500 4072 201552 4078
rect 201500 4014 201552 4020
rect 200304 3936 200356 3942
rect 200304 3878 200356 3884
rect 199108 3324 199160 3330
rect 199108 3266 199160 3272
rect 197912 3256 197964 3262
rect 197912 3198 197964 3204
rect 197924 480 197952 3198
rect 199120 480 199148 3266
rect 200316 480 200344 3878
rect 201512 480 201540 4014
rect 202696 3392 202748 3398
rect 202696 3334 202748 3340
rect 202708 480 202736 3334
rect 203536 3194 203564 19926
rect 203812 12374 203840 41386
rect 203984 15904 204036 15910
rect 203984 15846 204036 15852
rect 203800 12368 203852 12374
rect 203800 12310 203852 12316
rect 203996 3738 204024 15846
rect 204272 6322 204300 46038
rect 204364 16046 204392 46378
rect 204444 46164 204496 46170
rect 204444 46106 204496 46112
rect 204456 16114 204484 46106
rect 204548 16182 204576 50079
rect 204628 48408 204680 48414
rect 204628 48350 204680 48356
rect 204640 46986 204668 48350
rect 204628 46980 204680 46986
rect 204628 46922 204680 46928
rect 204628 46776 204680 46782
rect 204628 46718 204680 46724
rect 204640 20058 204668 46718
rect 204732 46170 204760 50136
rect 204812 50118 204864 50124
rect 204720 46164 204772 46170
rect 204720 46106 204772 46112
rect 204824 46102 204852 50118
rect 204902 49872 204958 49881
rect 204902 49807 204958 49816
rect 204812 46096 204864 46102
rect 204812 46038 204864 46044
rect 204720 46028 204772 46034
rect 204720 45970 204772 45976
rect 204732 21554 204760 45970
rect 204916 41414 204944 49807
rect 205008 46442 205036 50186
rect 205100 50182 205128 51632
rect 205192 50182 205220 51700
rect 205088 50176 205140 50182
rect 205088 50118 205140 50124
rect 205180 50176 205232 50182
rect 205180 50118 205232 50124
rect 205284 48314 205312 51750
rect 205364 51672 205416 51678
rect 205364 51614 205416 51620
rect 205376 50046 205404 51614
rect 205468 50153 205496 51750
rect 205640 51740 205692 51746
rect 205560 51700 205640 51728
rect 205454 50144 205510 50153
rect 205454 50079 205510 50088
rect 205364 50040 205416 50046
rect 205364 49982 205416 49988
rect 205100 48286 205312 48314
rect 205362 48376 205418 48385
rect 205362 48311 205418 48320
rect 204996 46436 205048 46442
rect 204996 46378 205048 46384
rect 205100 46034 205128 48286
rect 205376 48226 205404 48311
rect 205560 48226 205588 51700
rect 205640 51682 205692 51688
rect 205640 51604 205692 51610
rect 205640 51546 205692 51552
rect 205652 50590 205680 51546
rect 205640 50584 205692 50590
rect 205640 50526 205692 50532
rect 205640 50176 205692 50182
rect 205640 50118 205692 50124
rect 205376 48198 205588 48226
rect 205652 48074 205680 50118
rect 205744 48754 205772 51750
rect 205916 51604 205968 51610
rect 206066 51592 206094 52020
rect 206158 51955 206186 52020
rect 206144 51946 206200 51955
rect 206250 51950 206278 52020
rect 206342 51955 206370 52020
rect 206144 51881 206200 51890
rect 206238 51944 206290 51950
rect 206238 51886 206290 51892
rect 206328 51946 206384 51955
rect 206328 51881 206384 51890
rect 206434 51882 206462 52020
rect 206422 51876 206474 51882
rect 206422 51818 206474 51824
rect 206526 51728 206554 52020
rect 206618 51950 206646 52020
rect 206710 51950 206738 52020
rect 206606 51944 206658 51950
rect 206606 51886 206658 51892
rect 206698 51944 206750 51950
rect 206698 51886 206750 51892
rect 206802 51882 206830 52020
rect 206894 51955 206922 52020
rect 206880 51946 206936 51955
rect 206986 51950 207014 52020
rect 206790 51876 206842 51882
rect 206880 51881 206936 51890
rect 206974 51944 207026 51950
rect 207078 51921 207106 52020
rect 207170 51950 207198 52020
rect 207158 51944 207210 51950
rect 206974 51886 207026 51892
rect 207064 51912 207120 51921
rect 207158 51886 207210 51892
rect 207064 51847 207120 51856
rect 206790 51818 206842 51824
rect 207262 51814 207290 52020
rect 206606 51808 206658 51814
rect 206928 51808 206980 51814
rect 206606 51750 206658 51756
rect 206848 51756 206928 51762
rect 206848 51750 206980 51756
rect 207250 51808 207302 51814
rect 207354 51785 207382 52020
rect 207446 51882 207474 52020
rect 207434 51876 207486 51882
rect 207434 51818 207486 51824
rect 207250 51750 207302 51756
rect 207340 51776 207396 51785
rect 206480 51700 206554 51728
rect 205916 51546 205968 51552
rect 206020 51564 206094 51592
rect 206192 51604 206244 51610
rect 205928 50232 205956 51546
rect 205836 50204 205956 50232
rect 205732 48748 205784 48754
rect 205732 48690 205784 48696
rect 205640 48068 205692 48074
rect 205640 48010 205692 48016
rect 205836 47462 205864 50204
rect 205916 50040 205968 50046
rect 205916 49982 205968 49988
rect 205824 47456 205876 47462
rect 205824 47398 205876 47404
rect 205180 46980 205232 46986
rect 205180 46922 205232 46928
rect 205088 46028 205140 46034
rect 205088 45970 205140 45976
rect 204824 41386 204944 41414
rect 204824 23050 204852 41386
rect 204812 23044 204864 23050
rect 204812 22986 204864 22992
rect 204720 21548 204772 21554
rect 204720 21490 204772 21496
rect 205192 20194 205220 46922
rect 205272 46504 205324 46510
rect 205272 46446 205324 46452
rect 205284 32570 205312 46446
rect 205732 46164 205784 46170
rect 205732 46106 205784 46112
rect 205272 32564 205324 32570
rect 205272 32506 205324 32512
rect 205180 20188 205232 20194
rect 205180 20130 205232 20136
rect 204628 20052 204680 20058
rect 204628 19994 204680 20000
rect 204536 16176 204588 16182
rect 204536 16118 204588 16124
rect 204444 16108 204496 16114
rect 204444 16050 204496 16056
rect 204352 16040 204404 16046
rect 204352 15982 204404 15988
rect 205744 12102 205772 46106
rect 205824 46096 205876 46102
rect 205824 46038 205876 46044
rect 205732 12096 205784 12102
rect 205732 12038 205784 12044
rect 205836 12034 205864 46038
rect 205928 12238 205956 49982
rect 205916 12232 205968 12238
rect 205916 12174 205968 12180
rect 206020 12170 206048 51564
rect 206192 51546 206244 51552
rect 206376 51604 206428 51610
rect 206376 51546 206428 51552
rect 206100 50584 206152 50590
rect 206100 50526 206152 50532
rect 206112 50266 206140 50526
rect 206204 50368 206232 51546
rect 206284 51536 206336 51542
rect 206284 51478 206336 51484
rect 206296 50590 206324 51478
rect 206284 50584 206336 50590
rect 206284 50526 206336 50532
rect 206204 50340 206324 50368
rect 206112 50250 206232 50266
rect 206112 50244 206244 50250
rect 206112 50238 206192 50244
rect 206192 50186 206244 50192
rect 206100 50176 206152 50182
rect 206100 50118 206152 50124
rect 206112 14754 206140 50118
rect 206190 50008 206246 50017
rect 206190 49943 206246 49952
rect 206204 14822 206232 49943
rect 206296 48686 206324 50340
rect 206388 50182 206416 51546
rect 206376 50176 206428 50182
rect 206376 50118 206428 50124
rect 206284 48680 206336 48686
rect 206284 48622 206336 48628
rect 206480 48532 206508 51700
rect 206618 51626 206646 51750
rect 206744 51740 206796 51746
rect 206744 51682 206796 51688
rect 206848 51734 206968 51750
rect 206296 48504 206508 48532
rect 206572 51598 206646 51626
rect 206296 19990 206324 48504
rect 206466 48376 206522 48385
rect 206466 48311 206522 48320
rect 206480 46170 206508 48311
rect 206468 46164 206520 46170
rect 206468 46106 206520 46112
rect 206572 46102 206600 51598
rect 206652 49292 206704 49298
rect 206652 49234 206704 49240
rect 206560 46096 206612 46102
rect 206560 46038 206612 46044
rect 206284 19984 206336 19990
rect 206284 19926 206336 19932
rect 206664 18766 206692 49234
rect 206652 18760 206704 18766
rect 206652 18702 206704 18708
rect 206192 14816 206244 14822
rect 206192 14758 206244 14764
rect 206100 14748 206152 14754
rect 206100 14690 206152 14696
rect 206008 12164 206060 12170
rect 206008 12106 206060 12112
rect 205824 12028 205876 12034
rect 205824 11970 205876 11976
rect 206192 10328 206244 10334
rect 206192 10270 206244 10276
rect 204260 6316 204312 6322
rect 204260 6258 204312 6264
rect 205088 4004 205140 4010
rect 205088 3946 205140 3952
rect 203892 3732 203944 3738
rect 203892 3674 203944 3680
rect 203984 3732 204036 3738
rect 203984 3674 204036 3680
rect 203524 3188 203576 3194
rect 203524 3130 203576 3136
rect 203904 480 203932 3674
rect 205100 480 205128 3946
rect 206204 480 206232 10270
rect 206756 9110 206784 51682
rect 206848 50017 206876 51734
rect 207340 51711 207396 51720
rect 206928 51672 206980 51678
rect 207538 51660 207566 52020
rect 207630 51785 207658 52020
rect 207722 51882 207750 52020
rect 207710 51876 207762 51882
rect 207710 51818 207762 51824
rect 207814 51796 207842 52020
rect 207906 51950 207934 52020
rect 207894 51944 207946 51950
rect 207894 51886 207946 51892
rect 207616 51776 207672 51785
rect 207814 51768 207888 51796
rect 207616 51711 207672 51720
rect 207756 51672 207808 51678
rect 207538 51632 207612 51660
rect 206928 51614 206980 51620
rect 206940 50153 206968 51614
rect 207020 51604 207072 51610
rect 207020 51546 207072 51552
rect 207204 51604 207256 51610
rect 207204 51546 207256 51552
rect 206926 50144 206982 50153
rect 206926 50079 206982 50088
rect 206834 50008 206890 50017
rect 206834 49943 206890 49952
rect 207032 11966 207060 51546
rect 207112 50380 207164 50386
rect 207112 50322 207164 50328
rect 207124 49978 207152 50322
rect 207216 50046 207244 51546
rect 207388 51536 207440 51542
rect 207388 51478 207440 51484
rect 207480 51536 207532 51542
rect 207480 51478 207532 51484
rect 207296 50380 207348 50386
rect 207296 50322 207348 50328
rect 207204 50040 207256 50046
rect 207204 49982 207256 49988
rect 207112 49972 207164 49978
rect 207112 49914 207164 49920
rect 207112 46164 207164 46170
rect 207112 46106 207164 46112
rect 207124 14550 207152 46106
rect 207308 46050 207336 50322
rect 207400 50153 207428 51478
rect 207492 50386 207520 51478
rect 207480 50380 207532 50386
rect 207480 50322 207532 50328
rect 207480 50244 207532 50250
rect 207480 50186 207532 50192
rect 207386 50144 207442 50153
rect 207386 50079 207442 50088
rect 207388 50040 207440 50046
rect 207388 49982 207440 49988
rect 207216 46022 207336 46050
rect 207216 14686 207244 46022
rect 207296 45960 207348 45966
rect 207296 45902 207348 45908
rect 207204 14680 207256 14686
rect 207204 14622 207256 14628
rect 207308 14618 207336 45902
rect 207400 17814 207428 49982
rect 207388 17808 207440 17814
rect 207388 17750 207440 17756
rect 207492 17678 207520 50186
rect 207584 17746 207612 51632
rect 207756 51614 207808 51620
rect 207664 51604 207716 51610
rect 207664 51546 207716 51552
rect 207676 38146 207704 51546
rect 207768 45966 207796 51614
rect 207860 50250 207888 51768
rect 207998 51762 208026 52020
rect 208090 51785 208118 52020
rect 208182 51921 208210 52020
rect 208274 51950 208302 52020
rect 208366 51950 208394 52020
rect 208458 51950 208486 52020
rect 208262 51944 208314 51950
rect 208168 51912 208224 51921
rect 208262 51886 208314 51892
rect 208354 51944 208406 51950
rect 208354 51886 208406 51892
rect 208446 51944 208498 51950
rect 208446 51886 208498 51892
rect 208550 51882 208578 52020
rect 208734 51932 208762 52020
rect 208688 51904 208762 51932
rect 208168 51847 208224 51856
rect 208538 51876 208590 51882
rect 208538 51818 208590 51824
rect 207952 51734 208026 51762
rect 208076 51776 208132 51785
rect 207848 50244 207900 50250
rect 207848 50186 207900 50192
rect 207848 49768 207900 49774
rect 207848 49710 207900 49716
rect 207756 45960 207808 45966
rect 207756 45902 207808 45908
rect 207664 38140 207716 38146
rect 207664 38082 207716 38088
rect 207572 17740 207624 17746
rect 207572 17682 207624 17688
rect 207480 17672 207532 17678
rect 207480 17614 207532 17620
rect 207296 14612 207348 14618
rect 207296 14554 207348 14560
rect 207112 14544 207164 14550
rect 207112 14486 207164 14492
rect 207020 11960 207072 11966
rect 207020 11902 207072 11908
rect 206744 9104 206796 9110
rect 206744 9046 206796 9052
rect 207018 4856 207074 4865
rect 207018 4791 207074 4800
rect 207032 2854 207060 4791
rect 207860 3806 207888 49710
rect 207952 46170 207980 51734
rect 208688 51746 208716 51904
rect 208826 51864 208854 52020
rect 208918 51882 208946 52020
rect 209010 51921 209038 52020
rect 209102 51950 209130 52020
rect 209090 51944 209142 51950
rect 208996 51912 209052 51921
rect 208780 51836 208854 51864
rect 208906 51876 208958 51882
rect 208076 51711 208132 51720
rect 208216 51740 208268 51746
rect 208216 51682 208268 51688
rect 208308 51740 208360 51746
rect 208308 51682 208360 51688
rect 208676 51740 208728 51746
rect 208676 51682 208728 51688
rect 208032 50584 208084 50590
rect 208032 50526 208084 50532
rect 208044 50368 208072 50526
rect 208044 50340 208164 50368
rect 208032 50244 208084 50250
rect 208032 50186 208084 50192
rect 208044 49881 208072 50186
rect 208030 49872 208086 49881
rect 208030 49807 208086 49816
rect 208032 49700 208084 49706
rect 208032 49642 208084 49648
rect 207940 46164 207992 46170
rect 207940 46106 207992 46112
rect 208044 41414 208072 49642
rect 208136 48482 208164 50340
rect 208228 49230 208256 51682
rect 208320 50250 208348 51682
rect 208400 51672 208452 51678
rect 208400 51614 208452 51620
rect 208308 50244 208360 50250
rect 208308 50186 208360 50192
rect 208412 50182 208440 51614
rect 208676 51604 208728 51610
rect 208676 51546 208728 51552
rect 208492 50244 208544 50250
rect 208492 50186 208544 50192
rect 208400 50176 208452 50182
rect 208306 50144 208362 50153
rect 208400 50118 208452 50124
rect 208306 50079 208362 50088
rect 208320 49298 208348 50079
rect 208400 50040 208452 50046
rect 208400 49982 208452 49988
rect 208308 49292 208360 49298
rect 208308 49234 208360 49240
rect 208216 49224 208268 49230
rect 208216 49166 208268 49172
rect 208306 48648 208362 48657
rect 208306 48583 208362 48592
rect 208320 48550 208348 48583
rect 208308 48544 208360 48550
rect 208308 48486 208360 48492
rect 208124 48476 208176 48482
rect 208124 48418 208176 48424
rect 207952 41386 208072 41414
rect 207952 31210 207980 41386
rect 207940 31204 207992 31210
rect 207940 31146 207992 31152
rect 208412 4894 208440 49982
rect 208504 8974 208532 50186
rect 208584 50176 208636 50182
rect 208584 50118 208636 50124
rect 208596 9042 208624 50118
rect 208688 10402 208716 51546
rect 208780 44062 208808 51836
rect 209090 51886 209142 51892
rect 208996 51847 209052 51856
rect 208906 51818 208958 51824
rect 208950 51776 209006 51785
rect 208872 51734 208950 51762
rect 208768 44056 208820 44062
rect 208768 43998 208820 44004
rect 208768 43920 208820 43926
rect 208768 43862 208820 43868
rect 208780 11898 208808 43862
rect 208872 15978 208900 51734
rect 209194 51762 209222 52020
rect 209286 51921 209314 52020
rect 209272 51912 209328 51921
rect 209272 51847 209328 51856
rect 209378 51762 209406 52020
rect 209470 51950 209498 52020
rect 209458 51944 209510 51950
rect 209458 51886 209510 51892
rect 209562 51785 209590 52020
rect 209654 51955 209682 52020
rect 209640 51946 209696 51955
rect 209640 51881 209696 51890
rect 208950 51711 209006 51720
rect 209148 51734 209222 51762
rect 209332 51734 209406 51762
rect 209548 51776 209604 51785
rect 208952 51672 209004 51678
rect 208952 51614 209004 51620
rect 209044 51672 209096 51678
rect 209044 51614 209096 51620
rect 208964 24274 208992 51614
rect 209056 35358 209084 51614
rect 209148 50046 209176 51734
rect 209332 51592 209360 51734
rect 209548 51711 209604 51720
rect 209504 51672 209556 51678
rect 209240 51564 209360 51592
rect 209424 51632 209504 51660
rect 209136 50040 209188 50046
rect 209136 49982 209188 49988
rect 209136 48952 209188 48958
rect 209134 48920 209136 48929
rect 209188 48920 209190 48929
rect 209134 48855 209190 48864
rect 209240 44146 209268 51564
rect 209424 50250 209452 51632
rect 209746 51660 209774 52020
rect 209838 51728 209866 52020
rect 209930 51882 209958 52020
rect 210022 51950 210050 52020
rect 210010 51944 210062 51950
rect 210010 51886 210062 51892
rect 209918 51876 209970 51882
rect 209918 51818 209970 51824
rect 210114 51728 210142 52020
rect 210206 51796 210234 52020
rect 210298 51921 210326 52020
rect 210284 51912 210340 51921
rect 210284 51847 210340 51856
rect 210206 51768 210280 51796
rect 209838 51700 210004 51728
rect 210114 51700 210188 51728
rect 209746 51632 209820 51660
rect 209504 51614 209556 51620
rect 209596 51604 209648 51610
rect 209596 51546 209648 51552
rect 209412 50244 209464 50250
rect 209412 50186 209464 50192
rect 209608 50153 209636 51546
rect 209688 51536 209740 51542
rect 209688 51478 209740 51484
rect 209318 50144 209374 50153
rect 209318 50079 209374 50088
rect 209594 50144 209650 50153
rect 209594 50079 209650 50088
rect 209148 44118 209268 44146
rect 209044 35352 209096 35358
rect 209044 35294 209096 35300
rect 209148 35290 209176 44118
rect 209228 44056 209280 44062
rect 209228 43998 209280 44004
rect 209240 38214 209268 43998
rect 209332 43926 209360 50079
rect 209594 49736 209650 49745
rect 209594 49671 209650 49680
rect 209608 49094 209636 49671
rect 209700 49502 209728 51478
rect 209792 50017 209820 51632
rect 209778 50008 209834 50017
rect 209778 49943 209834 49952
rect 209870 49736 209926 49745
rect 209870 49671 209926 49680
rect 209688 49496 209740 49502
rect 209688 49438 209740 49444
rect 209596 49088 209648 49094
rect 209596 49030 209648 49036
rect 209778 49056 209834 49065
rect 209778 48991 209834 49000
rect 209792 48958 209820 48991
rect 209780 48952 209832 48958
rect 209780 48894 209832 48900
rect 209778 48784 209834 48793
rect 209778 48719 209834 48728
rect 209320 43920 209372 43926
rect 209320 43862 209372 43868
rect 209228 38208 209280 38214
rect 209228 38150 209280 38156
rect 209136 35284 209188 35290
rect 209136 35226 209188 35232
rect 208952 24268 209004 24274
rect 208952 24210 209004 24216
rect 208860 15972 208912 15978
rect 208860 15914 208912 15920
rect 208768 11892 208820 11898
rect 208768 11834 208820 11840
rect 208676 10396 208728 10402
rect 208676 10338 208728 10344
rect 208584 9036 208636 9042
rect 208584 8978 208636 8984
rect 208492 8968 208544 8974
rect 208492 8910 208544 8916
rect 209792 6254 209820 48719
rect 209884 7682 209912 49671
rect 209976 13190 210004 51700
rect 210056 51604 210108 51610
rect 210056 51546 210108 51552
rect 210068 48929 210096 51546
rect 210054 48920 210110 48929
rect 210054 48855 210110 48864
rect 210056 48816 210108 48822
rect 210056 48758 210108 48764
rect 210160 48770 210188 51700
rect 210252 48958 210280 51768
rect 210390 51660 210418 52020
rect 210482 51762 210510 52020
rect 210574 51921 210602 52020
rect 210666 51950 210694 52020
rect 210654 51944 210706 51950
rect 210560 51912 210616 51921
rect 210654 51886 210706 51892
rect 210560 51847 210616 51856
rect 210608 51808 210660 51814
rect 210482 51734 210556 51762
rect 210608 51750 210660 51756
rect 210758 51762 210786 52020
rect 210850 51882 210878 52020
rect 210942 51921 210970 52020
rect 210928 51912 210984 51921
rect 210838 51876 210890 51882
rect 210928 51847 210984 51856
rect 210838 51818 210890 51824
rect 210390 51632 210464 51660
rect 210332 51536 210384 51542
rect 210332 51478 210384 51484
rect 210344 50318 210372 51478
rect 210332 50312 210384 50318
rect 210332 50254 210384 50260
rect 210240 48952 210292 48958
rect 210240 48894 210292 48900
rect 210436 48822 210464 51632
rect 210424 48816 210476 48822
rect 210330 48784 210386 48793
rect 210068 15910 210096 48758
rect 210160 48742 210280 48770
rect 210148 48544 210200 48550
rect 210148 48486 210200 48492
rect 210160 17882 210188 48486
rect 210252 22982 210280 48742
rect 210424 48758 210476 48764
rect 210330 48719 210386 48728
rect 210240 22976 210292 22982
rect 210240 22918 210292 22924
rect 210344 22914 210372 48719
rect 210424 46164 210476 46170
rect 210424 46106 210476 46112
rect 210436 32502 210464 46106
rect 210528 38010 210556 51734
rect 210620 50386 210648 51750
rect 210758 51734 210924 51762
rect 210792 51672 210844 51678
rect 210792 51614 210844 51620
rect 210608 50380 210660 50386
rect 210608 50322 210660 50328
rect 210700 50380 210752 50386
rect 210700 50322 210752 50328
rect 210608 48952 210660 48958
rect 210608 48894 210660 48900
rect 210620 38078 210648 48894
rect 210712 46170 210740 50322
rect 210804 48793 210832 51614
rect 210896 50386 210924 51734
rect 211034 51660 211062 52020
rect 211126 51955 211154 52020
rect 211112 51946 211168 51955
rect 211112 51881 211168 51890
rect 211218 51728 211246 52020
rect 211172 51700 211246 51728
rect 211310 51728 211338 52020
rect 211402 51950 211430 52020
rect 211390 51944 211442 51950
rect 211390 51886 211442 51892
rect 211494 51814 211522 52020
rect 211482 51808 211534 51814
rect 211482 51750 211534 51756
rect 211310 51700 211384 51728
rect 211034 51632 211108 51660
rect 210976 51536 211028 51542
rect 210976 51478 211028 51484
rect 210884 50380 210936 50386
rect 210884 50322 210936 50328
rect 210884 48884 210936 48890
rect 210884 48826 210936 48832
rect 210790 48784 210846 48793
rect 210790 48719 210846 48728
rect 210896 48414 210924 48826
rect 210988 48550 211016 51478
rect 211080 50153 211108 51632
rect 211066 50144 211122 50153
rect 211066 50079 211122 50088
rect 210976 48544 211028 48550
rect 210976 48486 211028 48492
rect 210884 48408 210936 48414
rect 210884 48350 210936 48356
rect 211068 46572 211120 46578
rect 211068 46514 211120 46520
rect 210700 46164 210752 46170
rect 210700 46106 210752 46112
rect 211080 43382 211108 46514
rect 211172 46442 211200 51700
rect 211252 51604 211304 51610
rect 211252 51546 211304 51552
rect 211264 49910 211292 51546
rect 211356 50153 211384 51700
rect 211586 51660 211614 52020
rect 211678 51785 211706 52020
rect 211770 51882 211798 52020
rect 211758 51876 211810 51882
rect 211758 51818 211810 51824
rect 211664 51776 211720 51785
rect 211664 51711 211720 51720
rect 211540 51632 211614 51660
rect 211712 51672 211764 51678
rect 211436 51604 211488 51610
rect 211436 51546 211488 51552
rect 211342 50144 211398 50153
rect 211342 50079 211398 50088
rect 211252 49904 211304 49910
rect 211252 49846 211304 49852
rect 211344 46504 211396 46510
rect 211344 46446 211396 46452
rect 211160 46436 211212 46442
rect 211160 46378 211212 46384
rect 211356 45914 211384 46446
rect 211172 45886 211384 45914
rect 211068 43376 211120 43382
rect 211068 43318 211120 43324
rect 210608 38072 210660 38078
rect 210608 38014 210660 38020
rect 210516 38004 210568 38010
rect 210516 37946 210568 37952
rect 210424 32496 210476 32502
rect 210424 32438 210476 32444
rect 210332 22908 210384 22914
rect 210332 22850 210384 22856
rect 210148 17876 210200 17882
rect 210148 17818 210200 17824
rect 210422 17232 210478 17241
rect 210422 17167 210478 17176
rect 210056 15904 210108 15910
rect 210056 15846 210108 15852
rect 209964 13184 210016 13190
rect 209964 13126 210016 13132
rect 209872 7676 209924 7682
rect 209872 7618 209924 7624
rect 209780 6248 209832 6254
rect 209780 6190 209832 6196
rect 208400 4888 208452 4894
rect 208400 4830 208452 4836
rect 207388 3800 207440 3806
rect 207388 3742 207440 3748
rect 207848 3800 207900 3806
rect 207848 3742 207900 3748
rect 207020 2848 207072 2854
rect 207020 2790 207072 2796
rect 207400 480 207428 3742
rect 210436 3398 210464 17167
rect 211172 11762 211200 45886
rect 211344 45824 211396 45830
rect 211250 45792 211306 45801
rect 211344 45766 211396 45772
rect 211250 45727 211306 45736
rect 211264 11830 211292 45727
rect 211356 17474 211384 45766
rect 211448 17610 211476 51546
rect 211540 48822 211568 51632
rect 211862 51660 211890 52020
rect 211954 51728 211982 52020
rect 212046 51882 212074 52020
rect 212034 51876 212086 51882
rect 212034 51818 212086 51824
rect 212138 51728 212166 52020
rect 212230 51785 212258 52020
rect 212322 51955 212350 52020
rect 212308 51946 212364 51955
rect 212308 51881 212364 51890
rect 212414 51796 212442 52020
rect 212506 51921 212534 52020
rect 212492 51912 212548 51921
rect 212598 51882 212626 52020
rect 212492 51847 212548 51856
rect 212586 51876 212638 51882
rect 212586 51818 212638 51824
rect 211954 51700 212028 51728
rect 211862 51632 211936 51660
rect 211712 51614 211764 51620
rect 211620 51536 211672 51542
rect 211620 51478 211672 51484
rect 211528 48816 211580 48822
rect 211528 48758 211580 48764
rect 211528 43376 211580 43382
rect 211528 43318 211580 43324
rect 211436 17604 211488 17610
rect 211436 17546 211488 17552
rect 211540 17542 211568 43318
rect 211632 21486 211660 51478
rect 211724 46578 211752 51614
rect 211804 50380 211856 50386
rect 211804 50322 211856 50328
rect 211712 46572 211764 46578
rect 211712 46514 211764 46520
rect 211816 46510 211844 50322
rect 211804 46504 211856 46510
rect 211804 46446 211856 46452
rect 211712 46436 211764 46442
rect 211712 46378 211764 46384
rect 211724 22846 211752 46378
rect 211804 46164 211856 46170
rect 211804 46106 211856 46112
rect 211816 31074 211844 46106
rect 211908 36990 211936 51632
rect 212000 50386 212028 51700
rect 212092 51700 212166 51728
rect 212216 51776 212272 51785
rect 212216 51711 212272 51720
rect 212368 51768 212442 51796
rect 211988 50380 212040 50386
rect 211988 50322 212040 50328
rect 211988 50244 212040 50250
rect 211988 50186 212040 50192
rect 212000 49978 212028 50186
rect 211988 49972 212040 49978
rect 211988 49914 212040 49920
rect 211988 49360 212040 49366
rect 211988 49302 212040 49308
rect 212000 49026 212028 49302
rect 211988 49020 212040 49026
rect 211988 48962 212040 48968
rect 211988 48816 212040 48822
rect 211988 48758 212040 48764
rect 212000 37058 212028 48758
rect 212092 46170 212120 51700
rect 212172 51604 212224 51610
rect 212172 51546 212224 51552
rect 212080 46164 212132 46170
rect 212080 46106 212132 46112
rect 212184 45830 212212 51546
rect 212368 50674 212396 51768
rect 212540 51740 212592 51746
rect 212690 51728 212718 52020
rect 212782 51950 212810 52020
rect 212874 51950 212902 52020
rect 212966 51950 212994 52020
rect 212770 51944 212822 51950
rect 212770 51886 212822 51892
rect 212862 51944 212914 51950
rect 212862 51886 212914 51892
rect 212954 51944 213006 51950
rect 212954 51886 213006 51892
rect 213058 51882 213086 52020
rect 213046 51876 213098 51882
rect 213046 51818 213098 51824
rect 212816 51808 212868 51814
rect 212816 51750 212868 51756
rect 212540 51682 212592 51688
rect 212644 51700 212718 51728
rect 212448 51536 212500 51542
rect 212448 51478 212500 51484
rect 212276 50646 212396 50674
rect 212276 48793 212304 50646
rect 212262 48784 212318 48793
rect 212262 48719 212318 48728
rect 212460 46170 212488 51478
rect 212552 49774 212580 51682
rect 212644 49842 212672 51700
rect 212724 51604 212776 51610
rect 212724 51546 212776 51552
rect 212736 50046 212764 51546
rect 212724 50040 212776 50046
rect 212724 49982 212776 49988
rect 212632 49836 212684 49842
rect 212632 49778 212684 49784
rect 212540 49768 212592 49774
rect 212540 49710 212592 49716
rect 212724 49768 212776 49774
rect 212724 49710 212776 49716
rect 212540 48544 212592 48550
rect 212540 48486 212592 48492
rect 212448 46164 212500 46170
rect 212448 46106 212500 46112
rect 212172 45824 212224 45830
rect 212172 45766 212224 45772
rect 211988 37052 212040 37058
rect 211988 36994 212040 37000
rect 211896 36984 211948 36990
rect 211896 36926 211948 36932
rect 211804 31068 211856 31074
rect 211804 31010 211856 31016
rect 211712 22840 211764 22846
rect 211712 22782 211764 22788
rect 211620 21480 211672 21486
rect 211620 21422 211672 21428
rect 211802 17776 211858 17785
rect 211802 17711 211858 17720
rect 211528 17536 211580 17542
rect 211528 17478 211580 17484
rect 211344 17468 211396 17474
rect 211344 17410 211396 17416
rect 211252 11824 211304 11830
rect 211252 11766 211304 11772
rect 211160 11756 211212 11762
rect 211160 11698 211212 11704
rect 210976 3868 211028 3874
rect 210976 3810 211028 3816
rect 210424 3392 210476 3398
rect 210424 3334 210476 3340
rect 208584 3188 208636 3194
rect 208584 3130 208636 3136
rect 208596 480 208624 3130
rect 209780 2848 209832 2854
rect 209780 2790 209832 2796
rect 209792 480 209820 2790
rect 210988 480 211016 3810
rect 211816 3534 211844 17711
rect 212552 14482 212580 48486
rect 212632 46436 212684 46442
rect 212632 46378 212684 46384
rect 212644 17338 212672 46378
rect 212736 17406 212764 49710
rect 212828 46442 212856 51750
rect 212908 51740 212960 51746
rect 213150 51728 213178 52020
rect 213242 51950 213270 52020
rect 213230 51944 213282 51950
rect 213334 51921 213362 52020
rect 213426 51950 213454 52020
rect 213414 51944 213466 51950
rect 213230 51886 213282 51892
rect 213320 51912 213376 51921
rect 213414 51886 213466 51892
rect 213518 51882 213546 52020
rect 213320 51847 213376 51856
rect 213506 51876 213558 51882
rect 213506 51818 213558 51824
rect 213366 51776 213422 51785
rect 213276 51740 213328 51746
rect 213150 51700 213224 51728
rect 212908 51682 212960 51688
rect 212920 49910 212948 51682
rect 213000 51604 213052 51610
rect 213000 51546 213052 51552
rect 212908 49904 212960 49910
rect 212908 49846 212960 49852
rect 212908 49768 212960 49774
rect 212908 49710 212960 49716
rect 212920 49434 212948 49710
rect 212908 49428 212960 49434
rect 212908 49370 212960 49376
rect 212816 46436 212868 46442
rect 212816 46378 212868 46384
rect 212816 46164 212868 46170
rect 212816 46106 212868 46112
rect 212724 17400 212776 17406
rect 212724 17342 212776 17348
rect 212632 17332 212684 17338
rect 212632 17274 212684 17280
rect 212828 17270 212856 46106
rect 213012 46050 213040 51546
rect 213092 50040 213144 50046
rect 213092 49982 213144 49988
rect 212920 46022 213040 46050
rect 212920 21418 212948 46022
rect 213000 43036 213052 43042
rect 213000 42978 213052 42984
rect 213012 25566 213040 42978
rect 213104 29782 213132 49982
rect 213196 48550 213224 51700
rect 213610 51728 213638 52020
rect 213702 51950 213730 52020
rect 213794 51950 213822 52020
rect 213690 51944 213742 51950
rect 213690 51886 213742 51892
rect 213782 51944 213834 51950
rect 213886 51921 213914 52020
rect 213978 51950 214006 52020
rect 213966 51944 214018 51950
rect 213782 51886 213834 51892
rect 213872 51912 213928 51921
rect 213966 51886 214018 51892
rect 214070 51882 214098 52020
rect 214162 51882 214190 52020
rect 213872 51847 213928 51856
rect 214058 51876 214110 51882
rect 214058 51818 214110 51824
rect 214150 51876 214202 51882
rect 214150 51818 214202 51824
rect 213690 51808 213742 51814
rect 213366 51711 213422 51720
rect 213276 51682 213328 51688
rect 213184 48544 213236 48550
rect 213184 48486 213236 48492
rect 213184 48340 213236 48346
rect 213184 48282 213236 48288
rect 213196 36854 213224 48282
rect 213288 36922 213316 51682
rect 213380 50130 213408 51711
rect 213472 51700 213638 51728
rect 213688 51776 213690 51785
rect 213742 51776 213744 51785
rect 213688 51711 213744 51720
rect 213826 51776 213882 51785
rect 213826 51711 213882 51720
rect 213920 51740 213972 51746
rect 213472 50454 213500 51700
rect 213552 51604 213604 51610
rect 213552 51546 213604 51552
rect 213644 51604 213696 51610
rect 213644 51546 213696 51552
rect 213460 50448 213512 50454
rect 213460 50390 213512 50396
rect 213380 50102 213500 50130
rect 213368 49904 213420 49910
rect 213368 49846 213420 49852
rect 213380 37942 213408 49846
rect 213472 45554 213500 50102
rect 213564 48346 213592 51546
rect 213656 50017 213684 51546
rect 213642 50008 213698 50017
rect 213642 49943 213698 49952
rect 213840 48929 213868 51711
rect 213920 51682 213972 51688
rect 214012 51740 214064 51746
rect 214012 51682 214064 51688
rect 213826 48920 213882 48929
rect 213826 48855 213882 48864
rect 213552 48340 213604 48346
rect 213552 48282 213604 48288
rect 213472 45526 213868 45554
rect 213840 43042 213868 45526
rect 213828 43036 213880 43042
rect 213828 42978 213880 42984
rect 213368 37936 213420 37942
rect 213368 37878 213420 37884
rect 213276 36916 213328 36922
rect 213276 36858 213328 36864
rect 213184 36848 213236 36854
rect 213184 36790 213236 36796
rect 213184 32428 213236 32434
rect 213184 32370 213236 32376
rect 213092 29776 213144 29782
rect 213092 29718 213144 29724
rect 213000 25560 213052 25566
rect 213000 25502 213052 25508
rect 212908 21412 212960 21418
rect 212908 21354 212960 21360
rect 212816 17264 212868 17270
rect 212816 17206 212868 17212
rect 212540 14476 212592 14482
rect 212540 14418 212592 14424
rect 213196 3942 213224 32370
rect 213932 6186 213960 51682
rect 214024 48958 214052 51682
rect 214104 51672 214156 51678
rect 214104 51614 214156 51620
rect 214012 48952 214064 48958
rect 214012 48894 214064 48900
rect 214116 48906 214144 51614
rect 214254 51592 214282 52020
rect 214346 51660 214374 52020
rect 214530 51762 214558 52020
rect 214484 51734 214558 51762
rect 214346 51632 214420 51660
rect 214254 51564 214328 51592
rect 214196 50448 214248 50454
rect 214196 50390 214248 50396
rect 214208 49745 214236 50390
rect 214194 49736 214250 49745
rect 214194 49671 214250 49680
rect 214116 48878 214236 48906
rect 214104 48816 214156 48822
rect 214104 48758 214156 48764
rect 214012 48748 214064 48754
rect 214012 48690 214064 48696
rect 214024 22778 214052 48690
rect 214116 24206 214144 48758
rect 214208 48550 214236 48878
rect 214300 48822 214328 51564
rect 214392 48822 214420 51632
rect 214288 48816 214340 48822
rect 214288 48758 214340 48764
rect 214380 48816 214432 48822
rect 214380 48758 214432 48764
rect 214484 48668 214512 51734
rect 214622 51524 214650 52020
rect 214714 51785 214742 52020
rect 214806 51955 214834 52020
rect 214792 51946 214848 51955
rect 214898 51950 214926 52020
rect 214792 51881 214848 51890
rect 214886 51944 214938 51950
rect 214886 51886 214938 51892
rect 214990 51796 215018 52020
rect 215082 51950 215110 52020
rect 215174 51950 215202 52020
rect 215266 51950 215294 52020
rect 215070 51944 215122 51950
rect 215070 51886 215122 51892
rect 215162 51944 215214 51950
rect 215162 51886 215214 51892
rect 215254 51944 215306 51950
rect 215254 51886 215306 51892
rect 215116 51808 215168 51814
rect 214700 51776 214756 51785
rect 214990 51768 215064 51796
rect 214700 51711 214756 51720
rect 214840 51740 214892 51746
rect 214840 51682 214892 51688
rect 214852 51626 214880 51682
rect 214576 51496 214650 51524
rect 214760 51598 214880 51626
rect 214932 51604 214984 51610
rect 214576 48770 214604 51496
rect 214576 48742 214696 48770
rect 214760 48754 214788 51598
rect 214932 51546 214984 51552
rect 214944 50674 214972 51546
rect 214852 50646 214972 50674
rect 214300 48640 214512 48668
rect 214196 48544 214248 48550
rect 214196 48486 214248 48492
rect 214194 48376 214250 48385
rect 214194 48311 214250 48320
rect 214104 24200 214156 24206
rect 214104 24142 214156 24148
rect 214208 24138 214236 48311
rect 214300 26994 214328 48640
rect 214472 48544 214524 48550
rect 214472 48486 214524 48492
rect 214380 48340 214432 48346
rect 214380 48282 214432 48288
rect 214392 28286 214420 48282
rect 214484 31142 214512 48486
rect 214562 47968 214618 47977
rect 214562 47903 214618 47912
rect 214576 33794 214604 47903
rect 214668 35222 214696 48742
rect 214748 48748 214800 48754
rect 214748 48690 214800 48696
rect 214852 48385 214880 50646
rect 214932 50584 214984 50590
rect 214932 50526 214984 50532
rect 214944 50318 214972 50526
rect 214932 50312 214984 50318
rect 214932 50254 214984 50260
rect 215036 48929 215064 51768
rect 215116 51750 215168 51756
rect 215208 51808 215260 51814
rect 215208 51750 215260 51756
rect 215022 48920 215078 48929
rect 215022 48855 215078 48864
rect 214932 48816 214984 48822
rect 214932 48758 214984 48764
rect 214838 48376 214894 48385
rect 214838 48311 214894 48320
rect 214944 41414 214972 48758
rect 215128 47977 215156 51750
rect 215220 48793 215248 51750
rect 215358 51626 215386 52020
rect 215450 51950 215478 52020
rect 215542 51955 215570 52020
rect 215438 51944 215490 51950
rect 215438 51886 215490 51892
rect 215528 51946 215584 51955
rect 215528 51881 215584 51890
rect 215634 51660 215662 52020
rect 215726 51950 215754 52020
rect 215818 51950 215846 52020
rect 215714 51944 215766 51950
rect 215714 51886 215766 51892
rect 215806 51944 215858 51950
rect 215806 51886 215858 51892
rect 215944 51944 215996 51950
rect 215944 51886 215996 51892
rect 215760 51808 215812 51814
rect 215760 51750 215812 51756
rect 215852 51808 215904 51814
rect 215852 51750 215904 51756
rect 215588 51632 215662 51660
rect 215358 51598 215432 51626
rect 215300 48884 215352 48890
rect 215300 48826 215352 48832
rect 215206 48784 215262 48793
rect 215206 48719 215262 48728
rect 215114 47968 215170 47977
rect 215114 47903 215170 47912
rect 214760 41386 214972 41414
rect 214760 36718 214788 41386
rect 214748 36712 214800 36718
rect 214748 36654 214800 36660
rect 214656 35216 214708 35222
rect 214656 35158 214708 35164
rect 214564 33788 214616 33794
rect 214564 33730 214616 33736
rect 214472 31136 214524 31142
rect 214472 31078 214524 31084
rect 214380 28280 214432 28286
rect 214380 28222 214432 28228
rect 214288 26988 214340 26994
rect 214288 26930 214340 26936
rect 214196 24132 214248 24138
rect 214196 24074 214248 24080
rect 214012 22772 214064 22778
rect 214012 22714 214064 22720
rect 213920 6180 213972 6186
rect 213920 6122 213972 6128
rect 215312 4826 215340 48826
rect 215404 7614 215432 51598
rect 215588 48906 215616 51632
rect 215496 48878 215616 48906
rect 215772 48890 215800 51750
rect 215760 48884 215812 48890
rect 215496 10334 215524 48878
rect 215760 48826 215812 48832
rect 215576 48816 215628 48822
rect 215576 48758 215628 48764
rect 215758 48784 215814 48793
rect 215588 13122 215616 48758
rect 215758 48719 215814 48728
rect 215668 48680 215720 48686
rect 215668 48622 215720 48628
rect 215680 26926 215708 48622
rect 215772 29714 215800 48719
rect 215864 32434 215892 51750
rect 215956 48686 215984 51886
rect 216048 48822 216076 52142
rect 216128 52148 216180 52154
rect 216128 52090 216180 52096
rect 216140 51678 216168 52090
rect 216128 51672 216180 51678
rect 216128 51614 216180 51620
rect 216232 51474 216260 52294
rect 216312 52216 216364 52222
rect 216312 52158 216364 52164
rect 216220 51468 216272 51474
rect 216220 51410 216272 51416
rect 216128 48952 216180 48958
rect 216128 48894 216180 48900
rect 216036 48816 216088 48822
rect 216036 48758 216088 48764
rect 215944 48680 215996 48686
rect 215944 48622 215996 48628
rect 215944 48476 215996 48482
rect 215944 48418 215996 48424
rect 215852 32428 215904 32434
rect 215852 32370 215904 32376
rect 215760 29708 215812 29714
rect 215760 29650 215812 29656
rect 215668 26920 215720 26926
rect 215668 26862 215720 26868
rect 215956 18698 215984 48418
rect 216140 41414 216168 48894
rect 216324 48346 216352 52158
rect 216588 51740 216640 51746
rect 216588 51682 216640 51688
rect 216404 51604 216456 51610
rect 216404 51546 216456 51552
rect 216416 49881 216444 51546
rect 216600 49978 216628 51682
rect 218072 50726 218100 703582
rect 218808 703474 218836 703582
rect 218950 703520 219062 704960
rect 234632 703582 235028 703610
rect 218992 703474 219020 703520
rect 218808 703446 219020 703474
rect 218704 700664 218756 700670
rect 218704 700606 218756 700612
rect 218152 700324 218204 700330
rect 218152 700266 218204 700272
rect 218060 50720 218112 50726
rect 218060 50662 218112 50668
rect 216588 49972 216640 49978
rect 216588 49914 216640 49920
rect 216402 49872 216458 49881
rect 216402 49807 216458 49816
rect 216680 48408 216732 48414
rect 216680 48350 216732 48356
rect 216312 48340 216364 48346
rect 216312 48282 216364 48288
rect 216048 41386 216168 41414
rect 216048 36786 216076 41386
rect 216036 36780 216088 36786
rect 216036 36722 216088 36728
rect 215944 18692 215996 18698
rect 215944 18634 215996 18640
rect 215576 13116 215628 13122
rect 215576 13058 215628 13064
rect 215484 10328 215536 10334
rect 215484 10270 215536 10276
rect 215392 7608 215444 7614
rect 215392 7550 215444 7556
rect 215300 4820 215352 4826
rect 215300 4762 215352 4768
rect 213184 3936 213236 3942
rect 213184 3878 213236 3884
rect 211804 3528 211856 3534
rect 211804 3470 211856 3476
rect 213368 3528 213420 3534
rect 213368 3470 213420 3476
rect 212172 3392 212224 3398
rect 212172 3334 212224 3340
rect 212184 480 212212 3334
rect 213380 480 213408 3470
rect 215668 3460 215720 3466
rect 215668 3402 215720 3408
rect 214472 2916 214524 2922
rect 214472 2858 214524 2864
rect 214484 480 214512 2858
rect 215680 480 215708 3402
rect 216692 2922 216720 48350
rect 217322 47560 217378 47569
rect 217322 47495 217378 47504
rect 216864 6860 216916 6866
rect 216864 6802 216916 6808
rect 216680 2916 216732 2922
rect 216680 2858 216732 2864
rect 216876 480 216904 6802
rect 217336 3534 217364 47495
rect 218164 47394 218192 700266
rect 218716 52193 218744 700606
rect 233884 700528 233936 700534
rect 233884 700470 233936 700476
rect 232504 700324 232556 700330
rect 232504 700266 232556 700272
rect 221464 683188 221516 683194
rect 221464 683130 221516 683136
rect 220084 632120 220136 632126
rect 220084 632062 220136 632068
rect 219716 413976 219768 413982
rect 219716 413918 219768 413924
rect 219728 413137 219756 413918
rect 219992 413908 220044 413914
rect 219992 413850 220044 413856
rect 219808 413772 219860 413778
rect 219808 413714 219860 413720
rect 219714 413128 219770 413137
rect 219714 413063 219770 413072
rect 219820 412729 219848 413714
rect 220004 413545 220032 413850
rect 219990 413536 220046 413545
rect 219990 413471 220046 413480
rect 219806 412720 219862 412729
rect 219806 412655 219862 412664
rect 220096 412634 220124 632062
rect 220176 590708 220228 590714
rect 220176 590650 220228 590656
rect 220004 412606 220124 412634
rect 219900 412140 219952 412146
rect 219900 412082 219952 412088
rect 219912 411505 219940 412082
rect 219898 411496 219954 411505
rect 219898 411431 219954 411440
rect 219808 411188 219860 411194
rect 219808 411130 219860 411136
rect 219820 410689 219848 411130
rect 219806 410680 219862 410689
rect 219806 410615 219862 410624
rect 219900 409692 219952 409698
rect 219900 409634 219952 409640
rect 219912 408649 219940 409634
rect 220004 409465 220032 412606
rect 220084 411936 220136 411942
rect 220082 411904 220084 411913
rect 220136 411904 220138 411913
rect 220082 411839 220138 411848
rect 220084 410984 220136 410990
rect 220084 410926 220136 410932
rect 220096 410281 220124 410926
rect 220082 410272 220138 410281
rect 220082 410207 220138 410216
rect 220084 409828 220136 409834
rect 220084 409770 220136 409776
rect 219990 409456 220046 409465
rect 219990 409391 220046 409400
rect 220096 409057 220124 409770
rect 220082 409048 220138 409057
rect 220082 408983 220138 408992
rect 219898 408640 219954 408649
rect 219898 408575 219954 408584
rect 220084 408468 220136 408474
rect 220084 408410 220136 408416
rect 219900 408400 219952 408406
rect 219900 408342 219952 408348
rect 219912 407833 219940 408342
rect 219898 407824 219954 407833
rect 219898 407759 219954 407768
rect 220096 407425 220124 408410
rect 220082 407416 220138 407425
rect 220082 407351 220138 407360
rect 220084 407108 220136 407114
rect 220084 407050 220136 407056
rect 219900 406428 219952 406434
rect 219900 406370 219952 406376
rect 219912 406201 219940 406370
rect 219898 406192 219954 406201
rect 219898 406127 219954 406136
rect 220096 405793 220124 407050
rect 220082 405784 220138 405793
rect 220082 405719 220138 405728
rect 220084 405680 220136 405686
rect 220084 405622 220136 405628
rect 219900 405340 219952 405346
rect 219900 405282 219952 405288
rect 219912 404977 219940 405282
rect 219898 404968 219954 404977
rect 219898 404903 219954 404912
rect 220096 404569 220124 405622
rect 220082 404560 220138 404569
rect 220082 404495 220138 404504
rect 219992 404320 220044 404326
rect 219992 404262 220044 404268
rect 220004 403345 220032 404262
rect 220084 404184 220136 404190
rect 220084 404126 220136 404132
rect 220096 403753 220124 404126
rect 220082 403744 220138 403753
rect 220082 403679 220138 403688
rect 219990 403336 220046 403345
rect 219990 403271 220046 403280
rect 220188 402974 220216 590650
rect 220268 581052 220320 581058
rect 220268 580994 220320 581000
rect 219716 402960 219768 402966
rect 219912 402946 220216 402974
rect 219716 402902 219768 402908
rect 219806 402928 219862 402937
rect 219728 402529 219756 402902
rect 219806 402863 219862 402872
rect 219820 402762 219848 402863
rect 219808 402756 219860 402762
rect 219808 402698 219860 402704
rect 219714 402520 219770 402529
rect 219714 402455 219770 402464
rect 219912 396001 219940 402946
rect 220176 402892 220228 402898
rect 220176 402834 220228 402840
rect 220188 401713 220216 402834
rect 220174 401704 220230 401713
rect 220174 401639 220230 401648
rect 220176 401532 220228 401538
rect 220176 401474 220228 401480
rect 220084 401328 220136 401334
rect 220082 401296 220084 401305
rect 220136 401296 220138 401305
rect 220082 401231 220138 401240
rect 220188 400489 220216 401474
rect 220174 400480 220230 400489
rect 220174 400415 220230 400424
rect 220084 400104 220136 400110
rect 219990 400072 220046 400081
rect 220084 400046 220136 400052
rect 219990 400007 220046 400016
rect 220004 399974 220032 400007
rect 219992 399968 220044 399974
rect 219992 399910 220044 399916
rect 220096 399265 220124 400046
rect 220176 400036 220228 400042
rect 220176 399978 220228 399984
rect 220082 399256 220138 399265
rect 220082 399191 220138 399200
rect 220188 398857 220216 399978
rect 220174 398848 220230 398857
rect 220084 398812 220136 398818
rect 220174 398783 220230 398792
rect 220084 398754 220136 398760
rect 220096 398041 220124 398754
rect 220176 398744 220228 398750
rect 220176 398686 220228 398692
rect 220082 398032 220138 398041
rect 220082 397967 220138 397976
rect 220188 397633 220216 398686
rect 220174 397624 220230 397633
rect 220174 397559 220230 397568
rect 220176 397384 220228 397390
rect 220176 397326 220228 397332
rect 220188 396409 220216 397326
rect 220174 396400 220230 396409
rect 220174 396335 220230 396344
rect 220084 396024 220136 396030
rect 219898 395992 219954 396001
rect 220084 395966 220136 395972
rect 219898 395927 219954 395936
rect 220096 395593 220124 395966
rect 220176 395956 220228 395962
rect 220176 395898 220228 395904
rect 220082 395584 220138 395593
rect 220082 395519 220138 395528
rect 220188 395185 220216 395898
rect 220174 395176 220230 395185
rect 220174 395111 220230 395120
rect 219992 394596 220044 394602
rect 219992 394538 220044 394544
rect 220004 393961 220032 394538
rect 220176 394528 220228 394534
rect 220176 394470 220228 394476
rect 219990 393952 220046 393961
rect 219990 393887 220046 393896
rect 220188 393553 220216 394470
rect 220174 393544 220230 393553
rect 220174 393479 220230 393488
rect 220176 393304 220228 393310
rect 220176 393246 220228 393252
rect 220188 392329 220216 393246
rect 220280 392737 220308 580994
rect 220360 571396 220412 571402
rect 220360 571338 220412 571344
rect 220266 392728 220322 392737
rect 220266 392663 220322 392672
rect 220174 392320 220230 392329
rect 220174 392255 220230 392264
rect 220176 392012 220228 392018
rect 220176 391954 220228 391960
rect 219992 390584 220044 390590
rect 219992 390526 220044 390532
rect 219900 390380 219952 390386
rect 219900 390322 219952 390328
rect 219912 389881 219940 390322
rect 219898 389872 219954 389881
rect 219898 389807 219954 389816
rect 219900 389224 219952 389230
rect 219900 389166 219952 389172
rect 219912 383738 219940 389166
rect 220004 383874 220032 390526
rect 220084 389020 220136 389026
rect 220084 388962 220136 388968
rect 220096 388249 220124 388962
rect 220082 388240 220138 388249
rect 220082 388175 220138 388184
rect 220188 387841 220216 391954
rect 220268 391944 220320 391950
rect 220268 391886 220320 391892
rect 220280 391105 220308 391886
rect 220266 391096 220322 391105
rect 220266 391031 220322 391040
rect 220372 389473 220400 571338
rect 220452 567248 220504 567254
rect 220452 567190 220504 567196
rect 220464 392018 220492 567190
rect 220544 550656 220596 550662
rect 220544 550598 220596 550604
rect 220452 392012 220504 392018
rect 220452 391954 220504 391960
rect 220452 391808 220504 391814
rect 220452 391750 220504 391756
rect 220464 390697 220492 391750
rect 220450 390688 220506 390697
rect 220450 390623 220506 390632
rect 220358 389464 220414 389473
rect 220358 389399 220414 389408
rect 220452 389088 220504 389094
rect 220452 389030 220504 389036
rect 220464 388657 220492 389030
rect 220450 388648 220506 388657
rect 220450 388583 220506 388592
rect 220174 387832 220230 387841
rect 220174 387767 220230 387776
rect 220452 387796 220504 387802
rect 220452 387738 220504 387744
rect 220268 387660 220320 387666
rect 220268 387602 220320 387608
rect 220280 387025 220308 387602
rect 220266 387016 220322 387025
rect 220266 386951 220322 386960
rect 220464 386617 220492 387738
rect 220450 386608 220506 386617
rect 220450 386543 220506 386552
rect 220176 386300 220228 386306
rect 220176 386242 220228 386248
rect 220188 385801 220216 386242
rect 220452 386232 220504 386238
rect 220452 386174 220504 386180
rect 220174 385792 220230 385801
rect 220174 385727 220230 385736
rect 220464 385393 220492 386174
rect 220450 385384 220506 385393
rect 220450 385319 220506 385328
rect 220268 385008 220320 385014
rect 220268 384950 220320 384956
rect 220358 384976 220414 384985
rect 220280 384169 220308 384950
rect 220358 384911 220414 384920
rect 220372 384810 220400 384911
rect 220452 384872 220504 384878
rect 220452 384814 220504 384820
rect 220360 384804 220412 384810
rect 220360 384746 220412 384752
rect 220266 384160 220322 384169
rect 220266 384095 220322 384104
rect 220004 383846 220308 383874
rect 219912 383710 220216 383738
rect 220084 383648 220136 383654
rect 220084 383590 220136 383596
rect 220096 383353 220124 383590
rect 220082 383344 220138 383353
rect 220082 383279 220138 383288
rect 219716 380724 219768 380730
rect 219716 380666 219768 380672
rect 219728 380089 219756 380666
rect 219714 380080 219770 380089
rect 219714 380015 219770 380024
rect 220084 378208 220136 378214
rect 220084 378150 220136 378156
rect 219992 376644 220044 376650
rect 219992 376586 220044 376592
rect 219900 376032 219952 376038
rect 220004 376009 220032 376586
rect 219900 375974 219952 375980
rect 219990 376000 220046 376009
rect 219440 374876 219492 374882
rect 219440 374818 219492 374824
rect 219452 374785 219480 374818
rect 219438 374776 219494 374785
rect 219438 374711 219494 374720
rect 219912 373561 219940 375974
rect 219990 375935 220046 375944
rect 219992 375896 220044 375902
rect 219992 375838 220044 375844
rect 220004 375601 220032 375838
rect 219990 375592 220046 375601
rect 219990 375527 220046 375536
rect 219898 373552 219954 373561
rect 219898 373487 219954 373496
rect 219992 372564 220044 372570
rect 219992 372506 220044 372512
rect 218796 371884 218848 371890
rect 218796 371826 218848 371832
rect 218702 52184 218758 52193
rect 218702 52119 218758 52128
rect 218244 49360 218296 49366
rect 218244 49302 218296 49308
rect 218152 47388 218204 47394
rect 218152 47330 218204 47336
rect 218256 6914 218284 49302
rect 218808 48521 218836 371826
rect 220004 371521 220032 372506
rect 219990 371512 220046 371521
rect 219990 371447 220046 371456
rect 219716 370524 219768 370530
rect 219716 370466 219768 370472
rect 219728 368665 219756 370466
rect 219992 369164 220044 369170
rect 219992 369106 220044 369112
rect 219714 368656 219770 368665
rect 219714 368591 219770 368600
rect 219900 368076 219952 368082
rect 219900 368018 219952 368024
rect 219624 367804 219676 367810
rect 219624 367746 219676 367752
rect 219440 366376 219492 366382
rect 219440 366318 219492 366324
rect 219452 358465 219480 366318
rect 219636 365809 219664 367746
rect 219912 367441 219940 368018
rect 219898 367432 219954 367441
rect 219898 367367 219954 367376
rect 219622 365800 219678 365809
rect 219622 365735 219678 365744
rect 219716 365628 219768 365634
rect 219716 365570 219768 365576
rect 219728 364585 219756 365570
rect 220004 365401 220032 369106
rect 219990 365392 220046 365401
rect 219990 365327 220046 365336
rect 219714 364576 219770 364585
rect 219714 364511 219770 364520
rect 219900 361140 219952 361146
rect 219900 361082 219952 361088
rect 219912 360505 219940 361082
rect 219898 360496 219954 360505
rect 219898 360431 219954 360440
rect 219716 360120 219768 360126
rect 219716 360062 219768 360068
rect 219728 358873 219756 360062
rect 219900 359508 219952 359514
rect 219900 359450 219952 359456
rect 219714 358864 219770 358873
rect 219714 358799 219770 358808
rect 219438 358456 219494 358465
rect 219438 358391 219494 358400
rect 219912 356833 219940 359450
rect 219992 358692 220044 358698
rect 219992 358634 220044 358640
rect 220004 357649 220032 358634
rect 219990 357640 220046 357649
rect 219990 357575 220046 357584
rect 219898 356824 219954 356833
rect 219898 356759 219954 356768
rect 219900 356720 219952 356726
rect 219900 356662 219952 356668
rect 219808 355836 219860 355842
rect 219808 355778 219860 355784
rect 219820 354793 219848 355778
rect 219806 354784 219862 354793
rect 219806 354719 219862 354728
rect 219912 351937 219940 356662
rect 219898 351928 219954 351937
rect 219898 351863 219954 351872
rect 219992 351348 220044 351354
rect 219992 351290 220044 351296
rect 220004 351121 220032 351290
rect 219990 351112 220046 351121
rect 219900 351076 219952 351082
rect 219990 351047 220046 351056
rect 219900 351018 219952 351024
rect 219912 350713 219940 351018
rect 219898 350704 219954 350713
rect 219898 350639 219954 350648
rect 219900 350260 219952 350266
rect 219900 350202 219952 350208
rect 219912 349489 219940 350202
rect 219898 349480 219954 349489
rect 219898 349415 219954 349424
rect 219900 343936 219952 343942
rect 219900 343878 219952 343884
rect 219912 343777 219940 343878
rect 219898 343768 219954 343777
rect 219898 343703 219954 343712
rect 219808 341964 219860 341970
rect 219808 341906 219860 341912
rect 219820 341737 219848 341906
rect 219806 341728 219862 341737
rect 219806 341663 219862 341672
rect 219532 340876 219584 340882
rect 219532 340818 219584 340824
rect 219544 339697 219572 340818
rect 219900 340536 219952 340542
rect 219898 340504 219900 340513
rect 219952 340504 219954 340513
rect 219898 340439 219954 340448
rect 219530 339688 219586 339697
rect 219530 339623 219586 339632
rect 219898 338056 219954 338065
rect 219898 337991 219954 338000
rect 219912 334626 219940 337991
rect 219990 334792 220046 334801
rect 219990 334727 220046 334736
rect 219900 334620 219952 334626
rect 219900 334562 219952 334568
rect 220004 334082 220032 334727
rect 219992 334076 220044 334082
rect 219992 334018 220044 334024
rect 219806 333160 219862 333169
rect 219806 333095 219808 333104
rect 219860 333095 219862 333104
rect 219808 333066 219860 333072
rect 219898 332344 219954 332353
rect 219898 332279 219954 332288
rect 219912 331634 219940 332279
rect 219900 331628 219952 331634
rect 219900 331570 219952 331576
rect 219898 331528 219954 331537
rect 219898 331463 219900 331472
rect 219952 331463 219954 331472
rect 219900 331434 219952 331440
rect 219714 330712 219770 330721
rect 219714 330647 219770 330656
rect 219728 330002 219756 330647
rect 219716 329996 219768 330002
rect 219716 329938 219768 329944
rect 219530 329080 219586 329089
rect 219530 329015 219532 329024
rect 219584 329015 219586 329024
rect 219532 328986 219584 328992
rect 219530 327040 219586 327049
rect 219530 326975 219586 326984
rect 219544 324970 219572 326975
rect 219898 325000 219954 325009
rect 219532 324964 219584 324970
rect 219898 324935 219954 324944
rect 219532 324906 219584 324912
rect 219912 324358 219940 324935
rect 219900 324352 219952 324358
rect 219900 324294 219952 324300
rect 219714 323368 219770 323377
rect 219714 323303 219716 323312
rect 219768 323303 219770 323312
rect 219716 323274 219768 323280
rect 218980 320884 219032 320890
rect 218980 320826 219032 320832
rect 218794 48512 218850 48521
rect 218794 48447 218850 48456
rect 218992 48385 219020 320826
rect 219164 319456 219216 319462
rect 219164 319398 219216 319404
rect 219176 49201 219204 319398
rect 219990 318472 220046 318481
rect 219990 318407 219992 318416
rect 220044 318407 220046 318416
rect 219992 318378 220044 318384
rect 219990 315616 220046 315625
rect 219990 315551 220046 315560
rect 220004 314906 220032 315551
rect 219992 314900 220044 314906
rect 219992 314842 220044 314848
rect 219898 313168 219954 313177
rect 219898 313103 219954 313112
rect 219912 312254 219940 313103
rect 219900 312248 219952 312254
rect 219900 312190 219952 312196
rect 219714 309088 219770 309097
rect 219714 309023 219770 309032
rect 219728 307834 219756 309023
rect 219898 308680 219954 308689
rect 219898 308615 219954 308624
rect 219912 308038 219940 308615
rect 219900 308032 219952 308038
rect 219900 307974 219952 307980
rect 219716 307828 219768 307834
rect 219716 307770 219768 307776
rect 219898 302968 219954 302977
rect 219898 302903 219954 302912
rect 219912 302394 219940 302903
rect 219900 302388 219952 302394
rect 219900 302330 219952 302336
rect 219990 301336 220046 301345
rect 219990 301271 220046 301280
rect 220004 301102 220032 301271
rect 219992 301096 220044 301102
rect 219992 301038 220044 301044
rect 219990 298888 220046 298897
rect 219990 298823 220046 298832
rect 220004 298314 220032 298823
rect 219992 298308 220044 298314
rect 219992 298250 220044 298256
rect 219898 296032 219954 296041
rect 219898 295967 219954 295976
rect 219912 295526 219940 295967
rect 219900 295520 219952 295526
rect 219900 295462 219952 295468
rect 219898 294808 219954 294817
rect 219898 294743 219954 294752
rect 219912 294030 219940 294743
rect 219900 294024 219952 294030
rect 219900 293966 219952 293972
rect 219898 292360 219954 292369
rect 219898 292295 219954 292304
rect 219912 291378 219940 292295
rect 219900 291372 219952 291378
rect 219900 291314 219952 291320
rect 219530 288280 219586 288289
rect 219530 288215 219586 288224
rect 219544 287094 219572 288215
rect 219532 287088 219584 287094
rect 219532 287030 219584 287036
rect 219898 287056 219954 287065
rect 219898 286991 219954 287000
rect 219912 286754 219940 286991
rect 219900 286748 219952 286754
rect 219900 286690 219952 286696
rect 219898 286648 219954 286657
rect 219898 286583 219954 286592
rect 219912 286142 219940 286583
rect 219900 286136 219952 286142
rect 219900 286078 219952 286084
rect 220096 50794 220124 378150
rect 220188 340105 220216 383710
rect 220280 340921 220308 383846
rect 220464 383761 220492 384814
rect 220450 383752 220506 383761
rect 220450 383687 220506 383696
rect 220452 383308 220504 383314
rect 220452 383250 220504 383256
rect 220464 382945 220492 383250
rect 220450 382936 220506 382945
rect 220450 382871 220506 382880
rect 220556 382537 220584 550598
rect 220636 535492 220688 535498
rect 220636 535434 220688 535440
rect 220542 382528 220598 382537
rect 220542 382463 220598 382472
rect 220648 382242 220676 535434
rect 220726 413944 220782 413953
rect 220726 413879 220782 413888
rect 220740 413846 220768 413879
rect 220728 413840 220780 413846
rect 220728 413782 220780 413788
rect 220728 412616 220780 412622
rect 220728 412558 220780 412564
rect 220740 412321 220768 412558
rect 220726 412312 220782 412321
rect 220726 412247 220782 412256
rect 220728 411256 220780 411262
rect 220728 411198 220780 411204
rect 220740 411097 220768 411198
rect 220726 411088 220782 411097
rect 220726 411023 220782 411032
rect 220726 409864 220782 409873
rect 220726 409799 220782 409808
rect 220740 409766 220768 409799
rect 220728 409760 220780 409766
rect 220728 409702 220780 409708
rect 220728 408332 220780 408338
rect 220728 408274 220780 408280
rect 220740 408241 220768 408274
rect 220726 408232 220782 408241
rect 220726 408167 220782 408176
rect 220728 407040 220780 407046
rect 220726 407008 220728 407017
rect 220780 407008 220782 407017
rect 220726 406943 220782 406952
rect 220728 406700 220780 406706
rect 220728 406642 220780 406648
rect 220740 406609 220768 406642
rect 220726 406600 220782 406609
rect 220726 406535 220782 406544
rect 220728 405408 220780 405414
rect 220726 405376 220728 405385
rect 220780 405376 220782 405385
rect 220726 405311 220782 405320
rect 220728 404252 220780 404258
rect 220728 404194 220780 404200
rect 220740 404161 220768 404194
rect 220726 404152 220782 404161
rect 220726 404087 220782 404096
rect 220728 402824 220780 402830
rect 220728 402766 220780 402772
rect 220740 402121 220768 402766
rect 220726 402112 220782 402121
rect 220726 402047 220782 402056
rect 220728 401600 220780 401606
rect 220728 401542 220780 401548
rect 220740 400897 220768 401542
rect 220726 400888 220782 400897
rect 220726 400823 220782 400832
rect 220728 400172 220780 400178
rect 220728 400114 220780 400120
rect 220740 399673 220768 400114
rect 220726 399664 220782 399673
rect 220726 399599 220782 399608
rect 220728 398676 220780 398682
rect 220728 398618 220780 398624
rect 220740 398449 220768 398618
rect 220726 398440 220782 398449
rect 220726 398375 220782 398384
rect 220728 397452 220780 397458
rect 220728 397394 220780 397400
rect 220740 397225 220768 397394
rect 220726 397216 220782 397225
rect 220726 397151 220782 397160
rect 220728 396908 220780 396914
rect 220728 396850 220780 396856
rect 220740 396817 220768 396850
rect 220726 396808 220782 396817
rect 220726 396743 220782 396752
rect 220728 395888 220780 395894
rect 220728 395830 220780 395836
rect 220740 394777 220768 395830
rect 220726 394768 220782 394777
rect 220726 394703 220782 394712
rect 220728 394664 220780 394670
rect 220728 394606 220780 394612
rect 220740 394369 220768 394606
rect 220726 394360 220782 394369
rect 220726 394295 220782 394304
rect 220728 393236 220780 393242
rect 220728 393178 220780 393184
rect 220740 393145 220768 393178
rect 220726 393136 220782 393145
rect 220726 393071 220782 393080
rect 220726 391912 220782 391921
rect 220726 391847 220728 391856
rect 220780 391847 220782 391856
rect 220728 391818 220780 391824
rect 220728 391536 220780 391542
rect 220726 391504 220728 391513
rect 220780 391504 220782 391513
rect 220726 391439 220782 391448
rect 220728 390516 220780 390522
rect 220728 390458 220780 390464
rect 220740 390289 220768 390458
rect 220726 390280 220782 390289
rect 220726 390215 220782 390224
rect 220728 389156 220780 389162
rect 220728 389098 220780 389104
rect 220740 389065 220768 389098
rect 220726 389056 220782 389065
rect 220726 388991 220782 389000
rect 220728 387728 220780 387734
rect 220728 387670 220780 387676
rect 220740 387433 220768 387670
rect 220726 387424 220782 387433
rect 220726 387359 220782 387368
rect 220728 386368 220780 386374
rect 220728 386310 220780 386316
rect 220740 386209 220768 386310
rect 220726 386200 220782 386209
rect 220726 386135 220782 386144
rect 220728 384940 220780 384946
rect 220728 384882 220780 384888
rect 220740 384577 220768 384882
rect 220726 384568 220782 384577
rect 220726 384503 220782 384512
rect 220464 382214 220676 382242
rect 220728 382220 220780 382226
rect 220464 376825 220492 382214
rect 220728 382162 220780 382168
rect 220636 382152 220688 382158
rect 220740 382129 220768 382162
rect 220636 382094 220688 382100
rect 220726 382120 220782 382129
rect 220544 382084 220596 382090
rect 220544 382026 220596 382032
rect 220556 381313 220584 382026
rect 220648 381721 220676 382094
rect 220726 382055 220782 382064
rect 220634 381712 220690 381721
rect 220634 381647 220690 381656
rect 220542 381304 220598 381313
rect 220542 381239 220598 381248
rect 220726 380896 220782 380905
rect 220636 380860 220688 380866
rect 220726 380831 220782 380840
rect 220636 380802 220688 380808
rect 220648 379681 220676 380802
rect 220740 380798 220768 380831
rect 220728 380792 220780 380798
rect 220728 380734 220780 380740
rect 220728 380520 220780 380526
rect 220726 380488 220728 380497
rect 220780 380488 220782 380497
rect 220726 380423 220782 380432
rect 220634 379672 220690 379681
rect 220634 379607 220690 379616
rect 220728 379500 220780 379506
rect 220728 379442 220780 379448
rect 220636 379432 220688 379438
rect 220636 379374 220688 379380
rect 220544 379364 220596 379370
rect 220544 379306 220596 379312
rect 220556 378865 220584 379306
rect 220542 378856 220598 378865
rect 220542 378791 220598 378800
rect 220648 378457 220676 379374
rect 220740 379273 220768 379442
rect 220726 379264 220782 379273
rect 220726 379199 220782 379208
rect 220634 378448 220690 378457
rect 220634 378383 220690 378392
rect 220636 378140 220688 378146
rect 220636 378082 220688 378088
rect 220544 378004 220596 378010
rect 220544 377946 220596 377952
rect 220556 377233 220584 377946
rect 220648 377641 220676 378082
rect 220728 378072 220780 378078
rect 220726 378040 220728 378049
rect 220780 378040 220782 378049
rect 220726 377975 220782 377984
rect 220634 377632 220690 377641
rect 220634 377567 220690 377576
rect 220542 377224 220598 377233
rect 220542 377159 220598 377168
rect 220450 376816 220506 376825
rect 220450 376751 220506 376760
rect 220728 376712 220780 376718
rect 220728 376654 220780 376660
rect 220740 376417 220768 376654
rect 220726 376408 220782 376417
rect 220726 376343 220782 376352
rect 220636 375352 220688 375358
rect 220636 375294 220688 375300
rect 220648 374377 220676 375294
rect 220728 375284 220780 375290
rect 220728 375226 220780 375232
rect 220740 375193 220768 375226
rect 220726 375184 220782 375193
rect 220726 375119 220782 375128
rect 220634 374368 220690 374377
rect 220634 374303 220690 374312
rect 220728 373992 220780 373998
rect 220542 373960 220598 373969
rect 220728 373934 220780 373940
rect 220542 373895 220598 373904
rect 220636 373924 220688 373930
rect 220556 373862 220584 373895
rect 220636 373866 220688 373872
rect 220544 373856 220596 373862
rect 220544 373798 220596 373804
rect 220648 373153 220676 373866
rect 220634 373144 220690 373153
rect 220634 373079 220690 373088
rect 220740 372745 220768 373934
rect 220726 372736 220782 372745
rect 220726 372671 220782 372680
rect 220360 372360 220412 372366
rect 220358 372328 220360 372337
rect 220412 372328 220414 372337
rect 220358 372263 220414 372272
rect 220452 372020 220504 372026
rect 220452 371962 220504 371968
rect 220464 371929 220492 371962
rect 220450 371920 220506 371929
rect 220450 371855 220506 371864
rect 220544 371204 220596 371210
rect 220544 371146 220596 371152
rect 220556 370297 220584 371146
rect 220728 371136 220780 371142
rect 220634 371104 220690 371113
rect 220728 371078 220780 371084
rect 220634 371039 220636 371048
rect 220688 371039 220690 371048
rect 220636 371010 220688 371016
rect 220740 370705 220768 371078
rect 220726 370696 220782 370705
rect 220726 370631 220782 370640
rect 220542 370288 220598 370297
rect 220542 370223 220598 370232
rect 220544 370184 220596 370190
rect 220544 370126 220596 370132
rect 220556 369889 220584 370126
rect 220542 369880 220598 369889
rect 220542 369815 220598 369824
rect 220636 369640 220688 369646
rect 220636 369582 220688 369588
rect 220648 369481 220676 369582
rect 220634 369472 220690 369481
rect 220634 369407 220690 369416
rect 220636 369368 220688 369374
rect 220636 369310 220688 369316
rect 220648 369073 220676 369310
rect 220634 369064 220690 369073
rect 220634 368999 220690 369008
rect 220544 368484 220596 368490
rect 220544 368426 220596 368432
rect 220556 367849 220584 368426
rect 220728 368416 220780 368422
rect 220728 368358 220780 368364
rect 220740 368257 220768 368358
rect 220726 368248 220782 368257
rect 220726 368183 220782 368192
rect 220542 367840 220598 367849
rect 220542 367775 220598 367784
rect 220544 367056 220596 367062
rect 220544 366998 220596 367004
rect 220726 367024 220782 367033
rect 220556 366625 220584 366998
rect 220726 366959 220728 366968
rect 220780 366959 220782 366968
rect 220728 366930 220780 366936
rect 220636 366920 220688 366926
rect 220636 366862 220688 366868
rect 220542 366616 220598 366625
rect 220542 366551 220598 366560
rect 220648 366217 220676 366862
rect 220634 366208 220690 366217
rect 220634 366143 220690 366152
rect 220636 365696 220688 365702
rect 220636 365638 220688 365644
rect 220648 364993 220676 365638
rect 220634 364984 220690 364993
rect 220634 364919 220690 364928
rect 220636 364336 220688 364342
rect 220636 364278 220688 364284
rect 220544 364200 220596 364206
rect 220542 364168 220544 364177
rect 220596 364168 220598 364177
rect 220542 364103 220598 364112
rect 220648 363361 220676 364278
rect 220728 364268 220780 364274
rect 220728 364210 220780 364216
rect 220740 363769 220768 364210
rect 220726 363760 220782 363769
rect 220726 363695 220782 363704
rect 220634 363352 220690 363361
rect 220634 363287 220690 363296
rect 220726 362944 220782 362953
rect 220726 362879 220782 362888
rect 220636 362840 220688 362846
rect 220636 362782 220688 362788
rect 220544 362704 220596 362710
rect 220544 362646 220596 362652
rect 220452 362160 220504 362166
rect 220450 362128 220452 362137
rect 220504 362128 220506 362137
rect 220450 362063 220506 362072
rect 220556 361729 220584 362646
rect 220648 362545 220676 362782
rect 220740 362778 220768 362879
rect 220728 362772 220780 362778
rect 220728 362714 220780 362720
rect 220634 362536 220690 362545
rect 220634 362471 220690 362480
rect 220636 362228 220688 362234
rect 220636 362170 220688 362176
rect 220542 361720 220598 361729
rect 220542 361655 220598 361664
rect 220452 360936 220504 360942
rect 220450 360904 220452 360913
rect 220504 360904 220506 360913
rect 220360 360868 220412 360874
rect 220450 360839 220506 360848
rect 220360 360810 220412 360816
rect 220372 350305 220400 360810
rect 220648 360346 220676 362170
rect 220728 361548 220780 361554
rect 220728 361490 220780 361496
rect 220740 361321 220768 361490
rect 220726 361312 220782 361321
rect 220726 361247 220782 361256
rect 220464 360318 220676 360346
rect 220464 354674 220492 360318
rect 220636 360188 220688 360194
rect 220636 360130 220688 360136
rect 220648 360097 220676 360130
rect 220634 360088 220690 360097
rect 220634 360023 220690 360032
rect 220728 360052 220780 360058
rect 220728 359994 220780 360000
rect 220740 359689 220768 359994
rect 220726 359680 220782 359689
rect 220726 359615 220782 359624
rect 220728 359304 220780 359310
rect 220726 359272 220728 359281
rect 220780 359272 220782 359281
rect 220726 359207 220782 359216
rect 220636 358760 220688 358766
rect 220636 358702 220688 358708
rect 220544 358080 220596 358086
rect 220648 358057 220676 358702
rect 220544 358022 220596 358028
rect 220634 358048 220690 358057
rect 220556 355201 220584 358022
rect 220634 357983 220690 357992
rect 220728 357400 220780 357406
rect 220728 357342 220780 357348
rect 220636 357264 220688 357270
rect 220634 357232 220636 357241
rect 220688 357232 220690 357241
rect 220634 357167 220690 357176
rect 220740 356425 220768 357342
rect 220726 356416 220782 356425
rect 220726 356351 220782 356360
rect 220728 356040 220780 356046
rect 220726 356008 220728 356017
rect 220780 356008 220782 356017
rect 220726 355943 220782 355952
rect 220728 355768 220780 355774
rect 220728 355710 220780 355716
rect 220740 355609 220768 355710
rect 220726 355600 220782 355609
rect 220726 355535 220782 355544
rect 220542 355192 220598 355201
rect 220542 355127 220598 355136
rect 220728 354680 220780 354686
rect 220464 354646 220584 354674
rect 220556 353569 220584 354646
rect 220728 354622 220780 354628
rect 220636 354408 220688 354414
rect 220634 354376 220636 354385
rect 220688 354376 220690 354385
rect 220634 354311 220690 354320
rect 220636 354000 220688 354006
rect 220740 353977 220768 354622
rect 220636 353942 220688 353948
rect 220726 353968 220782 353977
rect 220542 353560 220598 353569
rect 220542 353495 220598 353504
rect 220452 352776 220504 352782
rect 220450 352744 220452 352753
rect 220504 352744 220506 352753
rect 220450 352679 220506 352688
rect 220452 352504 220504 352510
rect 220452 352446 220504 352452
rect 220464 352345 220492 352446
rect 220450 352336 220506 352345
rect 220450 352271 220506 352280
rect 220544 350532 220596 350538
rect 220544 350474 220596 350480
rect 220358 350296 220414 350305
rect 220358 350231 220414 350240
rect 220556 349897 220584 350474
rect 220542 349888 220598 349897
rect 220542 349823 220598 349832
rect 220648 349466 220676 353942
rect 220726 353903 220782 353912
rect 220728 353252 220780 353258
rect 220728 353194 220780 353200
rect 220740 353161 220768 353194
rect 220726 353152 220782 353161
rect 220726 353087 220782 353096
rect 220728 351892 220780 351898
rect 220728 351834 220780 351840
rect 220740 351529 220768 351834
rect 220726 351520 220782 351529
rect 220726 351455 220782 351464
rect 220728 349852 220780 349858
rect 220728 349794 220780 349800
rect 220372 349438 220676 349466
rect 220372 345001 220400 349438
rect 220636 349104 220688 349110
rect 220542 349072 220598 349081
rect 220636 349046 220688 349052
rect 220542 349007 220544 349016
rect 220596 349007 220598 349016
rect 220544 348978 220596 348984
rect 220544 348424 220596 348430
rect 220544 348366 220596 348372
rect 220452 348084 220504 348090
rect 220452 348026 220504 348032
rect 220464 347857 220492 348026
rect 220450 347848 220506 347857
rect 220450 347783 220506 347792
rect 220452 347744 220504 347750
rect 220452 347686 220504 347692
rect 220464 347041 220492 347686
rect 220450 347032 220506 347041
rect 220450 346967 220506 346976
rect 220358 344992 220414 345001
rect 220358 344927 220414 344936
rect 220452 342576 220504 342582
rect 220450 342544 220452 342553
rect 220504 342544 220506 342553
rect 220450 342479 220506 342488
rect 220556 341329 220584 348366
rect 220648 348265 220676 349046
rect 220740 348673 220768 349794
rect 220726 348664 220782 348673
rect 220726 348599 220782 348608
rect 220634 348256 220690 348265
rect 220634 348191 220690 348200
rect 220728 347676 220780 347682
rect 220728 347618 220780 347624
rect 220636 347608 220688 347614
rect 220636 347550 220688 347556
rect 220648 346633 220676 347550
rect 220740 347449 220768 347618
rect 220726 347440 220782 347449
rect 220726 347375 220782 347384
rect 220634 346624 220690 346633
rect 220634 346559 220690 346568
rect 220636 346384 220688 346390
rect 220636 346326 220688 346332
rect 220648 345409 220676 346326
rect 220728 346316 220780 346322
rect 220728 346258 220780 346264
rect 220740 346225 220768 346258
rect 220726 346216 220782 346225
rect 220726 346151 220782 346160
rect 220728 345976 220780 345982
rect 220728 345918 220780 345924
rect 220740 345817 220768 345918
rect 220726 345808 220782 345817
rect 220726 345743 220782 345752
rect 220634 345400 220690 345409
rect 220634 345335 220690 345344
rect 220636 345024 220688 345030
rect 220636 344966 220688 344972
rect 220648 344185 220676 344966
rect 220728 344956 220780 344962
rect 220728 344898 220780 344904
rect 220740 344593 220768 344898
rect 220726 344584 220782 344593
rect 220726 344519 220782 344528
rect 220634 344176 220690 344185
rect 220634 344111 220690 344120
rect 220728 343596 220780 343602
rect 220728 343538 220780 343544
rect 220636 343392 220688 343398
rect 220634 343360 220636 343369
rect 220688 343360 220690 343369
rect 220634 343295 220690 343304
rect 220740 342961 220768 343538
rect 220726 342952 220782 342961
rect 220726 342887 220782 342896
rect 220728 342168 220780 342174
rect 220726 342136 220728 342145
rect 220780 342136 220782 342145
rect 220726 342071 220782 342080
rect 220542 341320 220598 341329
rect 220542 341255 220598 341264
rect 220266 340912 220322 340921
rect 220266 340847 220322 340856
rect 220174 340096 220230 340105
rect 220174 340031 220230 340040
rect 220728 339448 220780 339454
rect 220728 339390 220780 339396
rect 220636 339380 220688 339386
rect 220636 339322 220688 339328
rect 220452 339312 220504 339318
rect 220452 339254 220504 339260
rect 220464 338473 220492 339254
rect 220648 338881 220676 339322
rect 220740 339289 220768 339390
rect 220726 339280 220782 339289
rect 220726 339215 220782 339224
rect 220634 338872 220690 338881
rect 220634 338807 220690 338816
rect 220450 338464 220506 338473
rect 220450 338399 220506 338408
rect 220634 337648 220690 337657
rect 220634 337583 220690 337592
rect 220544 336932 220596 336938
rect 220544 336874 220596 336880
rect 220556 336841 220584 336874
rect 220542 336832 220598 336841
rect 220648 336802 220676 337583
rect 220726 337240 220782 337249
rect 220726 337175 220782 337184
rect 220740 336870 220768 337175
rect 220728 336864 220780 336870
rect 220728 336806 220780 336812
rect 220542 336767 220598 336776
rect 220636 336796 220688 336802
rect 220636 336738 220688 336744
rect 220634 336424 220690 336433
rect 220634 336359 220690 336368
rect 220648 336122 220676 336359
rect 220636 336116 220688 336122
rect 220636 336058 220688 336064
rect 220542 336016 220598 336025
rect 220542 335951 220598 335960
rect 220556 335510 220584 335951
rect 220726 335608 220782 335617
rect 220726 335543 220728 335552
rect 220780 335543 220782 335552
rect 220728 335514 220780 335520
rect 220544 335504 220596 335510
rect 220544 335446 220596 335452
rect 220174 335200 220230 335209
rect 220174 335135 220230 335144
rect 220188 320074 220216 335135
rect 220358 334384 220414 334393
rect 220358 334319 220414 334328
rect 220372 334014 220400 334319
rect 220360 334008 220412 334014
rect 220360 333950 220412 333956
rect 220450 333976 220506 333985
rect 220450 333911 220506 333920
rect 220464 331906 220492 333911
rect 220634 333568 220690 333577
rect 220634 333503 220690 333512
rect 220648 332722 220676 333503
rect 220726 332752 220782 332761
rect 220636 332716 220688 332722
rect 220726 332687 220782 332696
rect 220636 332658 220688 332664
rect 220740 332654 220768 332687
rect 220728 332648 220780 332654
rect 220728 332590 220780 332596
rect 220542 331936 220598 331945
rect 220452 331900 220504 331906
rect 220542 331871 220598 331880
rect 220452 331842 220504 331848
rect 220556 331294 220584 331871
rect 220544 331288 220596 331294
rect 220544 331230 220596 331236
rect 220542 331120 220598 331129
rect 220542 331055 220598 331064
rect 220556 329934 220584 331055
rect 220726 330304 220782 330313
rect 220726 330239 220782 330248
rect 220544 329928 220596 329934
rect 220544 329870 220596 329876
rect 220634 329896 220690 329905
rect 220740 329866 220768 330239
rect 220634 329831 220690 329840
rect 220728 329860 220780 329866
rect 220542 329488 220598 329497
rect 220542 329423 220598 329432
rect 220556 328506 220584 329423
rect 220648 329118 220676 329831
rect 220728 329802 220780 329808
rect 220636 329112 220688 329118
rect 220636 329054 220688 329060
rect 220726 328672 220782 328681
rect 220726 328607 220782 328616
rect 220740 328574 220768 328607
rect 220728 328568 220780 328574
rect 220728 328510 220780 328516
rect 220544 328500 220596 328506
rect 220544 328442 220596 328448
rect 220266 328264 220322 328273
rect 220266 328199 220322 328208
rect 220280 327962 220308 328199
rect 220268 327956 220320 327962
rect 220268 327898 220320 327904
rect 220266 327856 220322 327865
rect 220266 327791 220322 327800
rect 220280 327214 220308 327791
rect 220726 327448 220782 327457
rect 220726 327383 220782 327392
rect 220268 327208 220320 327214
rect 220268 327150 220320 327156
rect 220740 327146 220768 327383
rect 220728 327140 220780 327146
rect 220728 327082 220780 327088
rect 220634 326632 220690 326641
rect 220634 326567 220690 326576
rect 220358 326224 220414 326233
rect 220358 326159 220414 326168
rect 220372 325922 220400 326159
rect 220360 325916 220412 325922
rect 220360 325858 220412 325864
rect 220648 325718 220676 326567
rect 220726 325816 220782 325825
rect 220726 325751 220728 325760
rect 220780 325751 220782 325760
rect 220728 325722 220780 325728
rect 220636 325712 220688 325718
rect 220636 325654 220688 325660
rect 220266 325408 220322 325417
rect 220266 325343 220322 325352
rect 220280 324494 220308 325343
rect 220728 324624 220780 324630
rect 220726 324592 220728 324601
rect 220780 324592 220782 324601
rect 220726 324527 220782 324536
rect 220268 324488 220320 324494
rect 220268 324430 220320 324436
rect 220360 324420 220412 324426
rect 220360 324362 220412 324368
rect 220266 324184 220322 324193
rect 220266 324119 220322 324128
rect 220280 323134 220308 324119
rect 220268 323128 220320 323134
rect 220268 323070 220320 323076
rect 220266 321328 220322 321337
rect 220266 321263 220322 321272
rect 220280 320618 220308 321263
rect 220268 320612 220320 320618
rect 220268 320554 220320 320560
rect 220266 320512 220322 320521
rect 220266 320447 220322 320456
rect 220280 320278 220308 320447
rect 220268 320272 220320 320278
rect 220268 320214 220320 320220
rect 220176 320068 220228 320074
rect 220176 320010 220228 320016
rect 220372 319954 220400 324362
rect 220634 323776 220690 323785
rect 220634 323711 220690 323720
rect 220648 322998 220676 323711
rect 220728 323060 220780 323066
rect 220728 323002 220780 323008
rect 220636 322992 220688 322998
rect 220740 322969 220768 323002
rect 220636 322934 220688 322940
rect 220726 322960 220782 322969
rect 220726 322895 220782 322904
rect 220542 322552 220598 322561
rect 220542 322487 220598 322496
rect 220556 321774 220584 322487
rect 220634 322144 220690 322153
rect 220634 322079 220690 322088
rect 220544 321768 220596 321774
rect 220544 321710 220596 321716
rect 220648 321638 220676 322079
rect 220726 321736 220782 321745
rect 220726 321671 220728 321680
rect 220780 321671 220782 321680
rect 220728 321642 220780 321648
rect 220636 321632 220688 321638
rect 220636 321574 220688 321580
rect 220726 320920 220782 320929
rect 220726 320855 220782 320864
rect 220740 320210 220768 320855
rect 220728 320204 220780 320210
rect 220728 320146 220780 320152
rect 220450 320104 220506 320113
rect 220450 320039 220506 320048
rect 220188 319926 220400 319954
rect 220188 50862 220216 319926
rect 220268 319864 220320 319870
rect 220268 319806 220320 319812
rect 220280 296682 220308 319806
rect 220464 319802 220492 320039
rect 220452 319796 220504 319802
rect 220452 319738 220504 319744
rect 220450 319696 220506 319705
rect 220450 319631 220506 319640
rect 220358 319288 220414 319297
rect 220358 319223 220414 319232
rect 220372 318850 220400 319223
rect 220464 318918 220492 319631
rect 220728 319048 220780 319054
rect 220728 318990 220780 318996
rect 220452 318912 220504 318918
rect 220740 318889 220768 318990
rect 220452 318854 220504 318860
rect 220726 318880 220782 318889
rect 220360 318844 220412 318850
rect 220726 318815 220782 318824
rect 220360 318786 220412 318792
rect 220634 318064 220690 318073
rect 220634 317999 220690 318008
rect 220648 317558 220676 317999
rect 220726 317656 220782 317665
rect 220726 317591 220782 317600
rect 220636 317552 220688 317558
rect 220636 317494 220688 317500
rect 220740 317490 220768 317591
rect 220728 317484 220780 317490
rect 220728 317426 220780 317432
rect 220726 317248 220782 317257
rect 220726 317183 220782 317192
rect 220634 316840 220690 316849
rect 220634 316775 220690 316784
rect 220648 316538 220676 316775
rect 220636 316532 220688 316538
rect 220636 316474 220688 316480
rect 220450 316432 220506 316441
rect 220450 316367 220506 316376
rect 220464 316130 220492 316367
rect 220452 316124 220504 316130
rect 220452 316066 220504 316072
rect 220740 316062 220768 317183
rect 220728 316056 220780 316062
rect 220634 316024 220690 316033
rect 220728 315998 220780 316004
rect 220634 315959 220690 315968
rect 220544 314832 220596 314838
rect 220542 314800 220544 314809
rect 220596 314800 220598 314809
rect 220648 314770 220676 315959
rect 220726 315208 220782 315217
rect 220726 315143 220782 315152
rect 220542 314735 220598 314744
rect 220636 314764 220688 314770
rect 220636 314706 220688 314712
rect 220740 314702 220768 315143
rect 220728 314696 220780 314702
rect 220728 314638 220780 314644
rect 220634 314392 220690 314401
rect 220634 314327 220690 314336
rect 220450 313984 220506 313993
rect 220450 313919 220506 313928
rect 220464 313410 220492 313919
rect 220452 313404 220504 313410
rect 220452 313346 220504 313352
rect 220648 313342 220676 314327
rect 220726 313576 220782 313585
rect 220726 313511 220782 313520
rect 220740 313478 220768 313511
rect 220728 313472 220780 313478
rect 220728 313414 220780 313420
rect 220636 313336 220688 313342
rect 220636 313278 220688 313284
rect 220450 312760 220506 312769
rect 220450 312695 220506 312704
rect 220464 312458 220492 312695
rect 220452 312452 220504 312458
rect 220452 312394 220504 312400
rect 220450 312352 220506 312361
rect 220450 312287 220506 312296
rect 220464 311914 220492 312287
rect 220728 311976 220780 311982
rect 220726 311944 220728 311953
rect 220780 311944 220782 311953
rect 220452 311908 220504 311914
rect 220726 311879 220782 311888
rect 220452 311850 220504 311856
rect 220634 311536 220690 311545
rect 220634 311471 220690 311480
rect 220542 310720 220598 310729
rect 220542 310655 220544 310664
rect 220596 310655 220598 310664
rect 220544 310626 220596 310632
rect 220648 310554 220676 311471
rect 220726 311128 220782 311137
rect 220726 311063 220782 311072
rect 220740 310622 220768 311063
rect 220728 310616 220780 310622
rect 220728 310558 220780 310564
rect 220636 310548 220688 310554
rect 220636 310490 220688 310496
rect 220726 310312 220782 310321
rect 220726 310247 220782 310256
rect 220542 309904 220598 309913
rect 220542 309839 220598 309848
rect 220556 309262 220584 309839
rect 220634 309496 220690 309505
rect 220634 309431 220636 309440
rect 220688 309431 220690 309440
rect 220636 309402 220688 309408
rect 220544 309256 220596 309262
rect 220544 309198 220596 309204
rect 220740 309194 220768 310247
rect 220728 309188 220780 309194
rect 220728 309130 220780 309136
rect 220634 308272 220690 308281
rect 220634 308207 220690 308216
rect 220648 307902 220676 308207
rect 220728 307964 220780 307970
rect 220728 307906 220780 307912
rect 220636 307896 220688 307902
rect 220740 307873 220768 307906
rect 220636 307838 220688 307844
rect 220726 307864 220782 307873
rect 220726 307799 220782 307808
rect 220542 307456 220598 307465
rect 220542 307391 220598 307400
rect 220556 306542 220584 307391
rect 220634 307048 220690 307057
rect 220634 306983 220690 306992
rect 220544 306536 220596 306542
rect 220544 306478 220596 306484
rect 220648 306406 220676 306983
rect 220726 306640 220782 306649
rect 220726 306575 220782 306584
rect 220740 306474 220768 306575
rect 220728 306468 220780 306474
rect 220728 306410 220780 306416
rect 220636 306400 220688 306406
rect 220636 306342 220688 306348
rect 220542 306232 220598 306241
rect 220542 306167 220598 306176
rect 220556 305046 220584 306167
rect 220634 305824 220690 305833
rect 220634 305759 220690 305768
rect 220648 305114 220676 305759
rect 220726 305416 220782 305425
rect 220726 305351 220728 305360
rect 220780 305351 220782 305360
rect 220728 305322 220780 305328
rect 220728 305176 220780 305182
rect 220728 305118 220780 305124
rect 220636 305108 220688 305114
rect 220636 305050 220688 305056
rect 220544 305040 220596 305046
rect 220740 305017 220768 305118
rect 220544 304982 220596 304988
rect 220726 305008 220782 305017
rect 220726 304943 220782 304952
rect 220450 304600 220506 304609
rect 220450 304535 220506 304544
rect 220464 303686 220492 304535
rect 220634 304192 220690 304201
rect 220634 304127 220690 304136
rect 220648 303822 220676 304127
rect 220636 303816 220688 303822
rect 220636 303758 220688 303764
rect 220726 303784 220782 303793
rect 220726 303719 220728 303728
rect 220780 303719 220782 303728
rect 220728 303690 220780 303696
rect 220452 303680 220504 303686
rect 220452 303622 220504 303628
rect 220542 303376 220598 303385
rect 220542 303311 220598 303320
rect 220556 302326 220584 303311
rect 220726 302560 220782 302569
rect 220726 302495 220782 302504
rect 220544 302320 220596 302326
rect 220544 302262 220596 302268
rect 220740 302258 220768 302495
rect 220728 302252 220780 302258
rect 220728 302194 220780 302200
rect 220634 302152 220690 302161
rect 220634 302087 220690 302096
rect 220542 301744 220598 301753
rect 220542 301679 220598 301688
rect 220556 300966 220584 301679
rect 220544 300960 220596 300966
rect 220544 300902 220596 300908
rect 220648 300898 220676 302087
rect 220728 301028 220780 301034
rect 220728 300970 220780 300976
rect 220740 300937 220768 300970
rect 220726 300928 220782 300937
rect 220636 300892 220688 300898
rect 220726 300863 220782 300872
rect 220636 300834 220688 300840
rect 220634 300112 220690 300121
rect 220634 300047 220690 300056
rect 220648 299606 220676 300047
rect 220726 299704 220782 299713
rect 220726 299639 220782 299648
rect 220636 299600 220688 299606
rect 220636 299542 220688 299548
rect 220740 299538 220768 299639
rect 220728 299532 220780 299538
rect 220728 299474 220780 299480
rect 220542 299296 220598 299305
rect 220542 299231 220598 299240
rect 220556 298246 220584 299231
rect 220726 298480 220782 298489
rect 220726 298415 220782 298424
rect 220544 298240 220596 298246
rect 220544 298182 220596 298188
rect 220740 298178 220768 298415
rect 220728 298172 220780 298178
rect 220728 298114 220780 298120
rect 220634 298072 220690 298081
rect 220634 298007 220690 298016
rect 220358 296848 220414 296857
rect 220358 296783 220414 296792
rect 220268 296676 220320 296682
rect 220268 296618 220320 296624
rect 220266 295216 220322 295225
rect 220266 295151 220322 295160
rect 220280 294234 220308 295151
rect 220268 294228 220320 294234
rect 220268 294170 220320 294176
rect 220266 290320 220322 290329
rect 220266 290255 220322 290264
rect 220280 77246 220308 290255
rect 220372 104854 220400 296783
rect 220648 296750 220676 298007
rect 220726 297664 220782 297673
rect 220726 297599 220728 297608
rect 220780 297599 220782 297608
rect 220728 297570 220780 297576
rect 220726 297256 220782 297265
rect 220726 297191 220782 297200
rect 220740 296818 220768 297191
rect 220728 296812 220780 296818
rect 220728 296754 220780 296760
rect 220636 296744 220688 296750
rect 220636 296686 220688 296692
rect 220634 296440 220690 296449
rect 220634 296375 220690 296384
rect 220648 295458 220676 296375
rect 220726 295624 220782 295633
rect 220726 295559 220782 295568
rect 220636 295452 220688 295458
rect 220636 295394 220688 295400
rect 220740 295390 220768 295559
rect 220728 295384 220780 295390
rect 220728 295326 220780 295332
rect 220726 294400 220782 294409
rect 220726 294335 220782 294344
rect 220740 294166 220768 294335
rect 220728 294160 220780 294166
rect 220728 294102 220780 294108
rect 220450 293992 220506 294001
rect 220450 293927 220506 293936
rect 220464 119882 220492 293927
rect 220634 293584 220690 293593
rect 220634 293519 220690 293528
rect 220542 292768 220598 292777
rect 220542 292703 220544 292712
rect 220596 292703 220598 292712
rect 220544 292674 220596 292680
rect 220648 292602 220676 293519
rect 220726 293176 220782 293185
rect 220726 293111 220782 293120
rect 220740 292670 220768 293111
rect 220728 292664 220780 292670
rect 220728 292606 220780 292612
rect 220636 292596 220688 292602
rect 220636 292538 220688 292544
rect 220634 291952 220690 291961
rect 220634 291887 220690 291896
rect 220648 291310 220676 291887
rect 220726 291544 220782 291553
rect 220726 291479 220782 291488
rect 220636 291304 220688 291310
rect 220636 291246 220688 291252
rect 220740 291242 220768 291479
rect 220728 291236 220780 291242
rect 220728 291178 220780 291184
rect 220726 291136 220782 291145
rect 220726 291071 220782 291080
rect 220634 290728 220690 290737
rect 220634 290663 220690 290672
rect 220648 289950 220676 290663
rect 220740 290018 220768 291071
rect 220728 290012 220780 290018
rect 220728 289954 220780 289960
rect 220636 289944 220688 289950
rect 220636 289886 220688 289892
rect 220726 289912 220782 289921
rect 220726 289847 220728 289856
rect 220780 289847 220782 289856
rect 220728 289818 220780 289824
rect 220542 289504 220598 289513
rect 220542 289439 220598 289448
rect 220556 288590 220584 289439
rect 220634 289096 220690 289105
rect 220634 289031 220690 289040
rect 220544 288584 220596 288590
rect 220544 288526 220596 288532
rect 220648 288522 220676 289031
rect 220726 288688 220782 288697
rect 220726 288623 220782 288632
rect 220636 288516 220688 288522
rect 220636 288458 220688 288464
rect 220740 288454 220768 288623
rect 220728 288448 220780 288454
rect 220728 288390 220780 288396
rect 220634 287872 220690 287881
rect 220634 287807 220690 287816
rect 220648 287162 220676 287807
rect 220726 287464 220782 287473
rect 220726 287399 220728 287408
rect 220780 287399 220782 287408
rect 220728 287370 220780 287376
rect 220636 287156 220688 287162
rect 220636 287098 220688 287104
rect 220634 286240 220690 286249
rect 220634 286175 220690 286184
rect 220648 285802 220676 286175
rect 220728 285932 220780 285938
rect 220728 285874 220780 285880
rect 220740 285841 220768 285874
rect 220726 285832 220782 285841
rect 220636 285796 220688 285802
rect 220726 285767 220782 285776
rect 220636 285738 220688 285744
rect 220452 119876 220504 119882
rect 220452 119818 220504 119824
rect 220360 104848 220412 104854
rect 220360 104790 220412 104796
rect 220268 77240 220320 77246
rect 220268 77182 220320 77188
rect 220820 51128 220872 51134
rect 220820 51070 220872 51076
rect 220176 50856 220228 50862
rect 220176 50798 220228 50804
rect 220084 50788 220136 50794
rect 220084 50730 220136 50736
rect 220176 49836 220228 49842
rect 220176 49778 220228 49784
rect 220188 49502 220216 49778
rect 220176 49496 220228 49502
rect 220176 49438 220228 49444
rect 219162 49192 219218 49201
rect 219162 49127 219218 49136
rect 218978 48376 219034 48385
rect 218978 48311 219034 48320
rect 220832 16574 220860 51070
rect 221476 50289 221504 683130
rect 231124 641776 231176 641782
rect 231124 641718 231176 641724
rect 224224 638988 224276 638994
rect 224224 638930 224276 638936
rect 222844 629332 222896 629338
rect 222844 629274 222896 629280
rect 221648 616888 221700 616894
rect 221648 616830 221700 616836
rect 221556 524476 221608 524482
rect 221556 524418 221608 524424
rect 221568 51649 221596 524418
rect 221660 405686 221688 616830
rect 221740 612808 221792 612814
rect 221740 612750 221792 612756
rect 221648 405680 221700 405686
rect 221648 405622 221700 405628
rect 221752 402762 221780 612750
rect 221832 607232 221884 607238
rect 221832 607174 221884 607180
rect 221740 402756 221792 402762
rect 221740 402698 221792 402704
rect 221844 401334 221872 607174
rect 221924 552084 221976 552090
rect 221924 552026 221976 552032
rect 221832 401328 221884 401334
rect 221832 401270 221884 401276
rect 221740 394732 221792 394738
rect 221740 394674 221792 394680
rect 221648 393372 221700 393378
rect 221648 393314 221700 393320
rect 221660 341970 221688 393314
rect 221752 342582 221780 394674
rect 221936 383314 221964 552026
rect 222016 438932 222068 438938
rect 222016 438874 222068 438880
rect 221924 383308 221976 383314
rect 221924 383250 221976 383256
rect 222028 357270 222056 438874
rect 222752 425128 222804 425134
rect 222752 425070 222804 425076
rect 222108 404388 222160 404394
rect 222108 404330 222160 404336
rect 222016 357264 222068 357270
rect 222016 357206 222068 357212
rect 222120 345982 222148 404330
rect 222764 352510 222792 425070
rect 222856 409698 222884 629274
rect 222936 622464 222988 622470
rect 222936 622406 222988 622412
rect 222844 409692 222896 409698
rect 222844 409634 222896 409640
rect 222948 406434 222976 622406
rect 223028 593428 223080 593434
rect 223028 593370 223080 593376
rect 222936 406428 222988 406434
rect 222936 406370 222988 406376
rect 222844 397520 222896 397526
rect 222844 397462 222896 397468
rect 222752 352504 222804 352510
rect 222752 352446 222804 352452
rect 222108 345976 222160 345982
rect 222108 345918 222160 345924
rect 222856 343398 222884 397462
rect 223040 396914 223068 593370
rect 223120 557592 223172 557598
rect 223120 557534 223172 557540
rect 223028 396908 223080 396914
rect 223028 396850 223080 396856
rect 223132 384810 223160 557534
rect 223304 477556 223356 477562
rect 223304 477498 223356 477504
rect 223212 476128 223264 476134
rect 223212 476070 223264 476076
rect 223120 384804 223172 384810
rect 223120 384746 223172 384752
rect 223224 369646 223252 476070
rect 223316 370190 223344 477498
rect 223396 454096 223448 454102
rect 223396 454038 223448 454044
rect 223304 370184 223356 370190
rect 223304 370126 223356 370132
rect 223212 369640 223264 369646
rect 223212 369582 223264 369588
rect 223408 362166 223436 454038
rect 223488 448588 223540 448594
rect 223488 448530 223540 448536
rect 223396 362160 223448 362166
rect 223396 362102 223448 362108
rect 223500 361146 223528 448530
rect 224132 431996 224184 432002
rect 224132 431938 224184 431944
rect 224040 415472 224092 415478
rect 224040 415414 224092 415420
rect 223948 411324 224000 411330
rect 223948 411266 224000 411272
rect 223488 361140 223540 361146
rect 223488 361082 223540 361088
rect 223960 348090 223988 411266
rect 224052 349042 224080 415414
rect 224144 355842 224172 431938
rect 224236 411942 224264 638930
rect 228364 637628 228416 637634
rect 228364 637570 228416 637576
rect 225604 633480 225656 633486
rect 225604 633422 225656 633428
rect 224316 618316 224368 618322
rect 224316 618258 224368 618264
rect 224224 411936 224276 411942
rect 224224 411878 224276 411884
rect 224328 405346 224356 618258
rect 224408 489932 224460 489938
rect 224408 489874 224460 489880
rect 224316 405340 224368 405346
rect 224316 405282 224368 405288
rect 224420 373862 224448 489874
rect 224500 484424 224552 484430
rect 224500 484366 224552 484372
rect 224408 373856 224460 373862
rect 224408 373798 224460 373804
rect 224512 372366 224540 484366
rect 224592 483064 224644 483070
rect 224592 483006 224644 483012
rect 224500 372360 224552 372366
rect 224500 372302 224552 372308
rect 224604 372026 224632 483006
rect 224776 481704 224828 481710
rect 224776 481646 224828 481652
rect 224684 480276 224736 480282
rect 224684 480218 224736 480224
rect 224592 372020 224644 372026
rect 224592 371962 224644 371968
rect 224696 371074 224724 480218
rect 224788 372570 224816 481646
rect 224868 472048 224920 472054
rect 224868 471990 224920 471996
rect 224776 372564 224828 372570
rect 224776 372506 224828 372512
rect 224684 371068 224736 371074
rect 224684 371010 224736 371016
rect 224880 368422 224908 471990
rect 225616 410990 225644 633422
rect 226984 619676 227036 619682
rect 226984 619618 227036 619624
rect 225696 568608 225748 568614
rect 225696 568550 225748 568556
rect 225604 410984 225656 410990
rect 225604 410926 225656 410932
rect 225708 389026 225736 568550
rect 225788 495508 225840 495514
rect 225788 495450 225840 495456
rect 225696 389020 225748 389026
rect 225696 388962 225748 388968
rect 225800 376650 225828 495450
rect 225880 494080 225932 494086
rect 225880 494022 225932 494028
rect 225788 376644 225840 376650
rect 225788 376586 225840 376592
rect 225892 375902 225920 494022
rect 225972 491360 226024 491366
rect 225972 491302 226024 491308
rect 225880 375896 225932 375902
rect 225880 375838 225932 375844
rect 225984 374882 226012 491302
rect 226064 459604 226116 459610
rect 226064 459546 226116 459552
rect 225972 374876 226024 374882
rect 225972 374818 226024 374824
rect 224868 368416 224920 368422
rect 224868 368358 224920 368364
rect 226076 364206 226104 459546
rect 226892 449948 226944 449954
rect 226892 449890 226944 449896
rect 226800 445800 226852 445806
rect 226800 445742 226852 445748
rect 226156 434784 226208 434790
rect 226156 434726 226208 434732
rect 226064 364200 226116 364206
rect 226064 364142 226116 364148
rect 224132 355836 224184 355842
rect 224132 355778 224184 355784
rect 226168 355774 226196 434726
rect 226248 419552 226300 419558
rect 226248 419494 226300 419500
rect 226156 355768 226208 355774
rect 226156 355710 226208 355716
rect 226260 351082 226288 419494
rect 226812 359310 226840 445742
rect 226904 360942 226932 449890
rect 226996 405414 227024 619618
rect 227076 603152 227128 603158
rect 227076 603094 227128 603100
rect 226984 405408 227036 405414
rect 226984 405350 227036 405356
rect 227088 399974 227116 603094
rect 227168 578264 227220 578270
rect 227168 578206 227220 578212
rect 227076 399968 227128 399974
rect 227076 399910 227128 399916
rect 226984 398880 227036 398886
rect 226984 398822 227036 398828
rect 226892 360936 226944 360942
rect 226892 360878 226944 360884
rect 226800 359304 226852 359310
rect 226800 359246 226852 359252
rect 226248 351076 226300 351082
rect 226248 351018 226300 351024
rect 224040 349036 224092 349042
rect 224040 348978 224092 348984
rect 223948 348084 224000 348090
rect 223948 348026 224000 348032
rect 226996 343942 227024 398822
rect 227180 391542 227208 578206
rect 227260 572756 227312 572762
rect 227260 572698 227312 572704
rect 227168 391536 227220 391542
rect 227168 391478 227220 391484
rect 227272 390386 227300 572698
rect 227352 545148 227404 545154
rect 227352 545090 227404 545096
rect 227260 390380 227312 390386
rect 227260 390322 227312 390328
rect 227076 383716 227128 383722
rect 227076 383658 227128 383664
rect 226984 343936 227036 343942
rect 226984 343878 227036 343884
rect 222844 343392 222896 343398
rect 222844 343334 222896 343340
rect 221740 342576 221792 342582
rect 221740 342518 221792 342524
rect 221648 341964 221700 341970
rect 221648 341906 221700 341912
rect 227088 340542 227116 383658
rect 227364 380526 227392 545090
rect 227444 543788 227496 543794
rect 227444 543730 227496 543736
rect 227456 380730 227484 543730
rect 227536 474768 227588 474774
rect 227536 474710 227588 474716
rect 227444 380724 227496 380730
rect 227444 380666 227496 380672
rect 227352 380520 227404 380526
rect 227352 380462 227404 380468
rect 227548 369374 227576 474710
rect 227628 469260 227680 469266
rect 227628 469202 227680 469208
rect 227536 369368 227588 369374
rect 227536 369310 227588 369316
rect 227640 368082 227668 469202
rect 228376 412146 228404 637570
rect 228456 632732 228508 632738
rect 228456 632674 228508 632680
rect 228364 412140 228416 412146
rect 228364 412082 228416 412088
rect 228468 409766 228496 632674
rect 228548 623824 228600 623830
rect 228548 623766 228600 623772
rect 228456 409760 228508 409766
rect 228456 409702 228508 409708
rect 228560 406706 228588 623766
rect 229744 610020 229796 610026
rect 229744 609962 229796 609968
rect 228640 440292 228692 440298
rect 228640 440234 228692 440240
rect 228548 406700 228600 406706
rect 228548 406642 228600 406648
rect 227628 368076 227680 368082
rect 227628 368018 227680 368024
rect 228652 358698 228680 440234
rect 228732 430636 228784 430642
rect 228732 430578 228784 430584
rect 228640 358692 228692 358698
rect 228640 358634 228692 358640
rect 228744 354414 228772 430578
rect 228824 426488 228876 426494
rect 228824 426430 228876 426436
rect 228732 354408 228784 354414
rect 228732 354350 228784 354356
rect 228836 352782 228864 426430
rect 228916 420980 228968 420986
rect 228916 420922 228968 420928
rect 228824 352776 228876 352782
rect 228824 352718 228876 352724
rect 228928 351354 228956 420922
rect 229008 415540 229060 415546
rect 229008 415482 229060 415488
rect 228916 351348 228968 351354
rect 228916 351290 228968 351296
rect 229020 350266 229048 415482
rect 229756 402830 229784 609962
rect 229836 608660 229888 608666
rect 229836 608602 229888 608608
rect 229848 402898 229876 608602
rect 229928 587920 229980 587926
rect 229928 587862 229980 587868
rect 229836 402892 229888 402898
rect 229836 402834 229888 402840
rect 229744 402824 229796 402830
rect 229744 402766 229796 402772
rect 229744 400920 229796 400926
rect 229744 400862 229796 400868
rect 229008 350260 229060 350266
rect 229008 350202 229060 350208
rect 229756 346322 229784 400862
rect 229940 395894 229968 587862
rect 230020 582412 230072 582418
rect 230020 582354 230072 582360
rect 229928 395888 229980 395894
rect 229928 395830 229980 395836
rect 230032 393242 230060 582354
rect 230112 470620 230164 470626
rect 230112 470562 230164 470568
rect 230020 393236 230072 393242
rect 230020 393178 230072 393184
rect 230124 368490 230152 470562
rect 230204 466472 230256 466478
rect 230204 466414 230256 466420
rect 230112 368484 230164 368490
rect 230112 368426 230164 368432
rect 230216 366926 230244 466414
rect 230296 439544 230348 439550
rect 230296 439486 230348 439492
rect 230204 366920 230256 366926
rect 230204 366862 230256 366868
rect 230308 365634 230336 439486
rect 231136 413778 231164 641718
rect 231216 627972 231268 627978
rect 231216 627914 231268 627920
rect 231124 413772 231176 413778
rect 231124 413714 231176 413720
rect 231228 408338 231256 627914
rect 231308 626612 231360 626618
rect 231308 626554 231360 626560
rect 231320 408406 231348 626554
rect 231400 574116 231452 574122
rect 231400 574058 231452 574064
rect 231308 408400 231360 408406
rect 231308 408342 231360 408348
rect 231216 408332 231268 408338
rect 231216 408274 231268 408280
rect 231032 407176 231084 407182
rect 231032 407118 231084 407124
rect 230296 365628 230348 365634
rect 230296 365570 230348 365576
rect 231044 347614 231072 407118
rect 231216 401668 231268 401674
rect 231216 401610 231268 401616
rect 231124 364404 231176 364410
rect 231124 364346 231176 364352
rect 231032 347608 231084 347614
rect 231032 347550 231084 347556
rect 229744 346316 229796 346322
rect 229744 346258 229796 346264
rect 227076 340536 227128 340542
rect 227076 340478 227128 340484
rect 227076 336932 227128 336938
rect 227076 336874 227128 336880
rect 223948 336116 224000 336122
rect 223948 336058 224000 336064
rect 222936 335572 222988 335578
rect 222936 335514 222988 335520
rect 222844 334076 222896 334082
rect 222844 334018 222896 334024
rect 222752 320612 222804 320618
rect 222752 320554 222804 320560
rect 221648 319524 221700 319530
rect 221648 319466 221700 319472
rect 221554 51640 221610 51649
rect 221554 51575 221610 51584
rect 221462 50280 221518 50289
rect 221462 50215 221518 50224
rect 221660 49473 221688 319466
rect 221832 318436 221884 318442
rect 221832 318378 221884 318384
rect 221740 286136 221792 286142
rect 221740 286078 221792 286084
rect 221752 56574 221780 286078
rect 221844 213926 221872 318378
rect 222764 227730 222792 320554
rect 222856 295322 222884 334018
rect 222948 299470 222976 335514
rect 223488 319796 223540 319802
rect 223488 319738 223540 319744
rect 223396 318912 223448 318918
rect 223396 318854 223448 318860
rect 223304 318844 223356 318850
rect 223304 318786 223356 318792
rect 223212 314832 223264 314838
rect 223212 314774 223264 314780
rect 222936 299464 222988 299470
rect 222936 299406 222988 299412
rect 223120 298308 223172 298314
rect 223120 298250 223172 298256
rect 223028 297628 223080 297634
rect 223028 297570 223080 297576
rect 222844 295316 222896 295322
rect 222844 295258 222896 295264
rect 222936 294024 222988 294030
rect 222936 293966 222988 293972
rect 222844 286748 222896 286754
rect 222844 286690 222896 286696
rect 222752 227724 222804 227730
rect 222752 227666 222804 227672
rect 221832 213920 221884 213926
rect 221832 213862 221884 213868
rect 222856 57934 222884 286690
rect 222948 95198 222976 293966
rect 223040 109002 223068 297570
rect 223132 115938 223160 298250
rect 223224 194546 223252 314774
rect 223316 218006 223344 318786
rect 223408 219434 223436 318854
rect 223500 220794 223528 319738
rect 223960 303618 223988 336058
rect 224132 331492 224184 331498
rect 224132 331434 224184 331440
rect 224040 323060 224092 323066
rect 224040 323002 224092 323008
rect 223948 303612 224000 303618
rect 223948 303554 224000 303560
rect 224052 283626 224080 323002
rect 224040 283620 224092 283626
rect 224040 283562 224092 283568
rect 224144 278730 224172 331434
rect 224868 329044 224920 329050
rect 224868 328986 224920 328992
rect 224776 325916 224828 325922
rect 224776 325858 224828 325864
rect 224684 324352 224736 324358
rect 224684 324294 224736 324300
rect 224592 323128 224644 323134
rect 224592 323070 224644 323076
rect 224500 312452 224552 312458
rect 224500 312394 224552 312400
rect 224408 309460 224460 309466
rect 224408 309402 224460 309408
rect 224316 305380 224368 305386
rect 224316 305322 224368 305328
rect 224224 302388 224276 302394
rect 224224 302330 224276 302336
rect 224132 278724 224184 278730
rect 224132 278666 224184 278672
rect 223488 220788 223540 220794
rect 223488 220730 223540 220736
rect 223396 219428 223448 219434
rect 223396 219370 223448 219376
rect 223304 218000 223356 218006
rect 223304 217942 223356 217948
rect 223212 194540 223264 194546
rect 223212 194482 223264 194488
rect 224236 135250 224264 302330
rect 224328 147626 224356 305322
rect 224420 168366 224448 309402
rect 224512 184890 224540 312394
rect 224604 241466 224632 323070
rect 224696 245614 224724 324294
rect 224788 252550 224816 325858
rect 224880 266354 224908 328986
rect 226064 327208 226116 327214
rect 226064 327150 226116 327156
rect 225972 324488 226024 324494
rect 225972 324430 226024 324436
rect 225880 316532 225932 316538
rect 225880 316474 225932 316480
rect 225788 311976 225840 311982
rect 225788 311918 225840 311924
rect 225696 308032 225748 308038
rect 225696 307974 225748 307980
rect 225604 294228 225656 294234
rect 225604 294170 225656 294176
rect 224868 266348 224920 266354
rect 224868 266290 224920 266296
rect 224776 252544 224828 252550
rect 224776 252486 224828 252492
rect 224684 245608 224736 245614
rect 224684 245550 224736 245556
rect 224592 241460 224644 241466
rect 224592 241402 224644 241408
rect 224500 184884 224552 184890
rect 224500 184826 224552 184832
rect 224408 168360 224460 168366
rect 224408 168302 224460 168308
rect 224316 147620 224368 147626
rect 224316 147562 224368 147568
rect 224224 135244 224276 135250
rect 224224 135186 224276 135192
rect 224224 119876 224276 119882
rect 224224 119818 224276 119824
rect 223120 115932 223172 115938
rect 223120 115874 223172 115880
rect 223028 108996 223080 109002
rect 223028 108938 223080 108944
rect 222936 95192 222988 95198
rect 222936 95134 222988 95140
rect 224236 91050 224264 119818
rect 225616 96626 225644 294170
rect 225708 164218 225736 307974
rect 225800 180810 225828 311918
rect 225892 205630 225920 316474
rect 225984 248402 226012 324430
rect 226076 260846 226104 327150
rect 226984 319592 227036 319598
rect 226984 319534 227036 319540
rect 226064 260840 226116 260846
rect 226064 260782 226116 260788
rect 225972 248396 226024 248402
rect 225972 248338 226024 248344
rect 225880 205624 225932 205630
rect 225880 205566 225932 205572
rect 225788 180804 225840 180810
rect 225788 180746 225840 180752
rect 225696 164212 225748 164218
rect 225696 164154 225748 164160
rect 225604 96620 225656 96626
rect 225604 96562 225656 96568
rect 224224 91044 224276 91050
rect 224224 90986 224276 90992
rect 224868 77240 224920 77246
rect 224868 77182 224920 77188
rect 224880 73166 224908 77182
rect 224868 73160 224920 73166
rect 224868 73102 224920 73108
rect 222844 57928 222896 57934
rect 222844 57870 222896 57876
rect 221740 56568 221792 56574
rect 221740 56510 221792 56516
rect 223580 50108 223632 50114
rect 223580 50050 223632 50056
rect 221646 49464 221702 49473
rect 221646 49399 221702 49408
rect 220832 16546 221136 16574
rect 220452 9444 220504 9450
rect 220452 9386 220504 9392
rect 218072 6886 218284 6914
rect 217324 3528 217376 3534
rect 217324 3470 217376 3476
rect 218072 480 218100 6886
rect 219256 3664 219308 3670
rect 219256 3606 219308 3612
rect 219268 480 219296 3606
rect 220464 480 220492 9386
rect 195164 354 195192 462
rect 195582 354 195694 480
rect 195164 326 195694 354
rect 195582 -960 195694 326
rect 196778 -960 196890 480
rect 197882 -960 197994 480
rect 199078 -960 199190 480
rect 200274 -960 200386 480
rect 201470 -960 201582 480
rect 202666 -960 202778 480
rect 203862 -960 203974 480
rect 205058 -960 205170 480
rect 206162 -960 206274 480
rect 207358 -960 207470 480
rect 208554 -960 208666 480
rect 209750 -960 209862 480
rect 210946 -960 211058 480
rect 212142 -960 212254 480
rect 213338 -960 213450 480
rect 214442 -960 214554 480
rect 215638 -960 215750 480
rect 216834 -960 216946 480
rect 218030 -960 218142 480
rect 219226 -960 219338 480
rect 220422 -960 220534 480
rect 221108 354 221136 16546
rect 222752 6792 222804 6798
rect 222752 6734 222804 6740
rect 222764 480 222792 6734
rect 221526 354 221638 480
rect 221108 326 221638 354
rect 221526 -960 221638 326
rect 222722 -960 222834 480
rect 223592 354 223620 50050
rect 226996 49337 227024 319534
rect 227088 312594 227116 336874
rect 229836 334620 229888 334626
rect 229836 334562 229888 334568
rect 227720 333124 227772 333130
rect 227720 333066 227772 333072
rect 227536 331628 227588 331634
rect 227536 331570 227588 331576
rect 227352 314900 227404 314906
rect 227352 314842 227404 314848
rect 227076 312588 227128 312594
rect 227076 312530 227128 312536
rect 227260 312248 227312 312254
rect 227260 312190 227312 312196
rect 227168 291372 227220 291378
rect 227168 291314 227220 291320
rect 227076 287428 227128 287434
rect 227076 287370 227128 287376
rect 227088 60722 227116 287370
rect 227180 82822 227208 291314
rect 227272 186318 227300 312190
rect 227364 198694 227392 314842
rect 227444 310684 227496 310690
rect 227444 310626 227496 310632
rect 227456 238066 227484 310626
rect 227548 282878 227576 331570
rect 227732 327758 227760 333066
rect 228916 329996 228968 330002
rect 228916 329938 228968 329944
rect 228824 327956 228876 327962
rect 228824 327898 228876 327904
rect 227720 327752 227772 327758
rect 227720 327694 227772 327700
rect 228732 325780 228784 325786
rect 228732 325722 228784 325728
rect 228640 323332 228692 323338
rect 228640 323274 228692 323280
rect 228364 320952 228416 320958
rect 228364 320894 228416 320900
rect 227536 282872 227588 282878
rect 227536 282814 227588 282820
rect 227444 238060 227496 238066
rect 227444 238002 227496 238008
rect 227352 198688 227404 198694
rect 227352 198630 227404 198636
rect 227260 186312 227312 186318
rect 227260 186254 227312 186260
rect 227168 82816 227220 82822
rect 227168 82758 227220 82764
rect 227076 60716 227128 60722
rect 227076 60658 227128 60664
rect 228376 49570 228404 320894
rect 228548 295520 228600 295526
rect 228548 295462 228600 295468
rect 228456 292732 228508 292738
rect 228456 292674 228508 292680
rect 228468 84182 228496 292674
rect 228560 100706 228588 295462
rect 228652 237386 228680 323274
rect 228744 249762 228772 325722
rect 228836 262206 228864 327898
rect 228928 274650 228956 329938
rect 229744 319660 229796 319666
rect 229744 319602 229796 319608
rect 228916 274644 228968 274650
rect 228916 274586 228968 274592
rect 228824 262200 228876 262206
rect 228824 262142 228876 262148
rect 228732 249756 228784 249762
rect 228732 249698 228784 249704
rect 228640 237380 228692 237386
rect 228640 237322 228692 237328
rect 228548 100700 228600 100706
rect 228548 100642 228600 100648
rect 228456 84176 228508 84182
rect 228456 84118 228508 84124
rect 228364 49564 228416 49570
rect 228364 49506 228416 49512
rect 226982 49328 227038 49337
rect 226982 49263 227038 49272
rect 229756 48793 229784 319602
rect 229848 311846 229876 334562
rect 229928 319728 229980 319734
rect 229928 319670 229980 319676
rect 229836 311840 229888 311846
rect 229836 311782 229888 311788
rect 229836 288584 229888 288590
rect 229836 288526 229888 288532
rect 229848 69018 229876 288526
rect 229836 69012 229888 69018
rect 229836 68954 229888 68960
rect 229940 49609 229968 319670
rect 230204 314764 230256 314770
rect 230204 314706 230256 314712
rect 230112 313472 230164 313478
rect 230112 313414 230164 313420
rect 230020 310616 230072 310622
rect 230020 310558 230072 310564
rect 230032 176662 230060 310558
rect 230124 189038 230152 313414
rect 230216 201482 230244 314706
rect 230204 201476 230256 201482
rect 230204 201418 230256 201424
rect 230112 189032 230164 189038
rect 230112 188974 230164 188980
rect 230020 176656 230072 176662
rect 230020 176598 230072 176604
rect 231136 50930 231164 364346
rect 231228 344962 231256 401610
rect 231412 390522 231440 574058
rect 231492 546508 231544 546514
rect 231492 546450 231544 546456
rect 231400 390516 231452 390522
rect 231400 390458 231452 390464
rect 231504 380798 231532 546450
rect 231584 447160 231636 447166
rect 231584 447102 231636 447108
rect 231492 380792 231544 380798
rect 231492 380734 231544 380740
rect 231596 360058 231624 447102
rect 231676 441652 231728 441658
rect 231676 441594 231728 441600
rect 231584 360052 231636 360058
rect 231584 359994 231636 360000
rect 231688 358766 231716 441594
rect 231768 436144 231820 436150
rect 231768 436086 231820 436092
rect 231676 358760 231728 358766
rect 231676 358702 231728 358708
rect 231780 357406 231808 436086
rect 231768 357400 231820 357406
rect 231768 357342 231820 357348
rect 231216 344956 231268 344962
rect 231216 344898 231268 344904
rect 231676 329928 231728 329934
rect 231676 329870 231728 329876
rect 231584 328568 231636 328574
rect 231584 328510 231636 328516
rect 231492 322992 231544 322998
rect 231492 322934 231544 322940
rect 231400 303816 231452 303822
rect 231400 303758 231452 303764
rect 231308 298240 231360 298246
rect 231308 298182 231360 298188
rect 231216 295452 231268 295458
rect 231216 295394 231268 295400
rect 231228 103494 231256 295394
rect 231320 117298 231348 298182
rect 231412 142118 231440 303758
rect 231504 240106 231532 322934
rect 231596 264926 231624 328510
rect 231688 276010 231716 329870
rect 231676 276004 231728 276010
rect 231676 275946 231728 275952
rect 231584 264920 231636 264926
rect 231584 264862 231636 264868
rect 231492 240100 231544 240106
rect 231492 240042 231544 240048
rect 231400 142112 231452 142118
rect 231400 142054 231452 142060
rect 231308 117292 231360 117298
rect 231308 117234 231360 117240
rect 231216 103488 231268 103494
rect 231216 103430 231268 103436
rect 232516 51513 232544 700266
rect 232596 630692 232648 630698
rect 232596 630634 232648 630640
rect 232608 409834 232636 630634
rect 232688 599004 232740 599010
rect 232688 598946 232740 598952
rect 232596 409828 232648 409834
rect 232596 409770 232648 409776
rect 232700 398682 232728 598946
rect 232780 583772 232832 583778
rect 232780 583714 232832 583720
rect 232688 398676 232740 398682
rect 232688 398618 232740 398624
rect 232792 394534 232820 583714
rect 232872 553444 232924 553450
rect 232872 553386 232924 553392
rect 232780 394528 232832 394534
rect 232780 394470 232832 394476
rect 232884 383654 232912 553386
rect 232964 547936 233016 547942
rect 232964 547878 233016 547884
rect 232872 383648 232924 383654
rect 232872 383590 232924 383596
rect 232976 382090 233004 547878
rect 233056 497480 233108 497486
rect 233056 497422 233108 497428
rect 232964 382084 233016 382090
rect 232964 382026 233016 382032
rect 233068 378010 233096 497422
rect 233056 378004 233108 378010
rect 233056 377946 233108 377952
rect 232688 307964 232740 307970
rect 232688 307906 232740 307912
rect 232596 301096 232648 301102
rect 232596 301038 232648 301044
rect 232608 126954 232636 301038
rect 232700 160070 232728 307906
rect 232872 306536 232924 306542
rect 232872 306478 232924 306484
rect 232780 285796 232832 285802
rect 232780 285738 232832 285744
rect 232792 233918 232820 285738
rect 232884 267034 232912 306478
rect 232872 267028 232924 267034
rect 232872 266970 232924 266976
rect 232780 233912 232832 233918
rect 232780 233854 232832 233860
rect 232688 160064 232740 160070
rect 232688 160006 232740 160012
rect 232596 126948 232648 126954
rect 232596 126890 232648 126896
rect 232502 51504 232558 51513
rect 232502 51439 232558 51448
rect 231124 50924 231176 50930
rect 231124 50866 231176 50872
rect 233896 50425 233924 700470
rect 234160 644564 234212 644570
rect 234160 644506 234212 644512
rect 233976 644496 234028 644502
rect 233976 644438 234028 644444
rect 233988 413914 234016 644438
rect 234068 510672 234120 510678
rect 234068 510614 234120 510620
rect 233976 413908 234028 413914
rect 233976 413850 234028 413856
rect 233976 409896 234028 409902
rect 233976 409838 234028 409844
rect 233988 347682 234016 409838
rect 233976 347676 234028 347682
rect 233976 347618 234028 347624
rect 233976 336864 234028 336870
rect 233976 336806 234028 336812
rect 233988 309806 234016 336806
rect 233976 309800 234028 309806
rect 233976 309742 234028 309748
rect 233976 301028 234028 301034
rect 233976 300970 234028 300976
rect 233988 125594 234016 300970
rect 233976 125588 234028 125594
rect 233976 125530 234028 125536
rect 234080 50561 234108 510614
rect 234172 413846 234200 644506
rect 234252 643136 234304 643142
rect 234252 643078 234304 643084
rect 234264 413982 234292 643078
rect 234344 568676 234396 568682
rect 234344 568618 234396 568624
rect 234252 413976 234304 413982
rect 234252 413918 234304 413924
rect 234160 413840 234212 413846
rect 234160 413782 234212 413788
rect 234160 408536 234212 408542
rect 234160 408478 234212 408484
rect 234172 347750 234200 408478
rect 234356 389094 234384 568618
rect 234436 564460 234488 564466
rect 234436 564402 234488 564408
rect 234344 389088 234396 389094
rect 234344 389030 234396 389036
rect 234448 387666 234476 564402
rect 234528 558952 234580 558958
rect 234528 558894 234580 558900
rect 234436 387660 234488 387666
rect 234436 387602 234488 387608
rect 234540 386238 234568 558894
rect 234528 386232 234580 386238
rect 234528 386174 234580 386180
rect 234252 382288 234304 382294
rect 234252 382230 234304 382236
rect 234160 347744 234212 347750
rect 234160 347686 234212 347692
rect 234264 339318 234292 382230
rect 234252 339312 234304 339318
rect 234252 339254 234304 339260
rect 234344 324964 234396 324970
rect 234344 324906 234396 324912
rect 234252 309256 234304 309262
rect 234252 309198 234304 309204
rect 234160 300960 234212 300966
rect 234160 300902 234212 300908
rect 234172 129742 234200 300902
rect 234264 171086 234292 309198
rect 234356 256698 234384 324906
rect 234344 256692 234396 256698
rect 234344 256634 234396 256640
rect 234252 171080 234304 171086
rect 234252 171022 234304 171028
rect 234160 129736 234212 129742
rect 234160 129678 234212 129684
rect 234066 50552 234122 50561
rect 234066 50487 234122 50496
rect 233882 50416 233938 50425
rect 233882 50351 233938 50360
rect 234632 49638 234660 703582
rect 235000 703474 235028 703582
rect 235142 703520 235254 704960
rect 251426 703520 251538 704960
rect 267618 703520 267730 704960
rect 283810 703520 283922 704960
rect 300094 703520 300206 704960
rect 316286 703520 316398 704960
rect 332478 703520 332590 704960
rect 348762 703520 348874 704960
rect 364954 703520 365066 704960
rect 381146 703520 381258 704960
rect 397430 703520 397542 704960
rect 413622 703520 413734 704960
rect 429814 703520 429926 704960
rect 446098 703520 446210 704960
rect 462290 703520 462402 704960
rect 478482 703520 478594 704960
rect 494766 703520 494878 704960
rect 510958 703520 511070 704960
rect 527150 703520 527262 704960
rect 543434 703520 543546 704960
rect 559626 703520 559738 704960
rect 575818 703520 575930 704960
rect 235184 703474 235212 703520
rect 235000 703446 235212 703474
rect 246396 701004 246448 701010
rect 246396 700946 246448 700952
rect 243636 700868 243688 700874
rect 243636 700810 243688 700816
rect 240784 700800 240836 700806
rect 240784 700742 240836 700748
rect 238024 700120 238076 700126
rect 238024 700062 238076 700068
rect 236644 623892 236696 623898
rect 236644 623834 236696 623840
rect 235264 614168 235316 614174
rect 235264 614110 235316 614116
rect 235276 404190 235304 614110
rect 235356 600364 235408 600370
rect 235356 600306 235408 600312
rect 235264 404184 235316 404190
rect 235264 404126 235316 404132
rect 235368 400042 235396 600306
rect 235448 548004 235500 548010
rect 235448 547946 235500 547952
rect 235356 400036 235408 400042
rect 235356 399978 235408 399984
rect 235460 382158 235488 547946
rect 235540 539640 235592 539646
rect 235540 539582 235592 539588
rect 235448 382152 235500 382158
rect 235448 382094 235500 382100
rect 235552 379370 235580 539582
rect 235632 538280 235684 538286
rect 235632 538222 235684 538228
rect 235540 379364 235592 379370
rect 235540 379306 235592 379312
rect 235644 378078 235672 538222
rect 235724 536852 235776 536858
rect 235724 536794 235776 536800
rect 235736 378146 235764 536794
rect 235816 534132 235868 534138
rect 235816 534074 235868 534080
rect 235828 379438 235856 534074
rect 236656 407046 236684 623834
rect 236736 565888 236788 565894
rect 236736 565830 236788 565836
rect 236644 407040 236696 407046
rect 236644 406982 236696 406988
rect 236644 392012 236696 392018
rect 236644 391954 236696 391960
rect 235816 379432 235868 379438
rect 235816 379374 235868 379380
rect 235724 378140 235776 378146
rect 235724 378082 235776 378088
rect 235632 378072 235684 378078
rect 235632 378014 235684 378020
rect 236656 348430 236684 391954
rect 236748 387734 236776 565830
rect 236828 560312 236880 560318
rect 236828 560254 236880 560260
rect 236736 387728 236788 387734
rect 236736 387670 236788 387676
rect 236840 386306 236868 560254
rect 236920 554804 236972 554810
rect 236920 554746 236972 554752
rect 236828 386300 236880 386306
rect 236828 386242 236880 386248
rect 236932 384878 236960 554746
rect 237012 460216 237064 460222
rect 237012 460158 237064 460164
rect 237024 398750 237052 460158
rect 237012 398744 237064 398750
rect 237012 398686 237064 398692
rect 236920 384872 236972 384878
rect 236920 384814 236972 384820
rect 236644 348424 236696 348430
rect 236644 348366 236696 348372
rect 235632 332716 235684 332722
rect 235632 332658 235684 332664
rect 235540 324420 235592 324426
rect 235540 324362 235592 324368
rect 235448 311908 235500 311914
rect 235448 311850 235500 311856
rect 235356 290012 235408 290018
rect 235356 289954 235408 289960
rect 235264 287156 235316 287162
rect 235264 287098 235316 287104
rect 235276 62082 235304 287098
rect 235368 77246 235396 289954
rect 235460 182170 235488 311850
rect 235552 244254 235580 324362
rect 235644 288386 235672 332658
rect 236920 325712 236972 325718
rect 236920 325654 236972 325660
rect 236828 321768 236880 321774
rect 236828 321710 236880 321716
rect 236644 299600 236696 299606
rect 236644 299542 236696 299548
rect 235632 288380 235684 288386
rect 235632 288322 235684 288328
rect 235540 244248 235592 244254
rect 235540 244190 235592 244196
rect 235448 182164 235500 182170
rect 235448 182106 235500 182112
rect 236656 121446 236684 299542
rect 236736 288516 236788 288522
rect 236736 288458 236788 288464
rect 236748 140078 236776 288458
rect 236840 233238 236868 321710
rect 236932 253910 236960 325654
rect 236920 253904 236972 253910
rect 236920 253846 236972 253852
rect 236828 233232 236880 233238
rect 236828 233174 236880 233180
rect 236736 140072 236788 140078
rect 236736 140014 236788 140020
rect 236644 121440 236696 121446
rect 236644 121382 236696 121388
rect 235356 77240 235408 77246
rect 235356 77182 235408 77188
rect 235264 62076 235316 62082
rect 235264 62018 235316 62024
rect 234712 51876 234764 51882
rect 234712 51818 234764 51824
rect 234620 49632 234672 49638
rect 229926 49600 229982 49609
rect 234620 49574 234672 49580
rect 229926 49535 229982 49544
rect 229742 48784 229798 48793
rect 229742 48719 229798 48728
rect 224224 47456 224276 47462
rect 224224 47398 224276 47404
rect 224236 3670 224264 47398
rect 227720 46368 227772 46374
rect 227720 46310 227772 46316
rect 231858 46336 231914 46345
rect 226340 45008 226392 45014
rect 226340 44950 226392 44956
rect 225144 3936 225196 3942
rect 225144 3878 225196 3884
rect 224224 3664 224276 3670
rect 224224 3606 224276 3612
rect 225156 480 225184 3878
rect 226352 3466 226380 44950
rect 227732 16574 227760 46310
rect 231858 46271 231914 46280
rect 230478 42120 230534 42129
rect 230478 42055 230534 42064
rect 230492 16574 230520 42055
rect 227732 16546 228312 16574
rect 230492 16546 231072 16574
rect 226432 6656 226484 6662
rect 226432 6598 226484 6604
rect 226340 3460 226392 3466
rect 226340 3402 226392 3408
rect 226444 3346 226472 6598
rect 227536 3460 227588 3466
rect 227536 3402 227588 3408
rect 226352 3318 226472 3346
rect 226352 480 226380 3318
rect 227548 480 227576 3402
rect 223918 354 224030 480
rect 223592 326 224030 354
rect 223918 -960 224030 326
rect 225114 -960 225226 480
rect 226310 -960 226422 480
rect 227506 -960 227618 480
rect 228284 354 228312 16546
rect 229836 6452 229888 6458
rect 229836 6394 229888 6400
rect 229848 480 229876 6394
rect 231044 480 231072 16546
rect 228702 354 228814 480
rect 228284 326 228814 354
rect 228702 -960 228814 326
rect 229806 -960 229918 480
rect 231002 -960 231114 480
rect 231872 354 231900 46271
rect 234724 16574 234752 51818
rect 238036 51270 238064 700062
rect 239404 696992 239456 696998
rect 239404 696934 239456 696940
rect 238116 611380 238168 611386
rect 238116 611322 238168 611328
rect 238128 402966 238156 611322
rect 238208 604512 238260 604518
rect 238208 604454 238260 604460
rect 238116 402960 238168 402966
rect 238116 402902 238168 402908
rect 238220 401538 238248 604454
rect 238300 569968 238352 569974
rect 238300 569910 238352 569916
rect 238208 401532 238260 401538
rect 238208 401474 238260 401480
rect 238312 389162 238340 569910
rect 238392 487212 238444 487218
rect 238392 487154 238444 487160
rect 238300 389156 238352 389162
rect 238300 389098 238352 389104
rect 238404 373930 238432 487154
rect 238484 456816 238536 456822
rect 238484 456758 238536 456764
rect 238392 373924 238444 373930
rect 238392 373866 238444 373872
rect 238496 362778 238524 456758
rect 238576 433356 238628 433362
rect 238576 433298 238628 433304
rect 238484 362772 238536 362778
rect 238484 362714 238536 362720
rect 238588 358086 238616 433298
rect 238576 358080 238628 358086
rect 238576 358022 238628 358028
rect 238300 327140 238352 327146
rect 238300 327082 238352 327088
rect 238208 307896 238260 307902
rect 238208 307838 238260 307844
rect 238116 306468 238168 306474
rect 238116 306410 238168 306416
rect 238128 154562 238156 306410
rect 238220 162858 238248 307838
rect 238312 258058 238340 327082
rect 238300 258052 238352 258058
rect 238300 257994 238352 258000
rect 238208 162852 238260 162858
rect 238208 162794 238260 162800
rect 238116 154556 238168 154562
rect 238116 154498 238168 154504
rect 238760 51740 238812 51746
rect 238760 51682 238812 51688
rect 238024 51264 238076 51270
rect 238024 51206 238076 51212
rect 237380 46300 237432 46306
rect 237380 46242 237432 46248
rect 236000 43648 236052 43654
rect 236000 43590 236052 43596
rect 236012 16574 236040 43590
rect 237392 16574 237420 46242
rect 238772 16574 238800 51682
rect 239416 50697 239444 696934
rect 239496 640348 239548 640354
rect 239496 640290 239548 640296
rect 239508 412622 239536 640290
rect 239588 615528 239640 615534
rect 239588 615470 239640 615476
rect 239496 412616 239548 412622
rect 239496 412558 239548 412564
rect 239600 404258 239628 615470
rect 239680 575544 239732 575550
rect 239680 575486 239732 575492
rect 239588 404252 239640 404258
rect 239588 404194 239640 404200
rect 239692 391814 239720 575486
rect 239772 479528 239824 479534
rect 239772 479470 239824 479476
rect 239680 391808 239732 391814
rect 239680 391750 239732 391756
rect 239784 371142 239812 479470
rect 239864 455456 239916 455462
rect 239864 455398 239916 455404
rect 239772 371136 239824 371142
rect 239772 371078 239824 371084
rect 239876 362846 239904 455398
rect 239956 427848 240008 427854
rect 239956 427790 240008 427796
rect 239864 362840 239916 362846
rect 239864 362782 239916 362788
rect 239968 362234 239996 427790
rect 239956 362228 240008 362234
rect 239956 362170 240008 362176
rect 239680 317552 239732 317558
rect 239680 317494 239732 317500
rect 239588 313404 239640 313410
rect 239588 313346 239640 313352
rect 239496 303748 239548 303754
rect 239496 303690 239548 303696
rect 239508 139398 239536 303690
rect 239600 190466 239628 313346
rect 239692 211138 239720 317494
rect 239680 211132 239732 211138
rect 239680 211074 239732 211080
rect 239588 190460 239640 190466
rect 239588 190402 239640 190408
rect 239496 139392 239548 139398
rect 239496 139334 239548 139340
rect 240796 51241 240824 700742
rect 243544 700460 243596 700466
rect 243544 700402 243596 700408
rect 240968 700392 241020 700398
rect 240968 700334 241020 700340
rect 240876 529236 240928 529242
rect 240876 529178 240928 529184
rect 240782 51232 240838 51241
rect 240782 51167 240838 51176
rect 239402 50688 239458 50697
rect 239402 50623 239458 50632
rect 240888 46850 240916 529178
rect 240980 51377 241008 700334
rect 242164 621036 242216 621042
rect 242164 620978 242216 620984
rect 241060 589348 241112 589354
rect 241060 589290 241112 589296
rect 241072 395962 241100 589290
rect 241152 488572 241204 488578
rect 241152 488514 241204 488520
rect 241060 395956 241112 395962
rect 241060 395898 241112 395904
rect 241164 376038 241192 488514
rect 241244 451308 241296 451314
rect 241244 451250 241296 451256
rect 241152 376032 241204 376038
rect 241152 375974 241204 375980
rect 241256 361554 241284 451250
rect 242176 407114 242204 620978
rect 242256 579692 242308 579698
rect 242256 579634 242308 579640
rect 242164 407108 242216 407114
rect 242164 407050 242216 407056
rect 242268 393310 242296 579634
rect 242348 563100 242400 563106
rect 242348 563042 242400 563048
rect 242256 393304 242308 393310
rect 242256 393246 242308 393252
rect 242360 387802 242388 563042
rect 242440 473408 242492 473414
rect 242440 473350 242492 473356
rect 242348 387796 242400 387802
rect 242348 387738 242400 387744
rect 242452 370530 242480 473350
rect 242532 444440 242584 444446
rect 242532 444382 242584 444388
rect 242440 370524 242492 370530
rect 242440 370466 242492 370472
rect 241244 361548 241296 361554
rect 241244 361490 241296 361496
rect 242544 360126 242572 444382
rect 242624 418192 242676 418198
rect 242624 418134 242676 418140
rect 242636 360874 242664 418134
rect 242624 360868 242676 360874
rect 242624 360810 242676 360816
rect 242532 360120 242584 360126
rect 242532 360062 242584 360068
rect 241244 329112 241296 329118
rect 241244 329054 241296 329060
rect 241152 302320 241204 302326
rect 241152 302262 241204 302268
rect 241060 302252 241112 302258
rect 241060 302194 241112 302200
rect 241072 133890 241100 302194
rect 241164 158030 241192 302262
rect 241256 270502 241284 329054
rect 242348 320272 242400 320278
rect 242348 320214 242400 320220
rect 242256 307828 242308 307834
rect 242256 307770 242308 307776
rect 242164 287088 242216 287094
rect 242164 287030 242216 287036
rect 241244 270496 241296 270502
rect 241244 270438 241296 270444
rect 241152 158024 241204 158030
rect 241152 157966 241204 157972
rect 241060 133884 241112 133890
rect 241060 133826 241112 133832
rect 242176 54534 242204 287030
rect 242268 167006 242296 307770
rect 242360 223582 242388 320214
rect 242348 223576 242400 223582
rect 242348 223518 242400 223524
rect 242256 167000 242308 167006
rect 242256 166942 242308 166948
rect 242164 54528 242216 54534
rect 242164 54470 242216 54476
rect 242900 51536 242952 51542
rect 242900 51478 242952 51484
rect 240966 51368 241022 51377
rect 240966 51303 241022 51312
rect 240876 46844 240928 46850
rect 240876 46786 240928 46792
rect 240140 43580 240192 43586
rect 240140 43522 240192 43528
rect 234724 16546 235856 16574
rect 236012 16546 236592 16574
rect 237392 16546 237696 16574
rect 238772 16546 239352 16574
rect 233422 6080 233478 6089
rect 233422 6015 233478 6024
rect 233436 480 233464 6015
rect 234620 3596 234672 3602
rect 234620 3538 234672 3544
rect 234632 480 234660 3538
rect 235828 480 235856 16546
rect 232198 354 232310 480
rect 231872 326 232310 354
rect 232198 -960 232310 326
rect 233394 -960 233506 480
rect 234590 -960 234702 480
rect 235786 -960 235898 480
rect 236564 354 236592 16546
rect 236982 354 237094 480
rect 236564 326 237094 354
rect 237668 354 237696 16546
rect 239324 480 239352 16546
rect 238086 354 238198 480
rect 237668 326 238198 354
rect 236982 -960 237094 326
rect 238086 -960 238198 326
rect 239282 -960 239394 480
rect 240152 354 240180 43522
rect 241704 9376 241756 9382
rect 241704 9318 241756 9324
rect 241716 480 241744 9318
rect 242912 480 242940 51478
rect 243556 48113 243584 700402
rect 243648 48210 243676 700810
rect 246302 700360 246358 700369
rect 246302 700295 246358 700304
rect 244924 634840 244976 634846
rect 244924 634782 244976 634788
rect 243728 592068 243780 592074
rect 243728 592010 243780 592016
rect 243740 397390 243768 592010
rect 243820 561740 243872 561746
rect 243820 561682 243872 561688
rect 243728 397384 243780 397390
rect 243728 397326 243780 397332
rect 243832 386374 243860 561682
rect 243912 492720 243964 492726
rect 243912 492662 243964 492668
rect 243820 386368 243872 386374
rect 243820 386310 243872 386316
rect 243924 375290 243952 492662
rect 244096 463752 244148 463758
rect 244096 463694 244148 463700
rect 244004 462392 244056 462398
rect 244004 462334 244056 462340
rect 243912 375284 243964 375290
rect 243912 375226 243964 375232
rect 244016 365702 244044 462334
rect 244108 369170 244136 463694
rect 244188 416832 244240 416838
rect 244188 416774 244240 416780
rect 244096 369164 244148 369170
rect 244096 369106 244148 369112
rect 244004 365696 244056 365702
rect 244004 365638 244056 365644
rect 244200 350538 244228 416774
rect 244936 411194 244964 634782
rect 245016 625184 245068 625190
rect 245016 625126 245068 625132
rect 244924 411188 244976 411194
rect 244924 411130 244976 411136
rect 245028 408474 245056 625126
rect 245108 585200 245160 585206
rect 245108 585142 245160 585148
rect 245016 408468 245068 408474
rect 245016 408410 245068 408416
rect 245120 394602 245148 585142
rect 245200 557660 245252 557666
rect 245200 557602 245252 557608
rect 245108 394596 245160 394602
rect 245108 394538 245160 394544
rect 245212 384946 245240 557602
rect 245292 469328 245344 469334
rect 245292 469270 245344 469276
rect 245200 384940 245252 384946
rect 245200 384882 245252 384888
rect 245304 366994 245332 469270
rect 246212 437504 246264 437510
rect 246212 437446 246264 437452
rect 245384 429208 245436 429214
rect 245384 429150 245436 429156
rect 245292 366988 245344 366994
rect 245292 366930 245344 366936
rect 245396 354686 245424 429150
rect 245476 426556 245528 426562
rect 245476 426498 245528 426504
rect 245384 354680 245436 354686
rect 245384 354622 245436 354628
rect 245488 353258 245516 426498
rect 245568 414044 245620 414050
rect 245568 413986 245620 413992
rect 245476 353252 245528 353258
rect 245476 353194 245528 353200
rect 244188 350532 244240 350538
rect 244188 350474 244240 350480
rect 245580 349858 245608 413986
rect 246224 359514 246252 437446
rect 246212 359508 246264 359514
rect 246212 359450 246264 359456
rect 245568 349852 245620 349858
rect 245568 349794 245620 349800
rect 244924 332648 244976 332654
rect 244924 332590 244976 332596
rect 243912 314696 243964 314702
rect 243912 314638 243964 314644
rect 243820 305176 243872 305182
rect 243820 305118 243872 305124
rect 243728 292664 243780 292670
rect 243728 292606 243780 292612
rect 243740 86970 243768 292606
rect 243832 146266 243860 305118
rect 243924 197334 243952 314638
rect 244936 305658 244964 332590
rect 245108 310548 245160 310554
rect 245108 310490 245160 310496
rect 244924 305652 244976 305658
rect 244924 305594 244976 305600
rect 245016 305108 245068 305114
rect 245016 305050 245068 305056
rect 244924 289944 244976 289950
rect 244924 289886 244976 289892
rect 243912 197328 243964 197334
rect 243912 197270 243964 197276
rect 243820 146260 243872 146266
rect 243820 146202 243872 146208
rect 243728 86964 243780 86970
rect 243728 86906 243780 86912
rect 244936 74526 244964 289886
rect 245028 150414 245056 305050
rect 245120 178022 245148 310490
rect 245108 178016 245160 178022
rect 245108 177958 245160 177964
rect 245016 150408 245068 150414
rect 245016 150350 245068 150356
rect 244924 74520 244976 74526
rect 244924 74462 244976 74468
rect 246316 48249 246344 700295
rect 246408 50998 246436 700946
rect 246488 700936 246540 700942
rect 246488 700878 246540 700884
rect 246500 51066 246528 700878
rect 253296 700732 253348 700738
rect 253296 700674 253348 700680
rect 249064 700596 249116 700602
rect 249064 700538 249116 700544
rect 246580 612876 246632 612882
rect 246580 612818 246632 612824
rect 246592 404326 246620 612818
rect 247776 597576 247828 597582
rect 247776 597518 247828 597524
rect 246672 590776 246724 590782
rect 246672 590718 246724 590724
rect 246580 404320 246632 404326
rect 246580 404262 246632 404268
rect 246684 396030 246712 590718
rect 246764 556232 246816 556238
rect 246764 556174 246816 556180
rect 246672 396024 246724 396030
rect 246672 395966 246724 395972
rect 246776 385014 246804 556174
rect 247684 529304 247736 529310
rect 247684 529246 247736 529252
rect 246856 485852 246908 485858
rect 246856 485794 246908 485800
rect 246764 385008 246816 385014
rect 246764 384950 246816 384956
rect 246868 373998 246896 485794
rect 246948 436212 247000 436218
rect 246948 436154 247000 436160
rect 246856 373992 246908 373998
rect 246856 373934 246908 373940
rect 246960 356046 246988 436154
rect 246948 356040 247000 356046
rect 246948 355982 247000 355988
rect 246580 335504 246632 335510
rect 246580 335446 246632 335452
rect 246592 300830 246620 335446
rect 246764 309188 246816 309194
rect 246764 309130 246816 309136
rect 246672 305040 246724 305046
rect 246672 304982 246724 304988
rect 246580 300824 246632 300830
rect 246580 300766 246632 300772
rect 246580 296812 246632 296818
rect 246580 296754 246632 296760
rect 246592 107642 246620 296754
rect 246684 151774 246712 304982
rect 246776 172514 246804 309130
rect 246764 172508 246816 172514
rect 246764 172450 246816 172456
rect 246672 151768 246724 151774
rect 246672 151710 246724 151716
rect 246580 107636 246632 107642
rect 246580 107578 246632 107584
rect 246488 51060 246540 51066
rect 246488 51002 246540 51008
rect 246396 50992 246448 50998
rect 246396 50934 246448 50940
rect 246302 48240 246358 48249
rect 243636 48204 243688 48210
rect 246302 48175 246358 48184
rect 243636 48146 243688 48152
rect 243542 48104 243598 48113
rect 243542 48039 243598 48048
rect 244280 48000 244332 48006
rect 244280 47942 244332 47948
rect 242992 43512 243044 43518
rect 242992 43454 243044 43460
rect 243004 16574 243032 43454
rect 244292 16574 244320 47942
rect 247696 46918 247724 529246
rect 247788 398818 247816 597518
rect 247868 594856 247920 594862
rect 247868 594798 247920 594804
rect 247776 398812 247828 398818
rect 247776 398754 247828 398760
rect 247880 397458 247908 594798
rect 247960 549296 248012 549302
rect 247960 549238 248012 549244
rect 247868 397452 247920 397458
rect 247868 397394 247920 397400
rect 247776 396092 247828 396098
rect 247776 396034 247828 396040
rect 247788 343602 247816 396034
rect 247972 382226 248000 549238
rect 248052 458244 248104 458250
rect 248052 458186 248104 458192
rect 247960 382220 248012 382226
rect 247960 382162 248012 382168
rect 248064 364274 248092 458186
rect 248972 423700 249024 423706
rect 248972 423642 249024 423648
rect 248144 412684 248196 412690
rect 248144 412626 248196 412632
rect 248052 364268 248104 364274
rect 248052 364210 248104 364216
rect 248156 349110 248184 412626
rect 248984 356726 249012 423642
rect 248972 356720 249024 356726
rect 248972 356662 249024 356668
rect 248144 349104 248196 349110
rect 248144 349046 248196 349052
rect 247776 343596 247828 343602
rect 247776 343538 247828 343544
rect 247776 336796 247828 336802
rect 247776 336738 247828 336744
rect 247788 309126 247816 336738
rect 248144 331900 248196 331906
rect 248144 331842 248196 331848
rect 248052 316124 248104 316130
rect 248052 316066 248104 316072
rect 247776 309120 247828 309126
rect 247776 309062 247828 309068
rect 247960 306400 248012 306406
rect 247960 306342 248012 306348
rect 247868 296744 247920 296750
rect 247868 296686 247920 296692
rect 247776 289876 247828 289882
rect 247776 289818 247828 289824
rect 247788 70378 247816 289818
rect 247880 111790 247908 296686
rect 247972 155922 248000 306342
rect 248064 202842 248092 316066
rect 248156 291174 248184 331842
rect 248144 291168 248196 291174
rect 248144 291110 248196 291116
rect 248052 202836 248104 202842
rect 248052 202778 248104 202784
rect 247960 155916 248012 155922
rect 247960 155858 248012 155864
rect 247868 111784 247920 111790
rect 247868 111726 247920 111732
rect 247776 70372 247828 70378
rect 247776 70314 247828 70320
rect 249076 50833 249104 700538
rect 253204 700256 253256 700262
rect 253204 700198 253256 700204
rect 251824 700188 251876 700194
rect 251824 700130 251876 700136
rect 251270 645824 251326 645833
rect 251270 645759 251326 645768
rect 251178 644600 251234 644609
rect 251284 644570 251312 645759
rect 251178 644535 251234 644544
rect 251272 644564 251324 644570
rect 251192 644502 251220 644535
rect 251272 644506 251324 644512
rect 251180 644496 251232 644502
rect 251180 644438 251232 644444
rect 251178 643376 251234 643385
rect 251178 643311 251234 643320
rect 251192 643142 251220 643311
rect 251180 643136 251232 643142
rect 251180 643078 251232 643084
rect 251178 642152 251234 642161
rect 251178 642087 251234 642096
rect 251192 641782 251220 642087
rect 251180 641776 251232 641782
rect 251180 641718 251232 641724
rect 251178 640928 251234 640937
rect 251178 640863 251234 640872
rect 251192 640354 251220 640863
rect 251180 640348 251232 640354
rect 251180 640290 251232 640296
rect 251178 639704 251234 639713
rect 251178 639639 251234 639648
rect 251192 638994 251220 639639
rect 251180 638988 251232 638994
rect 251180 638930 251232 638936
rect 251178 638480 251234 638489
rect 251178 638415 251234 638424
rect 251192 637634 251220 638415
rect 251180 637628 251232 637634
rect 251180 637570 251232 637576
rect 250442 637256 250498 637265
rect 250442 637191 250498 637200
rect 249156 601724 249208 601730
rect 249156 601666 249208 601672
rect 249168 400110 249196 601666
rect 249340 579760 249392 579766
rect 249340 579702 249392 579708
rect 249248 529372 249300 529378
rect 249248 529314 249300 529320
rect 249156 400104 249208 400110
rect 249156 400046 249208 400052
rect 249156 387864 249208 387870
rect 249156 387806 249208 387812
rect 249168 340882 249196 387806
rect 249156 340876 249208 340882
rect 249156 340818 249208 340824
rect 249156 291304 249208 291310
rect 249156 291246 249208 291252
rect 249168 80034 249196 291246
rect 249156 80028 249208 80034
rect 249156 79970 249208 79976
rect 249260 50969 249288 529314
rect 249352 391882 249380 579702
rect 249432 577040 249484 577046
rect 249432 576982 249484 576988
rect 249444 391950 249472 576982
rect 249524 541000 249576 541006
rect 249524 540942 249576 540948
rect 249432 391944 249484 391950
rect 249432 391886 249484 391892
rect 249340 391876 249392 391882
rect 249340 391818 249392 391824
rect 249536 379506 249564 540942
rect 249616 478916 249668 478922
rect 249616 478858 249668 478864
rect 249524 379500 249576 379506
rect 249524 379442 249576 379448
rect 249628 371210 249656 478858
rect 249708 465112 249760 465118
rect 249708 465054 249760 465060
rect 249616 371204 249668 371210
rect 249616 371146 249668 371152
rect 249720 367810 249748 465054
rect 250456 411262 250484 637191
rect 251178 636032 251234 636041
rect 251178 635967 251234 635976
rect 251192 634846 251220 635967
rect 251180 634840 251232 634846
rect 251180 634782 251232 634788
rect 251270 634808 251326 634817
rect 251270 634743 251326 634752
rect 251178 633584 251234 633593
rect 251178 633519 251234 633528
rect 251192 632738 251220 633519
rect 251284 633486 251312 634743
rect 251272 633480 251324 633486
rect 251272 633422 251324 633428
rect 251180 632732 251232 632738
rect 251180 632674 251232 632680
rect 251178 632360 251234 632369
rect 251178 632295 251234 632304
rect 251192 632126 251220 632295
rect 251180 632120 251232 632126
rect 251180 632062 251232 632068
rect 251178 631136 251234 631145
rect 251178 631071 251234 631080
rect 251192 630698 251220 631071
rect 251180 630692 251232 630698
rect 251180 630634 251232 630640
rect 251178 629912 251234 629921
rect 251178 629847 251234 629856
rect 251192 629338 251220 629847
rect 251180 629332 251232 629338
rect 251180 629274 251232 629280
rect 251178 628688 251234 628697
rect 251178 628623 251234 628632
rect 251192 627978 251220 628623
rect 251180 627972 251232 627978
rect 251180 627914 251232 627920
rect 251178 627464 251234 627473
rect 251178 627399 251234 627408
rect 251192 626618 251220 627399
rect 251180 626612 251232 626618
rect 251180 626554 251232 626560
rect 251178 626240 251234 626249
rect 251178 626175 251234 626184
rect 251192 625190 251220 626175
rect 251180 625184 251232 625190
rect 251180 625126 251232 625132
rect 251270 625016 251326 625025
rect 251270 624951 251326 624960
rect 251284 623898 251312 624951
rect 251272 623892 251324 623898
rect 251272 623834 251324 623840
rect 251180 623824 251232 623830
rect 251178 623792 251180 623801
rect 251232 623792 251234 623801
rect 251178 623727 251234 623736
rect 251178 622568 251234 622577
rect 251178 622503 251234 622512
rect 251192 622470 251220 622503
rect 251180 622464 251232 622470
rect 251180 622406 251232 622412
rect 251178 621344 251234 621353
rect 251178 621279 251234 621288
rect 251192 621042 251220 621279
rect 251180 621036 251232 621042
rect 251180 620978 251232 620984
rect 251178 620120 251234 620129
rect 251178 620055 251234 620064
rect 251192 619682 251220 620055
rect 251180 619676 251232 619682
rect 251180 619618 251232 619624
rect 251178 618896 251234 618905
rect 251178 618831 251234 618840
rect 251192 618322 251220 618831
rect 251180 618316 251232 618322
rect 251180 618258 251232 618264
rect 251178 617672 251234 617681
rect 251178 617607 251234 617616
rect 251192 616894 251220 617607
rect 251180 616888 251232 616894
rect 251180 616830 251232 616836
rect 251178 616448 251234 616457
rect 251178 616383 251234 616392
rect 251192 615534 251220 616383
rect 251180 615528 251232 615534
rect 251180 615470 251232 615476
rect 251178 615224 251234 615233
rect 251178 615159 251234 615168
rect 251192 614174 251220 615159
rect 251180 614168 251232 614174
rect 251180 614110 251232 614116
rect 251270 614000 251326 614009
rect 251270 613935 251326 613944
rect 251284 612882 251312 613935
rect 251272 612876 251324 612882
rect 251272 612818 251324 612824
rect 251180 612808 251232 612814
rect 251178 612776 251180 612785
rect 251232 612776 251234 612785
rect 251178 612711 251234 612720
rect 251178 611552 251234 611561
rect 251178 611487 251234 611496
rect 251192 611386 251220 611487
rect 251180 611380 251232 611386
rect 251180 611322 251232 611328
rect 251178 610328 251234 610337
rect 251178 610263 251234 610272
rect 251192 610026 251220 610263
rect 251180 610020 251232 610026
rect 251180 609962 251232 609968
rect 251178 609104 251234 609113
rect 251178 609039 251234 609048
rect 251192 608666 251220 609039
rect 251180 608660 251232 608666
rect 251180 608602 251232 608608
rect 251178 607880 251234 607889
rect 251178 607815 251234 607824
rect 251192 607238 251220 607815
rect 251180 607232 251232 607238
rect 251180 607174 251232 607180
rect 250534 606656 250590 606665
rect 250534 606591 250590 606600
rect 250444 411256 250496 411262
rect 250444 411198 250496 411204
rect 250548 401606 250576 606591
rect 251178 605432 251234 605441
rect 251178 605367 251234 605376
rect 251192 604518 251220 605367
rect 251180 604512 251232 604518
rect 251180 604454 251232 604460
rect 251178 604208 251234 604217
rect 251178 604143 251234 604152
rect 251192 603158 251220 604143
rect 251180 603152 251232 603158
rect 251180 603094 251232 603100
rect 251270 601760 251326 601769
rect 251270 601695 251272 601704
rect 251324 601695 251326 601704
rect 251272 601666 251324 601672
rect 251178 600536 251234 600545
rect 251178 600471 251234 600480
rect 251192 600370 251220 600471
rect 251180 600364 251232 600370
rect 251180 600306 251232 600312
rect 251178 599312 251234 599321
rect 251178 599247 251234 599256
rect 251192 599010 251220 599247
rect 251180 599004 251232 599010
rect 251180 598946 251232 598952
rect 251178 598088 251234 598097
rect 251178 598023 251234 598032
rect 251192 597582 251220 598023
rect 251180 597576 251232 597582
rect 251180 597518 251232 597524
rect 251178 595640 251234 595649
rect 251178 595575 251234 595584
rect 251192 594862 251220 595575
rect 251180 594856 251232 594862
rect 251180 594798 251232 594804
rect 251178 594416 251234 594425
rect 251178 594351 251234 594360
rect 251192 593434 251220 594351
rect 251180 593428 251232 593434
rect 251180 593370 251232 593376
rect 251178 593192 251234 593201
rect 251178 593127 251234 593136
rect 251192 592074 251220 593127
rect 251180 592068 251232 592074
rect 251180 592010 251232 592016
rect 251270 591968 251326 591977
rect 251270 591903 251326 591912
rect 251180 590776 251232 590782
rect 251178 590744 251180 590753
rect 251232 590744 251234 590753
rect 251284 590714 251312 591903
rect 251178 590679 251234 590688
rect 251272 590708 251324 590714
rect 251272 590650 251324 590656
rect 251178 589520 251234 589529
rect 251178 589455 251234 589464
rect 251192 589354 251220 589455
rect 251180 589348 251232 589354
rect 251180 589290 251232 589296
rect 251178 588296 251234 588305
rect 251178 588231 251234 588240
rect 251192 587926 251220 588231
rect 251180 587920 251232 587926
rect 251180 587862 251232 587868
rect 250626 587072 250682 587081
rect 250626 587007 250682 587016
rect 250536 401600 250588 401606
rect 250536 401542 250588 401548
rect 250640 394670 250668 587007
rect 251178 585848 251234 585857
rect 251178 585783 251234 585792
rect 251192 585206 251220 585783
rect 251180 585200 251232 585206
rect 251180 585142 251232 585148
rect 251178 584624 251234 584633
rect 251178 584559 251234 584568
rect 251192 583778 251220 584559
rect 251180 583772 251232 583778
rect 251180 583714 251232 583720
rect 251178 583400 251234 583409
rect 251178 583335 251234 583344
rect 251192 582418 251220 583335
rect 251180 582412 251232 582418
rect 251180 582354 251232 582360
rect 251178 582176 251234 582185
rect 251178 582111 251234 582120
rect 251192 581058 251220 582111
rect 251180 581052 251232 581058
rect 251180 580994 251232 581000
rect 251178 580952 251234 580961
rect 251178 580887 251234 580896
rect 251192 579698 251220 580887
rect 251272 579760 251324 579766
rect 251270 579728 251272 579737
rect 251324 579728 251326 579737
rect 251180 579692 251232 579698
rect 251270 579663 251326 579672
rect 251180 579634 251232 579640
rect 251178 578504 251234 578513
rect 251178 578439 251234 578448
rect 251192 578270 251220 578439
rect 251180 578264 251232 578270
rect 251180 578206 251232 578212
rect 251270 577280 251326 577289
rect 251270 577215 251326 577224
rect 251284 577046 251312 577215
rect 251272 577040 251324 577046
rect 251272 576982 251324 576988
rect 251178 576056 251234 576065
rect 251178 575991 251234 576000
rect 251192 575550 251220 575991
rect 251180 575544 251232 575550
rect 251180 575486 251232 575492
rect 251178 574832 251234 574841
rect 251178 574767 251234 574776
rect 251192 574122 251220 574767
rect 251180 574116 251232 574122
rect 251180 574058 251232 574064
rect 251178 573608 251234 573617
rect 251178 573543 251234 573552
rect 251192 572762 251220 573543
rect 251180 572756 251232 572762
rect 251180 572698 251232 572704
rect 251178 572384 251234 572393
rect 251178 572319 251234 572328
rect 251192 571402 251220 572319
rect 251180 571396 251232 571402
rect 251180 571338 251232 571344
rect 251178 571160 251234 571169
rect 251178 571095 251234 571104
rect 251192 569974 251220 571095
rect 251180 569968 251232 569974
rect 251180 569910 251232 569916
rect 251270 569936 251326 569945
rect 251270 569871 251326 569880
rect 251178 568712 251234 568721
rect 251284 568682 251312 569871
rect 251178 568647 251234 568656
rect 251272 568676 251324 568682
rect 251192 568614 251220 568647
rect 251272 568618 251324 568624
rect 251180 568608 251232 568614
rect 251180 568550 251232 568556
rect 251178 567488 251234 567497
rect 251178 567423 251234 567432
rect 251192 567254 251220 567423
rect 251180 567248 251232 567254
rect 251180 567190 251232 567196
rect 251178 566264 251234 566273
rect 251178 566199 251234 566208
rect 251192 565894 251220 566199
rect 251180 565888 251232 565894
rect 251180 565830 251232 565836
rect 251178 565040 251234 565049
rect 251178 564975 251234 564984
rect 251192 564466 251220 564975
rect 251180 564460 251232 564466
rect 251180 564402 251232 564408
rect 251178 563816 251234 563825
rect 251178 563751 251234 563760
rect 251192 563106 251220 563751
rect 251180 563100 251232 563106
rect 251180 563042 251232 563048
rect 251178 562592 251234 562601
rect 251178 562527 251234 562536
rect 251192 561746 251220 562527
rect 251180 561740 251232 561746
rect 251180 561682 251232 561688
rect 251178 561368 251234 561377
rect 251178 561303 251234 561312
rect 251192 560318 251220 561303
rect 251180 560312 251232 560318
rect 251180 560254 251232 560260
rect 251178 560144 251234 560153
rect 251178 560079 251234 560088
rect 251192 558958 251220 560079
rect 251180 558952 251232 558958
rect 251180 558894 251232 558900
rect 251270 558920 251326 558929
rect 251270 558855 251326 558864
rect 251178 557696 251234 557705
rect 251178 557631 251180 557640
rect 251232 557631 251234 557640
rect 251180 557602 251232 557608
rect 251284 557598 251312 558855
rect 251272 557592 251324 557598
rect 251272 557534 251324 557540
rect 251178 556472 251234 556481
rect 251178 556407 251234 556416
rect 251192 556238 251220 556407
rect 251180 556232 251232 556238
rect 251180 556174 251232 556180
rect 251178 555248 251234 555257
rect 251178 555183 251234 555192
rect 251192 554810 251220 555183
rect 251180 554804 251232 554810
rect 251180 554746 251232 554752
rect 251178 554024 251234 554033
rect 251178 553959 251234 553968
rect 251192 553450 251220 553959
rect 251180 553444 251232 553450
rect 251180 553386 251232 553392
rect 251178 552800 251234 552809
rect 251178 552735 251234 552744
rect 251192 552090 251220 552735
rect 251180 552084 251232 552090
rect 251180 552026 251232 552032
rect 251178 551576 251234 551585
rect 251178 551511 251234 551520
rect 251192 550662 251220 551511
rect 251180 550656 251232 550662
rect 251180 550598 251232 550604
rect 251178 550352 251234 550361
rect 251178 550287 251234 550296
rect 251192 549302 251220 550287
rect 251180 549296 251232 549302
rect 251180 549238 251232 549244
rect 251270 549128 251326 549137
rect 251270 549063 251326 549072
rect 251284 548010 251312 549063
rect 251272 548004 251324 548010
rect 251272 547946 251324 547952
rect 251180 547936 251232 547942
rect 251178 547904 251180 547913
rect 251232 547904 251234 547913
rect 251178 547839 251234 547848
rect 251178 546680 251234 546689
rect 251178 546615 251234 546624
rect 251192 546514 251220 546615
rect 251180 546508 251232 546514
rect 251180 546450 251232 546456
rect 251178 545456 251234 545465
rect 251178 545391 251234 545400
rect 251192 545154 251220 545391
rect 251180 545148 251232 545154
rect 251180 545090 251232 545096
rect 251178 544232 251234 544241
rect 251178 544167 251234 544176
rect 251192 543794 251220 544167
rect 251180 543788 251232 543794
rect 251180 543730 251232 543736
rect 250718 543008 250774 543017
rect 250718 542943 250774 542952
rect 250628 394664 250680 394670
rect 250628 394606 250680 394612
rect 250444 393916 250496 393922
rect 250444 393858 250496 393864
rect 249708 367804 249760 367810
rect 249708 367746 249760 367752
rect 250456 345030 250484 393858
rect 250732 380866 250760 542943
rect 251178 541784 251234 541793
rect 251178 541719 251234 541728
rect 251192 541006 251220 541719
rect 251180 541000 251232 541006
rect 251180 540942 251232 540948
rect 251178 540560 251234 540569
rect 251178 540495 251234 540504
rect 251192 539646 251220 540495
rect 251180 539640 251232 539646
rect 251180 539582 251232 539588
rect 251178 539336 251234 539345
rect 251178 539271 251234 539280
rect 251192 538286 251220 539271
rect 251180 538280 251232 538286
rect 251180 538222 251232 538228
rect 251178 538112 251234 538121
rect 251178 538047 251234 538056
rect 251192 536858 251220 538047
rect 251180 536852 251232 536858
rect 251180 536794 251232 536800
rect 251178 535664 251234 535673
rect 251178 535599 251234 535608
rect 251192 535498 251220 535599
rect 251180 535492 251232 535498
rect 251180 535434 251232 535440
rect 251178 534440 251234 534449
rect 251178 534375 251234 534384
rect 251192 534138 251220 534375
rect 251180 534132 251232 534138
rect 251180 534074 251232 534080
rect 251178 496224 251234 496233
rect 251178 496159 251234 496168
rect 251192 495514 251220 496159
rect 251180 495508 251232 495514
rect 251180 495450 251232 495456
rect 251178 495000 251234 495009
rect 251178 494935 251234 494944
rect 251192 494086 251220 494935
rect 251180 494080 251232 494086
rect 251180 494022 251232 494028
rect 251178 493776 251234 493785
rect 251178 493711 251234 493720
rect 251192 492726 251220 493711
rect 251180 492720 251232 492726
rect 251180 492662 251232 492668
rect 251178 492552 251234 492561
rect 251178 492487 251234 492496
rect 251192 491366 251220 492487
rect 251180 491360 251232 491366
rect 250810 491328 250866 491337
rect 251180 491302 251232 491308
rect 250810 491263 250866 491272
rect 250720 380860 250772 380866
rect 250720 380802 250772 380808
rect 250824 375358 250852 491263
rect 251178 490104 251234 490113
rect 251178 490039 251234 490048
rect 251192 489938 251220 490039
rect 251180 489932 251232 489938
rect 251180 489874 251232 489880
rect 251178 488880 251234 488889
rect 251178 488815 251234 488824
rect 251192 488578 251220 488815
rect 251180 488572 251232 488578
rect 251180 488514 251232 488520
rect 251178 487656 251234 487665
rect 251178 487591 251234 487600
rect 251192 487218 251220 487591
rect 251180 487212 251232 487218
rect 251180 487154 251232 487160
rect 251178 486432 251234 486441
rect 251178 486367 251234 486376
rect 251192 485858 251220 486367
rect 251180 485852 251232 485858
rect 251180 485794 251232 485800
rect 251178 485208 251234 485217
rect 251178 485143 251234 485152
rect 251192 484430 251220 485143
rect 251180 484424 251232 484430
rect 251180 484366 251232 484372
rect 251178 483984 251234 483993
rect 251178 483919 251234 483928
rect 251192 483070 251220 483919
rect 251180 483064 251232 483070
rect 251180 483006 251232 483012
rect 251178 482760 251234 482769
rect 251178 482695 251234 482704
rect 251192 481710 251220 482695
rect 251180 481704 251232 481710
rect 251180 481646 251232 481652
rect 251178 481536 251234 481545
rect 251178 481471 251234 481480
rect 251192 480282 251220 481471
rect 251180 480276 251232 480282
rect 251180 480218 251232 480224
rect 251178 479088 251234 479097
rect 251178 479023 251234 479032
rect 251192 478922 251220 479023
rect 251180 478916 251232 478922
rect 251180 478858 251232 478864
rect 251178 477864 251234 477873
rect 251178 477799 251234 477808
rect 251192 477562 251220 477799
rect 251180 477556 251232 477562
rect 251180 477498 251232 477504
rect 251178 476640 251234 476649
rect 251178 476575 251234 476584
rect 251192 476134 251220 476575
rect 251180 476128 251232 476134
rect 251180 476070 251232 476076
rect 251178 475416 251234 475425
rect 251178 475351 251234 475360
rect 251192 474774 251220 475351
rect 251180 474768 251232 474774
rect 251180 474710 251232 474716
rect 251178 474192 251234 474201
rect 251178 474127 251234 474136
rect 251192 473414 251220 474127
rect 251180 473408 251232 473414
rect 251180 473350 251232 473356
rect 251178 472968 251234 472977
rect 251178 472903 251234 472912
rect 251192 472054 251220 472903
rect 251180 472048 251232 472054
rect 251180 471990 251232 471996
rect 251178 471744 251234 471753
rect 251178 471679 251234 471688
rect 251192 470626 251220 471679
rect 251180 470620 251232 470626
rect 251180 470562 251232 470568
rect 251270 470520 251326 470529
rect 251270 470455 251326 470464
rect 251180 469328 251232 469334
rect 251178 469296 251180 469305
rect 251232 469296 251234 469305
rect 251284 469266 251312 470455
rect 251178 469231 251234 469240
rect 251272 469260 251324 469266
rect 251272 469202 251324 469208
rect 251178 466848 251234 466857
rect 251178 466783 251234 466792
rect 251192 466478 251220 466783
rect 251180 466472 251232 466478
rect 251180 466414 251232 466420
rect 251638 465624 251694 465633
rect 251638 465559 251694 465568
rect 251652 465118 251680 465559
rect 251640 465112 251692 465118
rect 251640 465054 251692 465060
rect 251178 464400 251234 464409
rect 251178 464335 251234 464344
rect 251192 463758 251220 464335
rect 251180 463752 251232 463758
rect 251180 463694 251232 463700
rect 251178 463176 251234 463185
rect 251178 463111 251234 463120
rect 251192 462398 251220 463111
rect 251180 462392 251232 462398
rect 251180 462334 251232 462340
rect 251178 460728 251234 460737
rect 251178 460663 251234 460672
rect 251192 459610 251220 460663
rect 251180 459604 251232 459610
rect 251180 459546 251232 459552
rect 251178 459504 251234 459513
rect 251178 459439 251234 459448
rect 251192 458250 251220 459439
rect 251180 458244 251232 458250
rect 251180 458186 251232 458192
rect 251178 457056 251234 457065
rect 251178 456991 251234 457000
rect 251192 456822 251220 456991
rect 251180 456816 251232 456822
rect 251180 456758 251232 456764
rect 251178 455832 251234 455841
rect 251178 455767 251234 455776
rect 251192 455462 251220 455767
rect 251180 455456 251232 455462
rect 251180 455398 251232 455404
rect 251178 454608 251234 454617
rect 251178 454543 251234 454552
rect 251192 454102 251220 454543
rect 251180 454096 251232 454102
rect 251180 454038 251232 454044
rect 251730 453384 251786 453393
rect 251730 453319 251786 453328
rect 251178 452160 251234 452169
rect 251178 452095 251234 452104
rect 251192 451314 251220 452095
rect 251180 451308 251232 451314
rect 251180 451250 251232 451256
rect 251178 450936 251234 450945
rect 251178 450871 251234 450880
rect 251192 449954 251220 450871
rect 251180 449948 251232 449954
rect 251180 449890 251232 449896
rect 251178 449712 251234 449721
rect 251178 449647 251234 449656
rect 251192 448594 251220 449647
rect 251180 448588 251232 448594
rect 251180 448530 251232 448536
rect 251178 447264 251234 447273
rect 251178 447199 251234 447208
rect 251192 447166 251220 447199
rect 251180 447160 251232 447166
rect 251180 447102 251232 447108
rect 251744 446486 251772 453319
rect 251732 446480 251784 446486
rect 251732 446422 251784 446428
rect 251732 446344 251784 446350
rect 251732 446286 251784 446292
rect 251178 446040 251234 446049
rect 251178 445975 251234 445984
rect 251192 445806 251220 445975
rect 251180 445800 251232 445806
rect 251180 445742 251232 445748
rect 251178 444816 251234 444825
rect 251178 444751 251234 444760
rect 251192 444446 251220 444751
rect 251180 444440 251232 444446
rect 251180 444382 251232 444388
rect 250902 443592 250958 443601
rect 250902 443527 250958 443536
rect 250812 375352 250864 375358
rect 250812 375294 250864 375300
rect 250916 366382 250944 443527
rect 251178 442368 251234 442377
rect 251178 442303 251234 442312
rect 251192 441658 251220 442303
rect 251180 441652 251232 441658
rect 251180 441594 251232 441600
rect 251178 441144 251234 441153
rect 251178 441079 251234 441088
rect 251192 440298 251220 441079
rect 251180 440292 251232 440298
rect 251180 440234 251232 440240
rect 251178 439920 251234 439929
rect 251178 439855 251234 439864
rect 251192 438938 251220 439855
rect 251744 439550 251772 446286
rect 251732 439544 251784 439550
rect 251732 439486 251784 439492
rect 251180 438932 251232 438938
rect 251180 438874 251232 438880
rect 251178 438696 251234 438705
rect 251178 438631 251234 438640
rect 251192 437510 251220 438631
rect 251180 437504 251232 437510
rect 251180 437446 251232 437452
rect 251270 437472 251326 437481
rect 251270 437407 251326 437416
rect 251178 436248 251234 436257
rect 251178 436183 251180 436192
rect 251232 436183 251234 436192
rect 251180 436154 251232 436160
rect 251284 436150 251312 437407
rect 251272 436144 251324 436150
rect 251272 436086 251324 436092
rect 251178 435024 251234 435033
rect 251178 434959 251234 434968
rect 251192 434790 251220 434959
rect 251180 434784 251232 434790
rect 251180 434726 251232 434732
rect 251178 433800 251234 433809
rect 251178 433735 251234 433744
rect 251192 433362 251220 433735
rect 251180 433356 251232 433362
rect 251180 433298 251232 433304
rect 251178 432576 251234 432585
rect 251178 432511 251234 432520
rect 251192 432002 251220 432511
rect 251180 431996 251232 432002
rect 251180 431938 251232 431944
rect 251178 431352 251234 431361
rect 251178 431287 251234 431296
rect 251192 430642 251220 431287
rect 251180 430636 251232 430642
rect 251180 430578 251232 430584
rect 251178 430128 251234 430137
rect 251178 430063 251234 430072
rect 251192 429214 251220 430063
rect 251180 429208 251232 429214
rect 251180 429150 251232 429156
rect 251178 428904 251234 428913
rect 251178 428839 251234 428848
rect 251192 427854 251220 428839
rect 251180 427848 251232 427854
rect 251180 427790 251232 427796
rect 251270 427680 251326 427689
rect 251270 427615 251326 427624
rect 251284 426562 251312 427615
rect 251272 426556 251324 426562
rect 251272 426498 251324 426504
rect 251180 426488 251232 426494
rect 251178 426456 251180 426465
rect 251232 426456 251234 426465
rect 251178 426391 251234 426400
rect 251178 425232 251234 425241
rect 251178 425167 251234 425176
rect 251192 425134 251220 425167
rect 251180 425128 251232 425134
rect 251180 425070 251232 425076
rect 251178 424008 251234 424017
rect 251178 423943 251234 423952
rect 251192 423706 251220 423943
rect 251180 423700 251232 423706
rect 251180 423642 251232 423648
rect 250994 422784 251050 422793
rect 250994 422719 251050 422728
rect 250904 366376 250956 366382
rect 250904 366318 250956 366324
rect 251008 351898 251036 422719
rect 251178 421560 251234 421569
rect 251178 421495 251234 421504
rect 251192 420986 251220 421495
rect 251180 420980 251232 420986
rect 251180 420922 251232 420928
rect 251178 420336 251234 420345
rect 251178 420271 251234 420280
rect 251192 419558 251220 420271
rect 251180 419552 251232 419558
rect 251180 419494 251232 419500
rect 251178 419112 251234 419121
rect 251178 419047 251234 419056
rect 251192 418198 251220 419047
rect 251180 418192 251232 418198
rect 251180 418134 251232 418140
rect 251178 417888 251234 417897
rect 251178 417823 251234 417832
rect 251192 416838 251220 417823
rect 251180 416832 251232 416838
rect 251180 416774 251232 416780
rect 251270 416664 251326 416673
rect 251270 416599 251326 416608
rect 251284 415546 251312 416599
rect 251272 415540 251324 415546
rect 251272 415482 251324 415488
rect 251180 415472 251232 415478
rect 251178 415440 251180 415449
rect 251232 415440 251234 415449
rect 251178 415375 251234 415384
rect 251178 414216 251234 414225
rect 251178 414151 251234 414160
rect 251192 414050 251220 414151
rect 251180 414044 251232 414050
rect 251180 413986 251232 413992
rect 251178 412992 251234 413001
rect 251178 412927 251234 412936
rect 251192 412690 251220 412927
rect 251180 412684 251232 412690
rect 251180 412626 251232 412632
rect 251178 411768 251234 411777
rect 251178 411703 251234 411712
rect 251192 411330 251220 411703
rect 251180 411324 251232 411330
rect 251180 411266 251232 411272
rect 251178 410544 251234 410553
rect 251178 410479 251234 410488
rect 251192 409902 251220 410479
rect 251180 409896 251232 409902
rect 251180 409838 251232 409844
rect 251178 409320 251234 409329
rect 251178 409255 251234 409264
rect 251192 408542 251220 409255
rect 251180 408536 251232 408542
rect 251180 408478 251232 408484
rect 251178 408096 251234 408105
rect 251178 408031 251234 408040
rect 251192 407182 251220 408031
rect 251180 407176 251232 407182
rect 251180 407118 251232 407124
rect 251638 406872 251694 406881
rect 251638 406807 251694 406816
rect 251178 405648 251234 405657
rect 251178 405583 251234 405592
rect 251192 404394 251220 405583
rect 251180 404388 251232 404394
rect 251180 404330 251232 404336
rect 251086 403200 251142 403209
rect 251086 403135 251142 403144
rect 251100 354006 251128 403135
rect 251178 401976 251234 401985
rect 251178 401911 251234 401920
rect 251192 401674 251220 401911
rect 251180 401668 251232 401674
rect 251180 401610 251232 401616
rect 251652 400926 251680 406807
rect 251730 404424 251786 404433
rect 251730 404359 251786 404368
rect 251640 400920 251692 400926
rect 251640 400862 251692 400868
rect 251548 400852 251600 400858
rect 251548 400794 251600 400800
rect 251560 400178 251588 400794
rect 251548 400172 251600 400178
rect 251548 400114 251600 400120
rect 251178 399528 251234 399537
rect 251178 399463 251234 399472
rect 251192 398886 251220 399463
rect 251180 398880 251232 398886
rect 251180 398822 251232 398828
rect 251178 398304 251234 398313
rect 251178 398239 251234 398248
rect 251192 397526 251220 398239
rect 251744 398138 251772 404359
rect 251732 398132 251784 398138
rect 251732 398074 251784 398080
rect 251180 397520 251232 397526
rect 251180 397462 251232 397468
rect 251178 397080 251234 397089
rect 251178 397015 251234 397024
rect 251192 396098 251220 397015
rect 251180 396092 251232 396098
rect 251180 396034 251232 396040
rect 251178 395856 251234 395865
rect 251178 395791 251234 395800
rect 251192 394738 251220 395791
rect 251180 394732 251232 394738
rect 251180 394674 251232 394680
rect 251638 394632 251694 394641
rect 251638 394567 251694 394576
rect 251178 393408 251234 393417
rect 251178 393343 251180 393352
rect 251232 393343 251234 393352
rect 251180 393314 251232 393320
rect 251178 392184 251234 392193
rect 251178 392119 251234 392128
rect 251192 392018 251220 392119
rect 251180 392012 251232 392018
rect 251180 391954 251232 391960
rect 251178 390960 251234 390969
rect 251178 390895 251234 390904
rect 251192 390590 251220 390895
rect 251180 390584 251232 390590
rect 251180 390526 251232 390532
rect 251178 389736 251234 389745
rect 251178 389671 251234 389680
rect 251192 389230 251220 389671
rect 251180 389224 251232 389230
rect 251180 389166 251232 389172
rect 251454 388512 251510 388521
rect 251652 388482 251680 394567
rect 251454 388447 251510 388456
rect 251640 388476 251692 388482
rect 251468 387870 251496 388447
rect 251640 388418 251692 388424
rect 251456 387864 251508 387870
rect 251456 387806 251508 387812
rect 251730 387288 251786 387297
rect 251730 387223 251786 387232
rect 251454 386064 251510 386073
rect 251454 385999 251510 386008
rect 251178 384840 251234 384849
rect 251178 384775 251234 384784
rect 251192 383722 251220 384775
rect 251180 383716 251232 383722
rect 251180 383658 251232 383664
rect 251468 383654 251496 385999
rect 251468 383626 251680 383654
rect 251178 383616 251234 383625
rect 251178 383551 251234 383560
rect 251192 382294 251220 383551
rect 251180 382288 251232 382294
rect 251180 382230 251232 382236
rect 251088 354000 251140 354006
rect 251088 353942 251140 353948
rect 250996 351892 251048 351898
rect 250996 351834 251048 351840
rect 250444 345024 250496 345030
rect 250444 344966 250496 344972
rect 251652 339386 251680 383626
rect 251744 339454 251772 387223
rect 251732 339448 251784 339454
rect 251732 339390 251784 339396
rect 251640 339380 251692 339386
rect 251640 339322 251692 339328
rect 249616 334008 249668 334014
rect 249616 333950 249668 333956
rect 249524 320204 249576 320210
rect 249524 320146 249576 320152
rect 249432 313336 249484 313342
rect 249432 313278 249484 313284
rect 249340 292596 249392 292602
rect 249340 292538 249392 292544
rect 249352 88330 249380 292538
rect 249444 193186 249472 313278
rect 249536 224942 249564 320146
rect 249628 292534 249656 333950
rect 250444 329860 250496 329866
rect 250444 329802 250496 329808
rect 250456 292806 250484 329802
rect 250720 321700 250772 321706
rect 250720 321642 250772 321648
rect 250628 303680 250680 303686
rect 250628 303622 250680 303628
rect 250444 292800 250496 292806
rect 250444 292742 250496 292748
rect 249616 292528 249668 292534
rect 249616 292470 249668 292476
rect 250536 291236 250588 291242
rect 250536 291178 250588 291184
rect 250444 288448 250496 288454
rect 250444 288390 250496 288396
rect 249524 224936 249576 224942
rect 249524 224878 249576 224884
rect 249432 193180 249484 193186
rect 249432 193122 249484 193128
rect 249340 88324 249392 88330
rect 249340 88266 249392 88272
rect 250456 64462 250484 288390
rect 250548 78674 250576 291178
rect 250640 143546 250668 303622
rect 250732 229022 250760 321642
rect 250720 229016 250772 229022
rect 250720 228958 250772 228964
rect 250628 143540 250680 143546
rect 250628 143482 250680 143488
rect 250536 78668 250588 78674
rect 250536 78610 250588 78616
rect 250444 64456 250496 64462
rect 250444 64398 250496 64404
rect 249246 50960 249302 50969
rect 249246 50895 249302 50904
rect 249062 50824 249118 50833
rect 249062 50759 249118 50768
rect 251836 48278 251864 700130
rect 251914 602984 251970 602993
rect 251914 602919 251970 602928
rect 251928 400858 251956 602919
rect 252098 596864 252154 596873
rect 252098 596799 252154 596808
rect 252006 533216 252062 533225
rect 252006 533151 252062 533160
rect 251916 400852 251968 400858
rect 251916 400794 251968 400800
rect 251914 400752 251970 400761
rect 251914 400687 251970 400696
rect 251928 393922 251956 400687
rect 251916 393916 251968 393922
rect 251916 393858 251968 393864
rect 251916 388476 251968 388482
rect 251916 388418 251968 388424
rect 251928 342174 251956 388418
rect 252020 376718 252048 533151
rect 252112 460222 252140 596799
rect 252190 536888 252246 536897
rect 252190 536823 252246 536832
rect 252204 497486 252232 536823
rect 252192 497480 252244 497486
rect 252192 497422 252244 497428
rect 252374 480312 252430 480321
rect 252374 480247 252430 480256
rect 252388 479534 252416 480247
rect 252376 479528 252428 479534
rect 252376 479470 252428 479476
rect 252190 468072 252246 468081
rect 252190 468007 252246 468016
rect 252100 460216 252152 460222
rect 252100 460158 252152 460164
rect 252098 458280 252154 458289
rect 252098 458215 252154 458224
rect 252008 376712 252060 376718
rect 252008 376654 252060 376660
rect 252112 364342 252140 458215
rect 252204 367062 252232 468007
rect 252466 461952 252522 461961
rect 252466 461887 252522 461896
rect 252374 448488 252430 448497
rect 252374 448423 252430 448432
rect 252284 446480 252336 446486
rect 252284 446422 252336 446428
rect 252192 367056 252244 367062
rect 252192 366998 252244 367004
rect 252100 364336 252152 364342
rect 252100 364278 252152 364284
rect 252296 362710 252324 446422
rect 252284 362704 252336 362710
rect 252284 362646 252336 362652
rect 252388 360194 252416 448423
rect 252480 446350 252508 461887
rect 252468 446344 252520 446350
rect 252468 446286 252520 446292
rect 252468 398132 252520 398138
rect 252468 398074 252520 398080
rect 252376 360188 252428 360194
rect 252376 360130 252428 360136
rect 252480 346390 252508 398074
rect 252468 346384 252520 346390
rect 252468 346326 252520 346332
rect 251916 342168 251968 342174
rect 251916 342110 251968 342116
rect 252008 319048 252060 319054
rect 252008 318990 252060 318996
rect 251916 299532 251968 299538
rect 251916 299474 251968 299480
rect 251928 120086 251956 299474
rect 252020 215286 252048 318990
rect 252008 215280 252060 215286
rect 252008 215222 252060 215228
rect 251916 120080 251968 120086
rect 251916 120022 251968 120028
rect 253216 51202 253244 700198
rect 253204 51196 253256 51202
rect 253204 51138 253256 51144
rect 253308 51105 253336 700674
rect 267660 700126 267688 703520
rect 283852 700194 283880 703520
rect 300136 700262 300164 703520
rect 332520 701010 332548 703520
rect 332508 701004 332560 701010
rect 332508 700946 332560 700952
rect 348804 700942 348832 703520
rect 348792 700936 348844 700942
rect 348792 700878 348844 700884
rect 364996 700874 365024 703520
rect 364984 700868 365036 700874
rect 364984 700810 365036 700816
rect 397472 700806 397500 703520
rect 397460 700800 397512 700806
rect 397460 700742 397512 700748
rect 413664 700670 413692 703520
rect 429856 700738 429884 703520
rect 429844 700732 429896 700738
rect 429844 700674 429896 700680
rect 413652 700664 413704 700670
rect 413652 700606 413704 700612
rect 462332 700602 462360 703520
rect 462320 700596 462372 700602
rect 462320 700538 462372 700544
rect 478524 700534 478552 703520
rect 478512 700528 478564 700534
rect 478512 700470 478564 700476
rect 494808 700466 494836 703520
rect 494796 700460 494848 700466
rect 494796 700402 494848 700408
rect 527192 700398 527220 703520
rect 527180 700392 527232 700398
rect 527180 700334 527232 700340
rect 543476 700330 543504 703520
rect 559668 700369 559696 703520
rect 559654 700360 559710 700369
rect 543464 700324 543516 700330
rect 559654 700295 559710 700304
rect 543464 700266 543516 700272
rect 300124 700256 300176 700262
rect 300124 700198 300176 700204
rect 283840 700188 283892 700194
rect 283840 700130 283892 700136
rect 267648 700120 267700 700126
rect 267648 700062 267700 700068
rect 580170 697232 580226 697241
rect 580170 697167 580226 697176
rect 580184 696998 580212 697167
rect 580172 696992 580224 696998
rect 580172 696934 580224 696940
rect 580170 683904 580226 683913
rect 580170 683839 580226 683848
rect 580184 683194 580212 683839
rect 580172 683188 580224 683194
rect 580172 683130 580224 683136
rect 580538 644056 580594 644065
rect 580538 643991 580594 644000
rect 580262 630864 580318 630873
rect 580262 630799 580318 630808
rect 580170 617536 580226 617545
rect 580170 617471 580226 617480
rect 580184 616894 580212 617471
rect 574744 616888 574796 616894
rect 574744 616830 574796 616836
rect 580172 616888 580224 616894
rect 580172 616830 580224 616836
rect 573364 456816 573416 456822
rect 573364 456758 573416 456764
rect 258724 351960 258776 351966
rect 258724 351902 258776 351908
rect 254952 331288 255004 331294
rect 254952 331230 255004 331236
rect 254584 318844 254636 318850
rect 254584 318786 254636 318792
rect 253388 52488 253440 52494
rect 253388 52430 253440 52436
rect 253294 51096 253350 51105
rect 253294 51031 253350 51040
rect 253204 50652 253256 50658
rect 253204 50594 253256 50600
rect 252560 50380 252612 50386
rect 252560 50322 252612 50328
rect 251824 48272 251876 48278
rect 251824 48214 251876 48220
rect 248420 47932 248472 47938
rect 248420 47874 248472 47880
rect 247684 46912 247736 46918
rect 247684 46854 247736 46860
rect 247038 43480 247094 43489
rect 247038 43415 247094 43424
rect 247052 16574 247080 43415
rect 243004 16546 244136 16574
rect 244292 16546 245240 16574
rect 247052 16546 247632 16574
rect 244108 480 244136 16546
rect 245212 480 245240 16546
rect 246396 3732 246448 3738
rect 246396 3674 246448 3680
rect 246408 480 246436 3674
rect 247604 480 247632 16546
rect 240478 354 240590 480
rect 240152 326 240590 354
rect 240478 -960 240590 326
rect 241674 -960 241786 480
rect 242870 -960 242982 480
rect 244066 -960 244178 480
rect 245170 -960 245282 480
rect 246366 -960 246478 480
rect 247562 -960 247674 480
rect 248432 354 248460 47874
rect 251180 47864 251232 47870
rect 251180 47806 251232 47812
rect 249800 44940 249852 44946
rect 249800 44882 249852 44888
rect 249812 16574 249840 44882
rect 249812 16546 250024 16574
rect 249996 480 250024 16546
rect 251192 3466 251220 47806
rect 252572 6914 252600 50322
rect 253216 9382 253244 50594
rect 253296 50516 253348 50522
rect 253296 50458 253348 50464
rect 253204 9376 253256 9382
rect 253204 9318 253256 9324
rect 253308 8906 253336 50458
rect 253296 8900 253348 8906
rect 253296 8842 253348 8848
rect 251270 6896 251326 6905
rect 252572 6886 253336 6914
rect 251270 6831 251326 6840
rect 251180 3460 251232 3466
rect 251180 3402 251232 3408
rect 251284 3346 251312 6831
rect 253308 3482 253336 6886
rect 253400 6050 253428 52430
rect 253572 51808 253624 51814
rect 253572 51750 253624 51756
rect 253480 51672 253532 51678
rect 253480 51614 253532 51620
rect 253492 9586 253520 51614
rect 253480 9580 253532 9586
rect 253480 9522 253532 9528
rect 253584 9450 253612 51750
rect 254596 48618 254624 318786
rect 254860 316056 254912 316062
rect 254860 315998 254912 316004
rect 254768 298172 254820 298178
rect 254768 298114 254820 298120
rect 254676 294160 254728 294166
rect 254676 294102 254728 294108
rect 254688 92478 254716 294102
rect 254780 112946 254808 298114
rect 254872 206990 254900 315998
rect 254964 280158 254992 331230
rect 255964 328500 256016 328506
rect 255964 328442 256016 328448
rect 255976 289814 256004 328442
rect 257344 327752 257396 327758
rect 257344 327694 257396 327700
rect 256332 321632 256384 321638
rect 256332 321574 256384 321580
rect 256240 317484 256292 317490
rect 256240 317426 256292 317432
rect 256148 300892 256200 300898
rect 256148 300834 256200 300840
rect 256056 295384 256108 295390
rect 256056 295326 256108 295332
rect 255964 289808 256016 289814
rect 255964 289750 256016 289756
rect 255964 285932 256016 285938
rect 255964 285874 256016 285880
rect 254952 280152 255004 280158
rect 254952 280094 255004 280100
rect 254860 206984 254912 206990
rect 254860 206926 254912 206932
rect 254768 112940 254820 112946
rect 254768 112882 254820 112888
rect 254676 92472 254728 92478
rect 254676 92414 254728 92420
rect 255872 52556 255924 52562
rect 255872 52498 255924 52504
rect 254584 48612 254636 48618
rect 254584 48554 254636 48560
rect 253664 48136 253716 48142
rect 253664 48078 253716 48084
rect 253676 12442 253704 48078
rect 255320 47592 255372 47598
rect 255320 47534 255372 47540
rect 253756 47524 253808 47530
rect 253756 47466 253808 47472
rect 253768 20466 253796 47466
rect 253940 44872 253992 44878
rect 253940 44814 253992 44820
rect 253756 20460 253808 20466
rect 253756 20402 253808 20408
rect 253952 16574 253980 44814
rect 255332 16574 255360 47534
rect 255884 17950 255912 52498
rect 255976 51066 256004 285874
rect 256068 98433 256096 295326
rect 256160 131073 256188 300834
rect 256252 208593 256280 317426
rect 256344 231033 256372 321574
rect 256700 311840 256752 311846
rect 256700 311782 256752 311788
rect 256712 310593 256740 311782
rect 256698 310584 256754 310593
rect 256698 310519 256754 310528
rect 256792 309800 256844 309806
rect 256792 309742 256844 309748
rect 256700 309120 256752 309126
rect 256700 309062 256752 309068
rect 256712 308553 256740 309062
rect 256698 308544 256754 308553
rect 256698 308479 256754 308488
rect 256804 306513 256832 309742
rect 256790 306504 256846 306513
rect 256790 306439 256846 306448
rect 256700 303612 256752 303618
rect 256700 303554 256752 303560
rect 256712 302433 256740 303554
rect 256698 302424 256754 302433
rect 256698 302359 256754 302368
rect 256700 300824 256752 300830
rect 256700 300766 256752 300772
rect 256712 300393 256740 300766
rect 256698 300384 256754 300393
rect 256698 300319 256754 300328
rect 256700 299464 256752 299470
rect 256700 299406 256752 299412
rect 256712 298353 256740 299406
rect 256698 298344 256754 298353
rect 256698 298279 256754 298288
rect 256700 296676 256752 296682
rect 256700 296618 256752 296624
rect 256712 296313 256740 296618
rect 256698 296304 256754 296313
rect 256698 296239 256754 296248
rect 256700 295316 256752 295322
rect 256700 295258 256752 295264
rect 256712 294273 256740 295258
rect 256698 294264 256754 294273
rect 256698 294199 256754 294208
rect 256700 292528 256752 292534
rect 256700 292470 256752 292476
rect 256712 292233 256740 292470
rect 256698 292224 256754 292233
rect 256698 292159 256754 292168
rect 256700 291168 256752 291174
rect 256700 291110 256752 291116
rect 256712 290193 256740 291110
rect 256698 290184 256754 290193
rect 256698 290119 256754 290128
rect 256700 288380 256752 288386
rect 256700 288322 256752 288328
rect 256712 288153 256740 288322
rect 256698 288144 256754 288153
rect 256698 288079 256754 288088
rect 257356 286113 257384 327694
rect 257712 312588 257764 312594
rect 257712 312530 257764 312536
rect 257620 305652 257672 305658
rect 257620 305594 257672 305600
rect 257436 292800 257488 292806
rect 257436 292742 257488 292748
rect 257342 286104 257398 286113
rect 257342 286039 257398 286048
rect 257344 283620 257396 283626
rect 257344 283562 257396 283568
rect 256700 282872 256752 282878
rect 256700 282814 256752 282820
rect 256712 282033 256740 282814
rect 256698 282024 256754 282033
rect 256698 281959 256754 281968
rect 256700 280152 256752 280158
rect 256700 280094 256752 280100
rect 256712 279993 256740 280094
rect 256698 279984 256754 279993
rect 256698 279919 256754 279928
rect 256700 278724 256752 278730
rect 256700 278666 256752 278672
rect 256712 277953 256740 278666
rect 256698 277944 256754 277953
rect 256698 277879 256754 277888
rect 256700 276004 256752 276010
rect 256700 275946 256752 275952
rect 256712 275913 256740 275946
rect 256698 275904 256754 275913
rect 256698 275839 256754 275848
rect 256700 274644 256752 274650
rect 256700 274586 256752 274592
rect 256712 273873 256740 274586
rect 256698 273864 256754 273873
rect 256698 273799 256754 273808
rect 256700 270496 256752 270502
rect 256700 270438 256752 270444
rect 256712 269793 256740 270438
rect 256698 269784 256754 269793
rect 256698 269719 256754 269728
rect 256700 266348 256752 266354
rect 256700 266290 256752 266296
rect 256712 265713 256740 266290
rect 256698 265704 256754 265713
rect 256698 265639 256754 265648
rect 256700 264920 256752 264926
rect 256700 264862 256752 264868
rect 256712 263673 256740 264862
rect 256698 263664 256754 263673
rect 256698 263599 256754 263608
rect 256700 262200 256752 262206
rect 256700 262142 256752 262148
rect 256712 261633 256740 262142
rect 256698 261624 256754 261633
rect 256698 261559 256754 261568
rect 256700 260840 256752 260846
rect 256700 260782 256752 260788
rect 256712 259593 256740 260782
rect 256698 259584 256754 259593
rect 256698 259519 256754 259528
rect 256700 258052 256752 258058
rect 256700 257994 256752 258000
rect 256712 257553 256740 257994
rect 256698 257544 256754 257553
rect 256698 257479 256754 257488
rect 256700 256692 256752 256698
rect 256700 256634 256752 256640
rect 256712 255513 256740 256634
rect 256698 255504 256754 255513
rect 256698 255439 256754 255448
rect 256700 253904 256752 253910
rect 256700 253846 256752 253852
rect 256712 253473 256740 253846
rect 256698 253464 256754 253473
rect 256698 253399 256754 253408
rect 256700 252544 256752 252550
rect 256700 252486 256752 252492
rect 256712 251433 256740 252486
rect 256698 251424 256754 251433
rect 256698 251359 256754 251368
rect 256700 249756 256752 249762
rect 256700 249698 256752 249704
rect 256712 249393 256740 249698
rect 256698 249384 256754 249393
rect 256698 249319 256754 249328
rect 256700 248396 256752 248402
rect 256700 248338 256752 248344
rect 256712 247353 256740 248338
rect 256698 247344 256754 247353
rect 256698 247279 256754 247288
rect 256700 245608 256752 245614
rect 256700 245550 256752 245556
rect 256712 245313 256740 245550
rect 256698 245304 256754 245313
rect 256698 245239 256754 245248
rect 256700 244248 256752 244254
rect 256700 244190 256752 244196
rect 256712 243273 256740 244190
rect 256698 243264 256754 243273
rect 256698 243199 256754 243208
rect 256700 241460 256752 241466
rect 256700 241402 256752 241408
rect 256712 241233 256740 241402
rect 256698 241224 256754 241233
rect 256698 241159 256754 241168
rect 256700 240100 256752 240106
rect 256700 240042 256752 240048
rect 256712 239193 256740 240042
rect 256698 239184 256754 239193
rect 256698 239119 256754 239128
rect 256700 237380 256752 237386
rect 256700 237322 256752 237328
rect 256712 237153 256740 237322
rect 256698 237144 256754 237153
rect 256698 237079 256754 237088
rect 257356 235113 257384 283562
rect 257448 271833 257476 292742
rect 257632 284073 257660 305594
rect 257724 304473 257752 312530
rect 257710 304464 257766 304473
rect 257710 304399 257766 304408
rect 257804 289808 257856 289814
rect 257804 289750 257856 289756
rect 257618 284064 257674 284073
rect 257618 283999 257674 284008
rect 257434 271824 257490 271833
rect 257434 271759 257490 271768
rect 257816 267753 257844 289750
rect 257802 267744 257858 267753
rect 257802 267679 257858 267688
rect 257436 267028 257488 267034
rect 257436 266970 257488 266976
rect 257342 235104 257398 235113
rect 257342 235039 257398 235048
rect 257344 233912 257396 233918
rect 257344 233854 257396 233860
rect 256700 233232 256752 233238
rect 256700 233174 256752 233180
rect 256712 233073 256740 233174
rect 256698 233064 256754 233073
rect 256698 232999 256754 233008
rect 256330 231024 256386 231033
rect 256330 230959 256386 230968
rect 256700 229016 256752 229022
rect 256698 228984 256700 228993
rect 256752 228984 256754 228993
rect 256698 228919 256754 228928
rect 256700 227724 256752 227730
rect 256700 227666 256752 227672
rect 256712 226953 256740 227666
rect 256698 226944 256754 226953
rect 256698 226879 256754 226888
rect 256700 224936 256752 224942
rect 256698 224904 256700 224913
rect 256752 224904 256754 224913
rect 256698 224839 256754 224848
rect 256700 223576 256752 223582
rect 256700 223518 256752 223524
rect 256712 222873 256740 223518
rect 256698 222864 256754 222873
rect 256698 222799 256754 222808
rect 256698 220824 256754 220833
rect 256698 220759 256700 220768
rect 256752 220759 256754 220768
rect 256700 220730 256752 220736
rect 256700 219428 256752 219434
rect 256700 219370 256752 219376
rect 256712 218793 256740 219370
rect 256698 218784 256754 218793
rect 256698 218719 256754 218728
rect 256700 218000 256752 218006
rect 256700 217942 256752 217948
rect 256712 216753 256740 217942
rect 256698 216744 256754 216753
rect 256698 216679 256754 216688
rect 256700 215280 256752 215286
rect 256700 215222 256752 215228
rect 256712 214713 256740 215222
rect 256698 214704 256754 214713
rect 256698 214639 256754 214648
rect 256700 213920 256752 213926
rect 256700 213862 256752 213868
rect 256712 212673 256740 213862
rect 256698 212664 256754 212673
rect 256698 212599 256754 212608
rect 256700 211132 256752 211138
rect 256700 211074 256752 211080
rect 256712 210633 256740 211074
rect 256698 210624 256754 210633
rect 256698 210559 256754 210568
rect 256238 208584 256294 208593
rect 256238 208519 256294 208528
rect 256700 206984 256752 206990
rect 256700 206926 256752 206932
rect 256712 206553 256740 206926
rect 256698 206544 256754 206553
rect 256698 206479 256754 206488
rect 256700 205624 256752 205630
rect 256700 205566 256752 205572
rect 256712 204513 256740 205566
rect 256698 204504 256754 204513
rect 256698 204439 256754 204448
rect 256700 202836 256752 202842
rect 256700 202778 256752 202784
rect 256712 202473 256740 202778
rect 256698 202464 256754 202473
rect 256698 202399 256754 202408
rect 256700 201476 256752 201482
rect 256700 201418 256752 201424
rect 256712 200433 256740 201418
rect 256698 200424 256754 200433
rect 256698 200359 256754 200368
rect 256700 198688 256752 198694
rect 256700 198630 256752 198636
rect 256712 198393 256740 198630
rect 256698 198384 256754 198393
rect 256698 198319 256754 198328
rect 256700 197328 256752 197334
rect 256700 197270 256752 197276
rect 256712 196353 256740 197270
rect 256698 196344 256754 196353
rect 256698 196279 256754 196288
rect 256700 194540 256752 194546
rect 256700 194482 256752 194488
rect 256712 194313 256740 194482
rect 256698 194304 256754 194313
rect 256698 194239 256754 194248
rect 256700 193180 256752 193186
rect 256700 193122 256752 193128
rect 256712 192273 256740 193122
rect 256698 192264 256754 192273
rect 256698 192199 256754 192208
rect 256700 190460 256752 190466
rect 256700 190402 256752 190408
rect 256712 190233 256740 190402
rect 256698 190224 256754 190233
rect 256698 190159 256754 190168
rect 256700 189032 256752 189038
rect 256700 188974 256752 188980
rect 256712 188193 256740 188974
rect 256698 188184 256754 188193
rect 256698 188119 256754 188128
rect 256700 186312 256752 186318
rect 256700 186254 256752 186260
rect 256712 186153 256740 186254
rect 256698 186144 256754 186153
rect 256698 186079 256754 186088
rect 256700 184884 256752 184890
rect 256700 184826 256752 184832
rect 256712 184113 256740 184826
rect 256698 184104 256754 184113
rect 256698 184039 256754 184048
rect 256700 182164 256752 182170
rect 256700 182106 256752 182112
rect 256712 182073 256740 182106
rect 256698 182064 256754 182073
rect 256698 181999 256754 182008
rect 256700 180804 256752 180810
rect 256700 180746 256752 180752
rect 256712 180033 256740 180746
rect 256698 180024 256754 180033
rect 256698 179959 256754 179968
rect 256700 178016 256752 178022
rect 256698 177984 256700 177993
rect 256752 177984 256754 177993
rect 256698 177919 256754 177928
rect 256700 176656 256752 176662
rect 256700 176598 256752 176604
rect 256712 175953 256740 176598
rect 256698 175944 256754 175953
rect 256698 175879 256754 175888
rect 256700 172508 256752 172514
rect 256700 172450 256752 172456
rect 256712 171873 256740 172450
rect 256698 171864 256754 171873
rect 256698 171799 256754 171808
rect 256700 171080 256752 171086
rect 256700 171022 256752 171028
rect 256712 169833 256740 171022
rect 256698 169824 256754 169833
rect 256698 169759 256754 169768
rect 256700 168360 256752 168366
rect 256700 168302 256752 168308
rect 256712 167793 256740 168302
rect 256698 167784 256754 167793
rect 256698 167719 256754 167728
rect 256700 167000 256752 167006
rect 256700 166942 256752 166948
rect 256712 165753 256740 166942
rect 256698 165744 256754 165753
rect 256698 165679 256754 165688
rect 256700 164212 256752 164218
rect 256700 164154 256752 164160
rect 256712 163713 256740 164154
rect 256698 163704 256754 163713
rect 256698 163639 256754 163648
rect 256700 162852 256752 162858
rect 256700 162794 256752 162800
rect 256712 161673 256740 162794
rect 256698 161664 256754 161673
rect 256698 161599 256754 161608
rect 256700 160064 256752 160070
rect 256700 160006 256752 160012
rect 256712 159633 256740 160006
rect 256698 159624 256754 159633
rect 256698 159559 256754 159568
rect 256700 155916 256752 155922
rect 256700 155858 256752 155864
rect 256712 155553 256740 155858
rect 256698 155544 256754 155553
rect 256698 155479 256754 155488
rect 256700 154556 256752 154562
rect 256700 154498 256752 154504
rect 256712 153513 256740 154498
rect 256698 153504 256754 153513
rect 256698 153439 256754 153448
rect 256700 151768 256752 151774
rect 256700 151710 256752 151716
rect 256712 151473 256740 151710
rect 256698 151464 256754 151473
rect 256698 151399 256754 151408
rect 256700 150408 256752 150414
rect 256700 150350 256752 150356
rect 256712 149433 256740 150350
rect 256698 149424 256754 149433
rect 256698 149359 256754 149368
rect 256700 147620 256752 147626
rect 256700 147562 256752 147568
rect 256712 147393 256740 147562
rect 256698 147384 256754 147393
rect 256698 147319 256754 147328
rect 256700 146260 256752 146266
rect 256700 146202 256752 146208
rect 256712 145353 256740 146202
rect 256698 145344 256754 145353
rect 256698 145279 256754 145288
rect 256700 143540 256752 143546
rect 256700 143482 256752 143488
rect 256712 143313 256740 143482
rect 256698 143304 256754 143313
rect 256698 143239 256754 143248
rect 256700 142112 256752 142118
rect 256700 142054 256752 142060
rect 256712 141273 256740 142054
rect 256698 141264 256754 141273
rect 256698 141199 256754 141208
rect 256700 139392 256752 139398
rect 256700 139334 256752 139340
rect 256712 139233 256740 139334
rect 256698 139224 256754 139233
rect 256698 139159 256754 139168
rect 256700 135244 256752 135250
rect 256700 135186 256752 135192
rect 256712 135153 256740 135186
rect 256698 135144 256754 135153
rect 256698 135079 256754 135088
rect 256700 133884 256752 133890
rect 256700 133826 256752 133832
rect 256712 133113 256740 133826
rect 256698 133104 256754 133113
rect 256698 133039 256754 133048
rect 256146 131064 256202 131073
rect 256146 130999 256202 131008
rect 256700 129736 256752 129742
rect 256700 129678 256752 129684
rect 256712 129033 256740 129678
rect 256698 129024 256754 129033
rect 256698 128959 256754 128968
rect 256698 126984 256754 126993
rect 256698 126919 256700 126928
rect 256752 126919 256754 126928
rect 256700 126890 256752 126896
rect 256700 125588 256752 125594
rect 256700 125530 256752 125536
rect 256712 124953 256740 125530
rect 256698 124944 256754 124953
rect 256698 124879 256754 124888
rect 256700 121440 256752 121446
rect 256700 121382 256752 121388
rect 256712 120873 256740 121382
rect 256698 120864 256754 120873
rect 256698 120799 256754 120808
rect 256700 120080 256752 120086
rect 256700 120022 256752 120028
rect 256712 118833 256740 120022
rect 256698 118824 256754 118833
rect 256698 118759 256754 118768
rect 256700 117292 256752 117298
rect 256700 117234 256752 117240
rect 256712 116793 256740 117234
rect 256698 116784 256754 116793
rect 256698 116719 256754 116728
rect 256700 115932 256752 115938
rect 256700 115874 256752 115880
rect 256712 114753 256740 115874
rect 256698 114744 256754 114753
rect 256698 114679 256754 114688
rect 256700 112940 256752 112946
rect 256700 112882 256752 112888
rect 256712 112713 256740 112882
rect 256698 112704 256754 112713
rect 256698 112639 256754 112648
rect 256700 111784 256752 111790
rect 256700 111726 256752 111732
rect 256712 110673 256740 111726
rect 256698 110664 256754 110673
rect 256698 110599 256754 110608
rect 256700 108996 256752 109002
rect 256700 108938 256752 108944
rect 256712 108633 256740 108938
rect 256698 108624 256754 108633
rect 256698 108559 256754 108568
rect 256700 107636 256752 107642
rect 256700 107578 256752 107584
rect 256712 106593 256740 107578
rect 256698 106584 256754 106593
rect 256698 106519 256754 106528
rect 256700 104848 256752 104854
rect 256700 104790 256752 104796
rect 256712 104553 256740 104790
rect 256698 104544 256754 104553
rect 256698 104479 256754 104488
rect 256700 103488 256752 103494
rect 256700 103430 256752 103436
rect 256712 102513 256740 103430
rect 256698 102504 256754 102513
rect 256698 102439 256754 102448
rect 256700 100700 256752 100706
rect 256700 100642 256752 100648
rect 256712 100473 256740 100642
rect 256698 100464 256754 100473
rect 256698 100399 256754 100408
rect 256054 98424 256110 98433
rect 256054 98359 256110 98368
rect 256700 96620 256752 96626
rect 256700 96562 256752 96568
rect 256712 96393 256740 96562
rect 256698 96384 256754 96393
rect 256698 96319 256754 96328
rect 256700 95192 256752 95198
rect 256700 95134 256752 95140
rect 256712 94353 256740 95134
rect 256698 94344 256754 94353
rect 256698 94279 256754 94288
rect 256700 92472 256752 92478
rect 256700 92414 256752 92420
rect 256712 92313 256740 92414
rect 256698 92304 256754 92313
rect 256698 92239 256754 92248
rect 256700 91044 256752 91050
rect 256700 90986 256752 90992
rect 256712 90273 256740 90986
rect 256698 90264 256754 90273
rect 256698 90199 256754 90208
rect 256700 88324 256752 88330
rect 256700 88266 256752 88272
rect 256712 88233 256740 88266
rect 256698 88224 256754 88233
rect 256698 88159 256754 88168
rect 256700 86964 256752 86970
rect 256700 86906 256752 86912
rect 256712 86193 256740 86906
rect 256698 86184 256754 86193
rect 256698 86119 256754 86128
rect 256700 84176 256752 84182
rect 256698 84144 256700 84153
rect 256752 84144 256754 84153
rect 256698 84079 256754 84088
rect 256700 82816 256752 82822
rect 256700 82758 256752 82764
rect 256712 82113 256740 82758
rect 256698 82104 256754 82113
rect 256698 82039 256754 82048
rect 256698 80064 256754 80073
rect 256698 79999 256700 80008
rect 256752 79999 256754 80008
rect 256700 79970 256752 79976
rect 256700 78668 256752 78674
rect 256700 78610 256752 78616
rect 256712 78033 256740 78610
rect 256698 78024 256754 78033
rect 256698 77959 256754 77968
rect 256700 77240 256752 77246
rect 256700 77182 256752 77188
rect 256712 75993 256740 77182
rect 256698 75984 256754 75993
rect 256698 75919 256754 75928
rect 256700 74520 256752 74526
rect 256700 74462 256752 74468
rect 256712 73953 256740 74462
rect 256698 73944 256754 73953
rect 256698 73879 256754 73888
rect 256700 73160 256752 73166
rect 256700 73102 256752 73108
rect 256712 71913 256740 73102
rect 256698 71904 256754 71913
rect 256698 71839 256754 71848
rect 256700 70372 256752 70378
rect 256700 70314 256752 70320
rect 256712 69873 256740 70314
rect 256698 69864 256754 69873
rect 256698 69799 256754 69808
rect 256700 69012 256752 69018
rect 256700 68954 256752 68960
rect 256712 67833 256740 68954
rect 256698 67824 256754 67833
rect 256698 67759 256754 67768
rect 256700 64456 256752 64462
rect 256700 64398 256752 64404
rect 256712 63753 256740 64398
rect 256698 63744 256754 63753
rect 256698 63679 256754 63688
rect 256700 62076 256752 62082
rect 256700 62018 256752 62024
rect 256712 61713 256740 62018
rect 256698 61704 256754 61713
rect 256698 61639 256754 61648
rect 256700 60716 256752 60722
rect 256700 60658 256752 60664
rect 256712 59673 256740 60658
rect 256698 59664 256754 59673
rect 256698 59599 256754 59608
rect 256700 57928 256752 57934
rect 256700 57870 256752 57876
rect 256712 57633 256740 57870
rect 256698 57624 256754 57633
rect 256698 57559 256754 57568
rect 256700 56568 256752 56574
rect 256700 56510 256752 56516
rect 256712 55593 256740 56510
rect 256698 55584 256754 55593
rect 256698 55519 256754 55528
rect 256700 54528 256752 54534
rect 256700 54470 256752 54476
rect 256712 51513 256740 54470
rect 257356 53553 257384 233854
rect 257448 157593 257476 266970
rect 257804 238060 257856 238066
rect 257804 238002 257856 238008
rect 257816 173913 257844 238002
rect 257802 173904 257858 173913
rect 257802 173839 257858 173848
rect 257528 158024 257580 158030
rect 257528 157966 257580 157972
rect 257434 157584 257490 157593
rect 257434 157519 257490 157528
rect 257436 140072 257488 140078
rect 257436 140014 257488 140020
rect 257448 65793 257476 140014
rect 257540 137193 257568 157966
rect 257526 137184 257582 137193
rect 257526 137119 257582 137128
rect 257434 65784 257490 65793
rect 257434 65719 257490 65728
rect 257342 53544 257398 53553
rect 257342 53479 257398 53488
rect 258736 52154 258764 351902
rect 551284 271924 551336 271930
rect 551284 271866 551336 271872
rect 550088 151836 550140 151842
rect 550088 151778 550140 151784
rect 258724 52148 258776 52154
rect 258724 52090 258776 52096
rect 258816 51604 258868 51610
rect 258816 51546 258868 51552
rect 256698 51504 256754 51513
rect 256332 51468 256384 51474
rect 256698 51439 256754 51448
rect 256332 51410 256384 51416
rect 256240 51400 256292 51406
rect 256240 51342 256292 51348
rect 256148 51332 256200 51338
rect 256148 51274 256200 51280
rect 255964 51060 256016 51066
rect 255964 51002 256016 51008
rect 256056 49768 256108 49774
rect 256056 49710 256108 49716
rect 255964 47728 256016 47734
rect 255964 47670 256016 47676
rect 255872 17944 255924 17950
rect 255872 17886 255924 17892
rect 253952 16546 254256 16574
rect 255332 16546 255912 16574
rect 253664 12436 253716 12442
rect 253664 12378 253716 12384
rect 253572 9444 253624 9450
rect 253572 9386 253624 9392
rect 253388 6044 253440 6050
rect 253388 5986 253440 5992
rect 252376 3460 252428 3466
rect 253308 3454 253520 3482
rect 252376 3402 252428 3408
rect 251192 3318 251312 3346
rect 251192 480 251220 3318
rect 252388 480 252416 3402
rect 253492 480 253520 3454
rect 248758 354 248870 480
rect 248432 326 248870 354
rect 248758 -960 248870 326
rect 249954 -960 250066 480
rect 251150 -960 251262 480
rect 252346 -960 252458 480
rect 253450 -960 253562 480
rect 254228 354 254256 16546
rect 255884 480 255912 16546
rect 255976 3262 256004 47670
rect 256068 3466 256096 49710
rect 256160 6118 256188 51274
rect 256252 6798 256280 51342
rect 256240 6792 256292 6798
rect 256240 6734 256292 6740
rect 256344 6458 256372 51410
rect 256700 51060 256752 51066
rect 256700 51002 256752 51008
rect 256608 50448 256660 50454
rect 256608 50390 256660 50396
rect 256424 47796 256476 47802
rect 256424 47738 256476 47744
rect 256332 6452 256384 6458
rect 256332 6394 256384 6400
rect 256148 6112 256200 6118
rect 256148 6054 256200 6060
rect 256056 3460 256108 3466
rect 256056 3402 256108 3408
rect 256436 3330 256464 47738
rect 256516 47660 256568 47666
rect 256516 47602 256568 47608
rect 256424 3324 256476 3330
rect 256424 3266 256476 3272
rect 255964 3256 256016 3262
rect 255964 3198 256016 3204
rect 256528 3194 256556 47602
rect 256620 6662 256648 50390
rect 256712 49473 256740 51002
rect 258724 50584 258776 50590
rect 258724 50526 258776 50532
rect 256698 49464 256754 49473
rect 256698 49399 256754 49408
rect 258632 49292 258684 49298
rect 258632 49234 258684 49240
rect 258080 43444 258132 43450
rect 258080 43386 258132 43392
rect 258092 16574 258120 43386
rect 258644 21622 258672 49234
rect 258632 21616 258684 21622
rect 258632 21558 258684 21564
rect 258092 16546 258304 16574
rect 256608 6656 256660 6662
rect 256608 6598 256660 6604
rect 257068 3392 257120 3398
rect 257068 3334 257120 3340
rect 256516 3188 256568 3194
rect 256516 3130 256568 3136
rect 257080 480 257108 3334
rect 258276 480 258304 16546
rect 258736 3602 258764 50526
rect 258828 4010 258856 51546
rect 260104 49428 260156 49434
rect 260104 49370 260156 49376
rect 259000 49360 259052 49366
rect 259000 49302 259052 49308
rect 260116 49314 260144 49370
rect 258908 49224 258960 49230
rect 258908 49166 258960 49172
rect 258816 4004 258868 4010
rect 258816 3946 258868 3952
rect 258920 3874 258948 49166
rect 258908 3868 258960 3874
rect 258908 3810 258960 3816
rect 259012 3738 259040 49302
rect 260116 49286 260236 49314
rect 259184 49156 259236 49162
rect 259184 49098 259236 49104
rect 259092 48068 259144 48074
rect 259092 48010 259144 48016
rect 259104 4078 259132 48010
rect 259196 13258 259224 49098
rect 259276 49088 259328 49094
rect 259276 49030 259328 49036
rect 259288 14890 259316 49030
rect 259368 49020 259420 49026
rect 259368 48962 259420 48968
rect 259380 20330 259408 48962
rect 259460 46232 259512 46238
rect 259460 46174 259512 46180
rect 260102 46200 260158 46209
rect 259368 20324 259420 20330
rect 259368 20266 259420 20272
rect 259276 14884 259328 14890
rect 259276 14826 259328 14832
rect 259184 13252 259236 13258
rect 259184 13194 259236 13200
rect 259092 4072 259144 4078
rect 259092 4014 259144 4020
rect 259000 3732 259052 3738
rect 259000 3674 259052 3680
rect 258724 3596 258776 3602
rect 258724 3538 258776 3544
rect 259472 480 259500 46174
rect 260102 46135 260158 46144
rect 260116 3942 260144 46135
rect 260208 18630 260236 49286
rect 550100 41177 550128 151778
rect 550180 111852 550232 111858
rect 550180 111794 550232 111800
rect 550086 41168 550142 41177
rect 550192 41138 550220 111794
rect 550086 41103 550142 41112
rect 550180 41132 550232 41138
rect 550180 41074 550232 41080
rect 287060 40860 287112 40866
rect 287060 40802 287112 40808
rect 266358 36544 266414 36553
rect 266358 36479 266414 36488
rect 260840 21684 260892 21690
rect 260840 21626 260892 21632
rect 260196 18624 260248 18630
rect 260196 18566 260248 18572
rect 260852 16574 260880 21626
rect 262220 20596 262272 20602
rect 262220 20538 262272 20544
rect 262232 16574 262260 20538
rect 266372 16574 266400 36479
rect 285678 35592 285734 35601
rect 285678 35527 285734 35536
rect 281540 28620 281592 28626
rect 281540 28562 281592 28568
rect 269764 20528 269816 20534
rect 269764 20470 269816 20476
rect 260852 16546 261800 16574
rect 262232 16546 262536 16574
rect 266372 16546 266584 16574
rect 260654 4040 260710 4049
rect 260654 3975 260710 3984
rect 260104 3936 260156 3942
rect 260104 3878 260156 3884
rect 260668 480 260696 3975
rect 261772 480 261800 16546
rect 254646 354 254758 480
rect 254228 326 254758 354
rect 254646 -960 254758 326
rect 255842 -960 255954 480
rect 257038 -960 257150 480
rect 258234 -960 258346 480
rect 259430 -960 259542 480
rect 260626 -960 260738 480
rect 261730 -960 261842 480
rect 262508 354 262536 16546
rect 264978 13560 265034 13569
rect 264978 13495 265034 13504
rect 264150 3904 264206 3913
rect 264150 3839 264206 3848
rect 264164 480 264192 3839
rect 262926 354 263038 480
rect 262508 326 263038 354
rect 262926 -960 263038 326
rect 264122 -960 264234 480
rect 264992 354 265020 13495
rect 266556 480 266584 16546
rect 268382 13424 268438 13433
rect 268382 13359 268438 13368
rect 267738 3768 267794 3777
rect 267738 3703 267794 3712
rect 267752 480 267780 3703
rect 265318 354 265430 480
rect 264992 326 265430 354
rect 265318 -960 265430 326
rect 266514 -960 266626 480
rect 267710 -960 267822 480
rect 268396 354 268424 13359
rect 269776 6866 269804 20470
rect 273260 19236 273312 19242
rect 273260 19178 273312 19184
rect 271142 14784 271198 14793
rect 271142 14719 271198 14728
rect 269764 6860 269816 6866
rect 269764 6802 269816 6808
rect 270040 6724 270092 6730
rect 270040 6666 270092 6672
rect 270052 480 270080 6666
rect 271156 3466 271184 14719
rect 272432 13320 272484 13326
rect 272432 13262 272484 13268
rect 271144 3460 271196 3466
rect 271144 3402 271196 3408
rect 271236 3188 271288 3194
rect 271236 3130 271288 3136
rect 271248 480 271276 3130
rect 272444 480 272472 13262
rect 268814 354 268926 480
rect 268396 326 268926 354
rect 268814 -960 268926 326
rect 270010 -960 270122 480
rect 271206 -960 271318 480
rect 272402 -960 272514 480
rect 273272 354 273300 19178
rect 276020 19168 276072 19174
rect 276020 19110 276072 19116
rect 276032 4214 276060 19110
rect 280160 19100 280212 19106
rect 280160 19042 280212 19048
rect 280172 16574 280200 19042
rect 280172 16546 280752 16574
rect 276112 11688 276164 11694
rect 276112 11630 276164 11636
rect 276020 4208 276072 4214
rect 276020 4150 276072 4156
rect 276124 3482 276152 11630
rect 279056 10600 279108 10606
rect 279056 10542 279108 10548
rect 276756 4208 276808 4214
rect 276756 4150 276808 4156
rect 276032 3454 276152 3482
rect 274824 3256 274876 3262
rect 274824 3198 274876 3204
rect 274836 480 274864 3198
rect 276032 480 276060 3454
rect 273598 354 273710 480
rect 273272 326 273710 354
rect 273598 -960 273710 326
rect 274794 -960 274906 480
rect 275990 -960 276102 480
rect 276768 354 276796 4150
rect 278318 3632 278374 3641
rect 278318 3567 278374 3576
rect 278332 480 278360 3567
rect 277094 354 277206 480
rect 276768 326 277206 354
rect 277094 -960 277206 326
rect 278290 -960 278402 480
rect 279068 354 279096 10542
rect 280724 480 280752 16546
rect 279486 354 279598 480
rect 279068 326 279598 354
rect 279486 -960 279598 326
rect 280682 -960 280794 480
rect 281552 354 281580 28562
rect 284298 24440 284354 24449
rect 284298 24375 284354 24384
rect 283102 13288 283158 13297
rect 283102 13223 283158 13232
rect 283116 480 283144 13223
rect 284312 4214 284340 24375
rect 284390 17640 284446 17649
rect 284390 17575 284446 17584
rect 284300 4208 284352 4214
rect 284300 4150 284352 4156
rect 284404 3482 284432 17575
rect 285692 16574 285720 35527
rect 287072 16574 287100 40802
rect 350540 40792 350592 40798
rect 350540 40734 350592 40740
rect 347780 39568 347832 39574
rect 347780 39510 347832 39516
rect 332600 38344 332652 38350
rect 332600 38286 332652 38292
rect 318798 37904 318854 37913
rect 318798 37839 318854 37848
rect 298100 35488 298152 35494
rect 298100 35430 298152 35436
rect 292672 27260 292724 27266
rect 292672 27202 292724 27208
rect 291200 19032 291252 19038
rect 291200 18974 291252 18980
rect 291212 16574 291240 18974
rect 292684 16574 292712 27202
rect 293960 18964 294012 18970
rect 293960 18906 294012 18912
rect 293972 16574 294000 18906
rect 285692 16546 286640 16574
rect 287072 16546 287376 16574
rect 291212 16546 291424 16574
rect 292684 16546 293264 16574
rect 293972 16546 294920 16574
rect 285036 4208 285088 4214
rect 285036 4150 285088 4156
rect 284312 3454 284432 3482
rect 284312 480 284340 3454
rect 281878 354 281990 480
rect 281552 326 281990 354
rect 281878 -960 281990 326
rect 283074 -960 283186 480
rect 284270 -960 284382 480
rect 285048 354 285076 4150
rect 286612 480 286640 16546
rect 285374 354 285486 480
rect 285048 326 285486 354
rect 285374 -960 285486 326
rect 286570 -960 286682 480
rect 287348 354 287376 16546
rect 290188 6044 290240 6050
rect 290188 5986 290240 5992
rect 288992 3324 289044 3330
rect 288992 3266 289044 3272
rect 289004 480 289032 3266
rect 290200 480 290228 5986
rect 291396 480 291424 16546
rect 292580 3392 292632 3398
rect 292580 3334 292632 3340
rect 292592 480 292620 3334
rect 287766 354 287878 480
rect 287348 326 287878 354
rect 287766 -960 287878 326
rect 288962 -960 289074 480
rect 290158 -960 290270 480
rect 291354 -960 291466 480
rect 292550 -960 292662 480
rect 293236 354 293264 16546
rect 294892 480 294920 16546
rect 297272 10532 297324 10538
rect 297272 10474 297324 10480
rect 296076 4140 296128 4146
rect 296076 4082 296128 4088
rect 296088 480 296116 4082
rect 297284 480 297312 10474
rect 293654 354 293766 480
rect 293236 326 293766 354
rect 293654 -960 293766 326
rect 294850 -960 294962 480
rect 296046 -960 296158 480
rect 297242 -960 297354 480
rect 298112 354 298140 35430
rect 303618 34232 303674 34241
rect 303618 34167 303674 34176
rect 299480 23384 299532 23390
rect 299480 23326 299532 23332
rect 299492 3398 299520 23326
rect 300858 18592 300914 18601
rect 300858 18527 300914 18536
rect 300872 16574 300900 18527
rect 303632 16574 303660 34167
rect 311900 31340 311952 31346
rect 311900 31282 311952 31288
rect 307760 28552 307812 28558
rect 307760 28494 307812 28500
rect 305000 18896 305052 18902
rect 305000 18838 305052 18844
rect 305012 16574 305040 18838
rect 300872 16546 301544 16574
rect 303632 16546 303936 16574
rect 305012 16546 305592 16574
rect 299664 6588 299716 6594
rect 299664 6530 299716 6536
rect 299480 3392 299532 3398
rect 299480 3334 299532 3340
rect 299676 480 299704 6530
rect 300768 3392 300820 3398
rect 300768 3334 300820 3340
rect 300780 480 300808 3334
rect 298438 354 298550 480
rect 298112 326 298550 354
rect 298438 -960 298550 326
rect 299634 -960 299746 480
rect 300738 -960 300850 480
rect 301516 354 301544 16546
rect 303158 6760 303214 6769
rect 303158 6695 303214 6704
rect 303172 480 303200 6695
rect 301934 354 302046 480
rect 301516 326 302046 354
rect 301934 -960 302046 326
rect 303130 -960 303242 480
rect 303908 354 303936 16546
rect 305564 480 305592 16546
rect 306748 6112 306800 6118
rect 306748 6054 306800 6060
rect 306760 480 306788 6054
rect 307772 3398 307800 28494
rect 309140 28484 309192 28490
rect 309140 28426 309192 28432
rect 309152 16574 309180 28426
rect 311912 16574 311940 31282
rect 313280 29980 313332 29986
rect 313280 29922 313332 29928
rect 313292 16574 313320 29922
rect 316040 24472 316092 24478
rect 316040 24414 316092 24420
rect 309152 16546 309824 16574
rect 311912 16546 312216 16574
rect 313292 16546 313872 16574
rect 307944 5160 307996 5166
rect 307944 5102 307996 5108
rect 307760 3392 307812 3398
rect 307760 3334 307812 3340
rect 307956 480 307984 5102
rect 309048 3392 309100 3398
rect 309048 3334 309100 3340
rect 309060 480 309088 3334
rect 304326 354 304438 480
rect 303908 326 304438 354
rect 304326 -960 304438 326
rect 305522 -960 305634 480
rect 306718 -960 306830 480
rect 307914 -960 308026 480
rect 309018 -960 309130 480
rect 309796 354 309824 16546
rect 311440 6520 311492 6526
rect 311440 6462 311492 6468
rect 311452 480 311480 6462
rect 310214 354 310326 480
rect 309796 326 310326 354
rect 310214 -960 310326 326
rect 311410 -960 311522 480
rect 312188 354 312216 16546
rect 313844 480 313872 16546
rect 315028 8016 315080 8022
rect 315028 7958 315080 7964
rect 315040 480 315068 7958
rect 316052 3398 316080 24414
rect 316132 17196 316184 17202
rect 316132 17138 316184 17144
rect 316144 16574 316172 17138
rect 318812 16574 318840 37839
rect 324320 33924 324372 33930
rect 324320 33866 324372 33872
rect 320178 29880 320234 29889
rect 320178 29815 320234 29824
rect 320192 16574 320220 29815
rect 316144 16546 316264 16574
rect 318812 16546 319760 16574
rect 320192 16546 320496 16574
rect 316040 3392 316092 3398
rect 316040 3334 316092 3340
rect 316236 480 316264 16546
rect 318062 13152 318118 13161
rect 318062 13087 318118 13096
rect 317328 3392 317380 3398
rect 317328 3334 317380 3340
rect 317340 480 317368 3334
rect 312606 354 312718 480
rect 312188 326 312718 354
rect 312606 -960 312718 326
rect 313802 -960 313914 480
rect 314998 -960 315110 480
rect 316194 -960 316306 480
rect 317298 -960 317410 480
rect 318076 354 318104 13087
rect 319732 480 319760 16546
rect 318494 354 318606 480
rect 318076 326 318606 354
rect 318494 -960 318606 326
rect 319690 -960 319802 480
rect 320468 354 320496 16546
rect 322110 14648 322166 14657
rect 322110 14583 322166 14592
rect 322124 480 322152 14583
rect 323308 5092 323360 5098
rect 323308 5034 323360 5040
rect 323320 480 323348 5034
rect 324332 3210 324360 33866
rect 324412 33856 324464 33862
rect 324412 33798 324464 33804
rect 324424 3398 324452 33798
rect 331220 31272 331272 31278
rect 331220 31214 331272 31220
rect 325700 23316 325752 23322
rect 325700 23258 325752 23264
rect 325712 16574 325740 23258
rect 329840 18828 329892 18834
rect 329840 18770 329892 18776
rect 329852 16574 329880 18770
rect 325712 16546 326384 16574
rect 329852 16546 330432 16574
rect 324412 3392 324464 3398
rect 324412 3334 324464 3340
rect 325608 3392 325660 3398
rect 325608 3334 325660 3340
rect 324332 3182 324452 3210
rect 324424 480 324452 3182
rect 325620 480 325648 3334
rect 320886 354 320998 480
rect 320468 326 320998 354
rect 320886 -960 320998 326
rect 322082 -960 322194 480
rect 323278 -960 323390 480
rect 324382 -960 324494 480
rect 325578 -960 325690 480
rect 326356 354 326384 16546
rect 328736 14340 328788 14346
rect 328736 14282 328788 14288
rect 328000 6792 328052 6798
rect 328000 6734 328052 6740
rect 328012 480 328040 6734
rect 326774 354 326886 480
rect 326356 326 326886 354
rect 326774 -960 326886 326
rect 327970 -960 328082 480
rect 328748 354 328776 14282
rect 330404 480 330432 16546
rect 329166 354 329278 480
rect 328748 326 329278 354
rect 329166 -960 329278 326
rect 330362 -960 330474 480
rect 331232 354 331260 31214
rect 332612 3398 332640 38286
rect 340880 29912 340932 29918
rect 340880 29854 340932 29860
rect 338118 29744 338174 29753
rect 338118 29679 338174 29688
rect 333980 25764 334032 25770
rect 333980 25706 334032 25712
rect 333992 16574 334020 25706
rect 336738 21856 336794 21865
rect 336738 21791 336794 21800
rect 336752 16574 336780 21791
rect 338132 16574 338160 29679
rect 340892 16574 340920 29854
rect 345020 27192 345072 27198
rect 345020 27134 345072 27140
rect 345032 16574 345060 27134
rect 347792 16574 347820 39510
rect 349160 23248 349212 23254
rect 349160 23190 349212 23196
rect 349172 16574 349200 23190
rect 350552 16574 350580 40734
rect 382280 40724 382332 40730
rect 382280 40666 382332 40672
rect 357440 39500 357492 39506
rect 357440 39442 357492 39448
rect 353298 21720 353354 21729
rect 353298 21655 353354 21664
rect 353312 16574 353340 21655
rect 333992 16546 334664 16574
rect 336752 16546 337056 16574
rect 338132 16546 338712 16574
rect 340892 16546 341012 16574
rect 345032 16546 345336 16574
rect 347792 16546 348096 16574
rect 349172 16546 349292 16574
rect 350552 16546 351224 16574
rect 353312 16546 353616 16574
rect 332692 14408 332744 14414
rect 332692 14350 332744 14356
rect 332600 3392 332652 3398
rect 332600 3334 332652 3340
rect 332704 480 332732 14350
rect 333888 3392 333940 3398
rect 333888 3334 333940 3340
rect 333900 480 333928 3334
rect 331558 354 331670 480
rect 331232 326 331670 354
rect 331558 -960 331670 326
rect 332662 -960 332774 480
rect 333858 -960 333970 480
rect 334636 354 334664 16546
rect 336280 15088 336332 15094
rect 336280 15030 336332 15036
rect 336292 480 336320 15030
rect 335054 354 335166 480
rect 334636 326 335166 354
rect 335054 -960 335166 326
rect 336250 -960 336362 480
rect 337028 354 337056 16546
rect 338684 480 338712 16546
rect 339500 15156 339552 15162
rect 339500 15098 339552 15104
rect 337446 354 337558 480
rect 337028 326 337558 354
rect 337446 -960 337558 326
rect 338642 -960 338754 480
rect 339512 354 339540 15098
rect 340984 480 341012 16546
rect 342904 15020 342956 15026
rect 342904 14962 342956 14968
rect 342168 6656 342220 6662
rect 342168 6598 342220 6604
rect 342180 480 342208 6598
rect 339838 354 339950 480
rect 339512 326 339950 354
rect 339838 -960 339950 326
rect 340942 -960 341054 480
rect 342138 -960 342250 480
rect 342916 354 342944 14962
rect 344560 9648 344612 9654
rect 344560 9590 344612 9596
rect 344572 480 344600 9590
rect 343334 354 343446 480
rect 342916 326 343446 354
rect 343334 -960 343446 326
rect 344530 -960 344642 480
rect 345308 354 345336 16546
rect 346952 14952 347004 14958
rect 346952 14894 347004 14900
rect 346964 480 346992 14894
rect 348068 480 348096 16546
rect 349264 480 349292 16546
rect 350448 7948 350500 7954
rect 350448 7890 350500 7896
rect 350460 480 350488 7890
rect 345726 354 345838 480
rect 345308 326 345838 354
rect 345726 -960 345838 326
rect 346922 -960 347034 480
rect 348026 -960 348138 480
rect 349222 -960 349334 480
rect 350418 -960 350530 480
rect 351196 354 351224 16546
rect 352840 7880 352892 7886
rect 352840 7822 352892 7828
rect 352852 480 352880 7822
rect 351614 354 351726 480
rect 351196 326 351726 354
rect 351614 -960 351726 326
rect 352810 -960 352922 480
rect 353588 354 353616 16546
rect 355230 16008 355286 16017
rect 355230 15943 355286 15952
rect 355244 480 355272 15943
rect 356334 6624 356390 6633
rect 356334 6559 356390 6568
rect 356348 480 356376 6559
rect 357452 3398 357480 39442
rect 365720 39432 365772 39438
rect 365720 39374 365772 39380
rect 361580 39364 361632 39370
rect 361580 39306 361632 39312
rect 357530 32736 357586 32745
rect 357530 32671 357586 32680
rect 357440 3392 357492 3398
rect 357440 3334 357492 3340
rect 357544 480 357572 32671
rect 358820 28416 358872 28422
rect 358820 28358 358872 28364
rect 358832 16574 358860 28358
rect 361592 16574 361620 39306
rect 364340 35420 364392 35426
rect 364340 35362 364392 35368
rect 362960 24404 363012 24410
rect 362960 24346 363012 24352
rect 362972 16574 363000 24346
rect 364352 16574 364380 35362
rect 365732 16574 365760 39374
rect 372620 32564 372672 32570
rect 372620 32506 372672 32512
rect 371238 31104 371294 31113
rect 371238 31039 371294 31048
rect 368480 25696 368532 25702
rect 368480 25638 368532 25644
rect 368492 16574 368520 25638
rect 358832 16546 359504 16574
rect 361592 16546 361896 16574
rect 362972 16546 363552 16574
rect 364352 16546 364656 16574
rect 365732 16546 365852 16574
rect 368492 16546 369440 16574
rect 358728 3392 358780 3398
rect 358728 3334 358780 3340
rect 358740 480 358768 3334
rect 354006 354 354118 480
rect 353588 326 354118 354
rect 354006 -960 354118 326
rect 355202 -960 355314 480
rect 356306 -960 356418 480
rect 357502 -960 357614 480
rect 358698 -960 358810 480
rect 359476 354 359504 16546
rect 361120 9512 361172 9518
rect 361120 9454 361172 9460
rect 361132 480 361160 9454
rect 359894 354 360006 480
rect 359476 326 360006 354
rect 359894 -960 360006 326
rect 361090 -960 361202 480
rect 361868 354 361896 16546
rect 363524 480 363552 16546
rect 364628 480 364656 16546
rect 365824 480 365852 16546
rect 367008 7812 367060 7818
rect 367008 7754 367060 7760
rect 367020 480 367048 7754
rect 368204 5024 368256 5030
rect 368204 4966 368256 4972
rect 368216 480 368244 4966
rect 369412 480 369440 16546
rect 370594 6488 370650 6497
rect 370594 6423 370650 6432
rect 370608 480 370636 6423
rect 362286 354 362398 480
rect 361868 326 362398 354
rect 362286 -960 362398 326
rect 363482 -960 363594 480
rect 364586 -960 364698 480
rect 365782 -960 365894 480
rect 366978 -960 367090 480
rect 368174 -960 368286 480
rect 369370 -960 369482 480
rect 370566 -960 370678 480
rect 371252 354 371280 31039
rect 372632 16574 372660 32506
rect 373998 28520 374054 28529
rect 373998 28455 374054 28464
rect 372632 16546 372936 16574
rect 372908 480 372936 16546
rect 374012 3398 374040 28455
rect 378140 27124 378192 27130
rect 378140 27066 378192 27072
rect 374090 21584 374146 21593
rect 374090 21519 374146 21528
rect 374000 3392 374052 3398
rect 374000 3334 374052 3340
rect 374104 480 374132 21519
rect 378152 16574 378180 27066
rect 379520 20392 379572 20398
rect 379520 20334 379572 20340
rect 378152 16546 378456 16574
rect 376024 12368 376076 12374
rect 376024 12310 376076 12316
rect 375288 3392 375340 3398
rect 375288 3334 375340 3340
rect 375300 480 375328 3334
rect 371670 354 371782 480
rect 371252 326 371782 354
rect 371670 -960 371782 326
rect 372866 -960 372978 480
rect 374062 -960 374174 480
rect 375258 -960 375370 480
rect 376036 354 376064 12310
rect 377680 6452 377732 6458
rect 377680 6394 377732 6400
rect 377692 480 377720 6394
rect 376454 354 376566 480
rect 376036 326 376566 354
rect 376454 -960 376566 326
rect 377650 -960 377762 480
rect 378428 354 378456 16546
rect 378846 354 378958 480
rect 378428 326 378958 354
rect 379532 354 379560 20334
rect 381176 8900 381228 8906
rect 381176 8842 381228 8848
rect 381188 480 381216 8842
rect 382292 3398 382320 40666
rect 551296 39778 551324 271866
rect 551376 258120 551428 258126
rect 551376 258062 551428 258068
rect 551284 39772 551336 39778
rect 551284 39714 551336 39720
rect 551388 39710 551416 258062
rect 551468 231872 551520 231878
rect 551468 231814 551520 231820
rect 551480 41070 551508 231814
rect 551560 218068 551612 218074
rect 551560 218010 551612 218016
rect 551468 41064 551520 41070
rect 551468 41006 551520 41012
rect 551572 39846 551600 218010
rect 552664 178084 552716 178090
rect 552664 178026 552716 178032
rect 551652 138032 551704 138038
rect 551652 137974 551704 137980
rect 551664 39914 551692 137974
rect 551744 59424 551796 59430
rect 551744 59366 551796 59372
rect 551756 39982 551784 59366
rect 552676 41313 552704 178026
rect 552662 41304 552718 41313
rect 552662 41239 552718 41248
rect 551744 39976 551796 39982
rect 551744 39918 551796 39924
rect 551652 39908 551704 39914
rect 551652 39850 551704 39856
rect 551560 39840 551612 39846
rect 551560 39782 551612 39788
rect 551376 39704 551428 39710
rect 551376 39646 551428 39652
rect 573376 38554 573404 456758
rect 574756 38622 574784 616830
rect 580170 537840 580226 537849
rect 580170 537775 580226 537784
rect 580184 529310 580212 537775
rect 580172 529304 580224 529310
rect 580172 529246 580224 529252
rect 580170 524512 580226 524521
rect 580170 524447 580172 524456
rect 580224 524447 580226 524456
rect 580172 524418 580224 524424
rect 580170 511320 580226 511329
rect 580170 511255 580226 511264
rect 580184 510678 580212 511255
rect 580172 510672 580224 510678
rect 580172 510614 580224 510620
rect 580170 458144 580226 458153
rect 580170 458079 580226 458088
rect 580184 456822 580212 458079
rect 580172 456816 580224 456822
rect 580172 456758 580224 456764
rect 579802 378448 579858 378457
rect 579802 378383 579858 378392
rect 579816 378214 579844 378383
rect 579804 378208 579856 378214
rect 579804 378150 579856 378156
rect 579986 365120 580042 365129
rect 579986 365055 580042 365064
rect 580000 364410 580028 365055
rect 579988 364404 580040 364410
rect 579988 364346 580040 364352
rect 580172 351960 580224 351966
rect 580170 351928 580172 351937
rect 580224 351928 580226 351937
rect 580170 351863 580226 351872
rect 580170 325272 580226 325281
rect 580170 325207 580226 325216
rect 580184 324358 580212 325207
rect 580172 324352 580224 324358
rect 580172 324294 580224 324300
rect 580276 319666 580304 630799
rect 580446 591016 580502 591025
rect 580446 590951 580502 590960
rect 580354 577688 580410 577697
rect 580354 577623 580410 577632
rect 580368 319734 580396 577623
rect 580460 371890 580488 590951
rect 580552 529242 580580 643991
rect 580630 564360 580686 564369
rect 580630 564295 580686 564304
rect 580644 529378 580672 564295
rect 580632 529372 580684 529378
rect 580632 529314 580684 529320
rect 580540 529236 580592 529242
rect 580540 529178 580592 529184
rect 580538 484664 580594 484673
rect 580538 484599 580594 484608
rect 580448 371884 580500 371890
rect 580448 371826 580500 371832
rect 580356 319728 580408 319734
rect 580356 319670 580408 319676
rect 580264 319660 580316 319666
rect 580264 319602 580316 319608
rect 580552 319598 580580 484599
rect 580630 471472 580686 471481
rect 580630 471407 580686 471416
rect 580540 319592 580592 319598
rect 580540 319534 580592 319540
rect 580644 319462 580672 471407
rect 580722 431624 580778 431633
rect 580722 431559 580778 431568
rect 580736 320890 580764 431559
rect 580814 418296 580870 418305
rect 580814 418231 580870 418240
rect 580724 320884 580776 320890
rect 580724 320826 580776 320832
rect 580828 319530 580856 418231
rect 580906 404968 580962 404977
rect 580906 404903 580962 404912
rect 580920 320958 580948 404903
rect 580908 320952 580960 320958
rect 580908 320894 580960 320900
rect 580816 319524 580868 319530
rect 580816 319466 580868 319472
rect 580632 319456 580684 319462
rect 580632 319398 580684 319404
rect 580448 318844 580500 318850
rect 580448 318786 580500 318792
rect 580460 312089 580488 318786
rect 580446 312080 580502 312089
rect 580446 312015 580502 312024
rect 580262 298752 580318 298761
rect 580262 298687 580318 298696
rect 580170 272232 580226 272241
rect 580170 272167 580226 272176
rect 580184 271930 580212 272167
rect 580172 271924 580224 271930
rect 580172 271866 580224 271872
rect 580170 258904 580226 258913
rect 580170 258839 580226 258848
rect 580184 258126 580212 258839
rect 580172 258120 580224 258126
rect 580172 258062 580224 258068
rect 579618 232384 579674 232393
rect 579618 232319 579674 232328
rect 579632 231878 579660 232319
rect 579620 231872 579672 231878
rect 579620 231814 579672 231820
rect 580170 219056 580226 219065
rect 580170 218991 580226 219000
rect 580184 218074 580212 218991
rect 580172 218068 580224 218074
rect 580172 218010 580224 218016
rect 580170 179208 580226 179217
rect 580170 179143 580226 179152
rect 580184 178090 580212 179143
rect 580172 178084 580224 178090
rect 580172 178026 580224 178032
rect 579986 152688 580042 152697
rect 579986 152623 580042 152632
rect 580000 151842 580028 152623
rect 579988 151836 580040 151842
rect 579988 151778 580040 151784
rect 580170 139360 580226 139369
rect 580170 139295 580226 139304
rect 580184 138038 580212 139295
rect 580172 138032 580224 138038
rect 580172 137974 580224 137980
rect 580170 112840 580226 112849
rect 580170 112775 580226 112784
rect 580184 111858 580212 112775
rect 580172 111852 580224 111858
rect 580172 111794 580224 111800
rect 580170 72992 580226 73001
rect 580170 72927 580226 72936
rect 580078 59664 580134 59673
rect 580078 59599 580134 59608
rect 580092 59430 580120 59599
rect 580080 59424 580132 59430
rect 580080 59366 580132 59372
rect 580080 50380 580132 50386
rect 580080 50322 580132 50328
rect 580092 40050 580120 50322
rect 580184 41410 580212 72927
rect 580172 41404 580224 41410
rect 580172 41346 580224 41352
rect 580276 41274 580304 298687
rect 580354 245576 580410 245585
rect 580354 245511 580410 245520
rect 580368 41342 580396 245511
rect 580446 205728 580502 205737
rect 580446 205663 580502 205672
rect 580460 41954 580488 205663
rect 580538 192536 580594 192545
rect 580538 192471 580594 192480
rect 580448 41948 580500 41954
rect 580448 41890 580500 41896
rect 580552 41886 580580 192471
rect 580630 165880 580686 165889
rect 580630 165815 580686 165824
rect 580644 41993 580672 165815
rect 580722 126032 580778 126041
rect 580722 125967 580778 125976
rect 580736 42022 580764 125967
rect 580814 99512 580870 99521
rect 580814 99447 580870 99456
rect 580828 50386 580856 99447
rect 580906 86184 580962 86193
rect 580906 86119 580962 86128
rect 580816 50380 580868 50386
rect 580816 50322 580868 50328
rect 580814 46336 580870 46345
rect 580814 46271 580870 46280
rect 580724 42016 580776 42022
rect 580630 41984 580686 41993
rect 580724 41958 580776 41964
rect 580630 41919 580686 41928
rect 580540 41880 580592 41886
rect 580540 41822 580592 41828
rect 580356 41336 580408 41342
rect 580356 41278 580408 41284
rect 580264 41268 580316 41274
rect 580264 41210 580316 41216
rect 580828 41206 580856 46271
rect 580920 42090 580948 86119
rect 580908 42084 580960 42090
rect 580908 42026 580960 42032
rect 580816 41200 580868 41206
rect 580816 41142 580868 41148
rect 580080 40044 580132 40050
rect 580080 39986 580132 39992
rect 574744 38616 574796 38622
rect 574744 38558 574796 38564
rect 573364 38548 573416 38554
rect 573364 38490 573416 38496
rect 400220 38276 400272 38282
rect 400220 38218 400272 38224
rect 385040 37120 385092 37126
rect 385040 37062 385092 37068
rect 383660 25628 383712 25634
rect 383660 25570 383712 25576
rect 382372 24336 382424 24342
rect 382372 24278 382424 24284
rect 382280 3392 382332 3398
rect 382280 3334 382332 3340
rect 382384 480 382412 24278
rect 383672 16574 383700 25570
rect 385052 16574 385080 37062
rect 390558 35456 390614 35465
rect 390558 35391 390614 35400
rect 386420 28348 386472 28354
rect 386420 28290 386472 28296
rect 386432 16574 386460 28290
rect 390572 16574 390600 35391
rect 394700 29844 394752 29850
rect 394700 29786 394752 29792
rect 394712 16574 394740 29786
rect 396080 23180 396132 23186
rect 396080 23122 396132 23128
rect 383672 16546 384344 16574
rect 385052 16546 386000 16574
rect 386432 16546 386736 16574
rect 390572 16546 390692 16574
rect 394712 16546 395384 16574
rect 383568 3392 383620 3398
rect 383568 3334 383620 3340
rect 383580 480 383608 3334
rect 379950 354 380062 480
rect 379532 326 380062 354
rect 378846 -960 378958 326
rect 379950 -960 380062 326
rect 381146 -960 381258 480
rect 382342 -960 382454 480
rect 383538 -960 383650 480
rect 384316 354 384344 16546
rect 385972 480 386000 16546
rect 384734 354 384846 480
rect 384316 326 384846 354
rect 384734 -960 384846 326
rect 385930 -960 386042 480
rect 386708 354 386736 16546
rect 389456 12300 389508 12306
rect 389456 12242 389508 12248
rect 388260 9308 388312 9314
rect 388260 9250 388312 9256
rect 388272 480 388300 9250
rect 389468 480 389496 12242
rect 390664 480 390692 16546
rect 392582 13016 392638 13025
rect 392582 12951 392638 12960
rect 391848 9240 391900 9246
rect 391848 9182 391900 9188
rect 391860 480 391888 9182
rect 387126 354 387238 480
rect 386708 326 387238 354
rect 387126 -960 387238 326
rect 388230 -960 388342 480
rect 389426 -960 389538 480
rect 390622 -960 390734 480
rect 391818 -960 391930 480
rect 392596 354 392624 12951
rect 394240 12436 394292 12442
rect 394240 12378 394292 12384
rect 394252 480 394280 12378
rect 395356 480 395384 16546
rect 393014 354 393126 480
rect 392596 326 393126 354
rect 393014 -960 393126 326
rect 394210 -960 394322 480
rect 395314 -960 395426 480
rect 396092 354 396120 23122
rect 398840 23112 398892 23118
rect 398840 23054 398892 23060
rect 397460 17944 397512 17950
rect 397460 17886 397512 17892
rect 397472 16574 397500 17886
rect 397472 16546 397776 16574
rect 397748 480 397776 16546
rect 398852 3210 398880 23054
rect 400232 16574 400260 38218
rect 462964 38208 463016 38214
rect 462964 38150 463016 38156
rect 450544 37052 450596 37058
rect 450544 36994 450596 37000
rect 407118 34096 407174 34105
rect 407118 34031 407174 34040
rect 404360 20256 404412 20262
rect 404360 20198 404412 20204
rect 400232 16546 400904 16574
rect 398932 10464 398984 10470
rect 398932 10406 398984 10412
rect 398944 3398 398972 10406
rect 398932 3392 398984 3398
rect 398932 3334 398984 3340
rect 400128 3392 400180 3398
rect 400128 3334 400180 3340
rect 398852 3182 398972 3210
rect 398944 480 398972 3182
rect 400140 480 400168 3334
rect 396510 354 396622 480
rect 396092 326 396622 354
rect 396510 -960 396622 326
rect 397706 -960 397818 480
rect 398902 -960 399014 480
rect 400098 -960 400210 480
rect 400876 354 400904 16546
rect 403624 6384 403676 6390
rect 403624 6326 403676 6332
rect 402520 4956 402572 4962
rect 402520 4898 402572 4904
rect 402532 480 402560 4898
rect 403636 480 403664 6326
rect 401294 354 401406 480
rect 400876 326 401406 354
rect 401294 -960 401406 326
rect 402490 -960 402602 480
rect 403594 -960 403706 480
rect 404372 354 404400 20198
rect 406016 7744 406068 7750
rect 406016 7686 406068 7692
rect 406028 480 406056 7686
rect 407132 3210 407160 34031
rect 425060 31204 425112 31210
rect 425060 31146 425112 31152
rect 423678 29608 423734 29617
rect 423678 29543 423734 29552
rect 415400 27056 415452 27062
rect 415400 26998 415452 27004
rect 411260 20460 411312 20466
rect 411260 20402 411312 20408
rect 407210 20088 407266 20097
rect 407210 20023 407266 20032
rect 407224 3398 407252 20023
rect 411272 16574 411300 20402
rect 411272 16546 411944 16574
rect 410798 14512 410854 14521
rect 410798 14447 410854 14456
rect 409602 6352 409658 6361
rect 409602 6287 409658 6296
rect 407212 3392 407264 3398
rect 407212 3334 407264 3340
rect 408408 3392 408460 3398
rect 408408 3334 408460 3340
rect 407132 3182 407252 3210
rect 407224 480 407252 3182
rect 408420 480 408448 3334
rect 409616 480 409644 6287
rect 410812 480 410840 14447
rect 411916 480 411944 16546
rect 414296 16380 414348 16386
rect 414296 16322 414348 16328
rect 413100 9580 413152 9586
rect 413100 9522 413152 9528
rect 413112 480 413140 9522
rect 414308 480 414336 16322
rect 415412 3398 415440 26998
rect 415492 20188 415544 20194
rect 415492 20130 415544 20136
rect 415400 3392 415452 3398
rect 415400 3334 415452 3340
rect 415504 480 415532 20130
rect 422300 20120 422352 20126
rect 422300 20062 422352 20068
rect 418160 18760 418212 18766
rect 418160 18702 418212 18708
rect 418172 16574 418200 18702
rect 422312 16574 422340 20062
rect 418172 16546 418568 16574
rect 422312 16546 422616 16574
rect 417424 16312 417476 16318
rect 417424 16254 417476 16260
rect 416688 3392 416740 3398
rect 416688 3334 416740 3340
rect 416700 480 416728 3334
rect 404790 354 404902 480
rect 404372 326 404902 354
rect 404790 -960 404902 326
rect 405986 -960 406098 480
rect 407182 -960 407294 480
rect 408378 -960 408490 480
rect 409574 -960 409686 480
rect 410770 -960 410882 480
rect 411874 -960 411986 480
rect 413070 -960 413182 480
rect 414266 -960 414378 480
rect 415462 -960 415574 480
rect 416658 -960 416770 480
rect 417436 354 417464 16254
rect 417854 354 417966 480
rect 417436 326 417966 354
rect 418540 354 418568 16546
rect 420920 16244 420972 16250
rect 420920 16186 420972 16192
rect 420184 9172 420236 9178
rect 420184 9114 420236 9120
rect 420196 480 420224 9114
rect 418958 354 419070 480
rect 418540 326 419070 354
rect 417854 -960 417966 326
rect 418958 -960 419070 326
rect 420154 -960 420266 480
rect 420932 354 420960 16186
rect 422588 480 422616 16546
rect 423692 3398 423720 29543
rect 425072 16574 425100 31146
rect 445758 27024 445814 27033
rect 445758 26959 445814 26968
rect 440332 23044 440384 23050
rect 440332 22986 440384 22992
rect 426438 21448 426494 21457
rect 426438 21383 426494 21392
rect 426452 16574 426480 21383
rect 429200 20052 429252 20058
rect 429200 19994 429252 20000
rect 425072 16546 425744 16574
rect 426452 16546 426848 16574
rect 423770 4992 423826 5001
rect 423770 4927 423826 4936
rect 423680 3392 423732 3398
rect 423680 3334 423732 3340
rect 423784 480 423812 4927
rect 424968 3392 425020 3398
rect 424968 3334 425020 3340
rect 424980 480 425008 3334
rect 421350 354 421462 480
rect 420932 326 421462 354
rect 421350 -960 421462 326
rect 422546 -960 422658 480
rect 423742 -960 423854 480
rect 424938 -960 425050 480
rect 425716 354 425744 16546
rect 426134 354 426246 480
rect 425716 326 426246 354
rect 426820 354 426848 16546
rect 428462 15872 428518 15881
rect 428462 15807 428518 15816
rect 428476 480 428504 15807
rect 427238 354 427350 480
rect 426820 326 427350 354
rect 426134 -960 426246 326
rect 427238 -960 427350 326
rect 428434 -960 428546 480
rect 429212 354 429240 19994
rect 436100 18692 436152 18698
rect 436100 18634 436152 18640
rect 436112 16574 436140 18634
rect 436112 16546 436784 16574
rect 432052 16176 432104 16182
rect 432052 16118 432104 16124
rect 430856 9444 430908 9450
rect 430856 9386 430908 9392
rect 430868 480 430896 9386
rect 432064 480 432092 16118
rect 435088 16108 435140 16114
rect 435088 16050 435140 16056
rect 434444 9376 434496 9382
rect 434444 9318 434496 9324
rect 433248 3800 433300 3806
rect 433248 3742 433300 3748
rect 433260 480 433288 3742
rect 434456 480 434484 9318
rect 429630 354 429742 480
rect 429212 326 429742 354
rect 429630 -960 429742 326
rect 430826 -960 430938 480
rect 432022 -960 432134 480
rect 433218 -960 433330 480
rect 434414 -960 434526 480
rect 435100 354 435128 16050
rect 436756 480 436784 16546
rect 439136 16040 439188 16046
rect 439136 15982 439188 15988
rect 437940 6316 437992 6322
rect 437940 6258 437992 6264
rect 437952 480 437980 6258
rect 439148 480 439176 15982
rect 440240 4072 440292 4078
rect 440240 4014 440292 4020
rect 440252 2122 440280 4014
rect 440344 3398 440372 22986
rect 441620 21548 441672 21554
rect 441620 21490 441672 21496
rect 441632 16574 441660 21490
rect 442998 19952 443054 19961
rect 442998 19887 443054 19896
rect 443012 16574 443040 19887
rect 441632 16546 442672 16574
rect 443012 16546 443408 16574
rect 440332 3392 440384 3398
rect 440332 3334 440384 3340
rect 441528 3392 441580 3398
rect 441528 3334 441580 3340
rect 440252 2094 440372 2122
rect 440344 480 440372 2094
rect 441540 480 441568 3334
rect 442644 480 442672 16546
rect 435518 354 435630 480
rect 435100 326 435630 354
rect 435518 -960 435630 326
rect 436714 -960 436826 480
rect 437910 -960 438022 480
rect 439106 -960 439218 480
rect 440302 -960 440414 480
rect 441498 -960 441610 480
rect 442602 -960 442714 480
rect 443380 354 443408 16546
rect 445022 9072 445078 9081
rect 445022 9007 445078 9016
rect 445036 480 445064 9007
rect 443798 354 443910 480
rect 443380 326 443910 354
rect 443798 -960 443910 326
rect 444994 -960 445106 480
rect 445772 354 445800 26959
rect 447416 14884 447468 14890
rect 447416 14826 447468 14832
rect 447428 480 447456 14826
rect 448612 12232 448664 12238
rect 448612 12174 448664 12180
rect 448520 4004 448572 4010
rect 448520 3946 448572 3952
rect 448532 1986 448560 3946
rect 448624 3398 448652 12174
rect 450556 3670 450584 36994
rect 454040 20324 454092 20330
rect 454040 20266 454092 20272
rect 453304 14816 453356 14822
rect 453304 14758 453356 14764
rect 451648 12164 451700 12170
rect 451648 12106 451700 12112
rect 450084 3664 450136 3670
rect 450084 3606 450136 3612
rect 450544 3664 450596 3670
rect 450544 3606 450596 3612
rect 448612 3392 448664 3398
rect 448612 3334 448664 3340
rect 449808 3392 449860 3398
rect 449808 3334 449860 3340
rect 448532 1958 448652 1986
rect 448624 480 448652 1958
rect 449820 480 449848 3334
rect 450096 2854 450124 3606
rect 450084 2848 450136 2854
rect 450084 2790 450136 2796
rect 450912 2848 450964 2854
rect 450912 2790 450964 2796
rect 450924 480 450952 2790
rect 446190 354 446302 480
rect 445772 326 446302 354
rect 446190 -960 446302 326
rect 447386 -960 447498 480
rect 448582 -960 448694 480
rect 449778 -960 449890 480
rect 450882 -960 450994 480
rect 451660 354 451688 12106
rect 453316 480 453344 14758
rect 452078 354 452190 480
rect 451660 326 452190 354
rect 452078 -960 452190 326
rect 453274 -960 453386 480
rect 454052 354 454080 20266
rect 456800 19984 456852 19990
rect 456800 19926 456852 19932
rect 455696 12096 455748 12102
rect 455696 12038 455748 12044
rect 455708 480 455736 12038
rect 456812 3398 456840 19926
rect 456892 14748 456944 14754
rect 456892 14690 456944 14696
rect 456800 3392 456852 3398
rect 456800 3334 456852 3340
rect 456904 480 456932 14690
rect 462318 12064 462374 12073
rect 459192 12028 459244 12034
rect 462318 11999 462374 12008
rect 459192 11970 459244 11976
rect 458088 3392 458140 3398
rect 458088 3334 458140 3340
rect 458100 480 458128 3334
rect 459204 480 459232 11970
rect 460388 9104 460440 9110
rect 460388 9046 460440 9052
rect 460400 480 460428 9046
rect 461584 3936 461636 3942
rect 461584 3878 461636 3884
rect 461596 480 461624 3878
rect 454470 354 454582 480
rect 454052 326 454582 354
rect 454470 -960 454582 326
rect 455666 -960 455778 480
rect 456862 -960 456974 480
rect 458058 -960 458170 480
rect 459162 -960 459274 480
rect 460358 -960 460470 480
rect 461554 -960 461666 480
rect 462332 354 462360 11999
rect 462976 4010 463004 38150
rect 474740 38140 474792 38146
rect 474740 38082 474792 38088
rect 471980 21616 472032 21622
rect 471980 21558 472032 21564
rect 468484 17876 468536 17882
rect 468484 17818 468536 17824
rect 466460 17808 466512 17814
rect 466460 17750 466512 17756
rect 463698 17504 463754 17513
rect 463698 17439 463754 17448
rect 463712 16574 463740 17439
rect 466472 16574 466500 17750
rect 463712 16546 464016 16574
rect 466472 16546 467512 16574
rect 462964 4004 463016 4010
rect 462964 3946 463016 3952
rect 463988 480 464016 16546
rect 465172 13252 465224 13258
rect 465172 13194 465224 13200
rect 465184 480 465212 13194
rect 465816 11960 465868 11966
rect 465816 11902 465868 11908
rect 462750 354 462862 480
rect 462332 326 462862 354
rect 462750 -960 462862 326
rect 463946 -960 464058 480
rect 465142 -960 465254 480
rect 465828 354 465856 11902
rect 467484 480 467512 16546
rect 468496 3942 468524 17818
rect 470600 17740 470652 17746
rect 470600 17682 470652 17688
rect 469864 14680 469916 14686
rect 469864 14622 469916 14628
rect 468484 3936 468536 3942
rect 468484 3878 468536 3884
rect 468666 3360 468722 3369
rect 468666 3295 468722 3304
rect 468680 480 468708 3295
rect 469876 480 469904 14622
rect 466246 354 466358 480
rect 465828 326 466358 354
rect 466246 -960 466358 326
rect 467442 -960 467554 480
rect 468638 -960 468750 480
rect 469834 -960 469946 480
rect 470612 354 470640 17682
rect 471992 16574 472020 21558
rect 473360 17672 473412 17678
rect 473360 17614 473412 17620
rect 471992 16546 472296 16574
rect 472268 480 472296 16546
rect 473372 3534 473400 17614
rect 474752 16574 474780 38082
rect 505100 38072 505152 38078
rect 505100 38014 505152 38020
rect 479524 36984 479576 36990
rect 479524 36926 479576 36932
rect 477498 17368 477554 17377
rect 477498 17303 477554 17312
rect 477512 16574 477540 17303
rect 474752 16546 475792 16574
rect 477512 16546 478184 16574
rect 473452 14612 473504 14618
rect 473452 14554 473504 14560
rect 473360 3528 473412 3534
rect 473360 3470 473412 3476
rect 473464 480 473492 14554
rect 474188 3528 474240 3534
rect 474188 3470 474240 3476
rect 471030 354 471142 480
rect 470612 326 471142 354
rect 471030 -960 471142 326
rect 472226 -960 472338 480
rect 473422 -960 473534 480
rect 474200 354 474228 3470
rect 475764 480 475792 16546
rect 476488 14544 476540 14550
rect 476488 14486 476540 14492
rect 474526 354 474638 480
rect 474200 326 474638 354
rect 474526 -960 474638 326
rect 475722 -960 475834 480
rect 476500 354 476528 14486
rect 478156 480 478184 16546
rect 479536 3806 479564 36926
rect 489920 35352 489972 35358
rect 489920 35294 489972 35300
rect 498198 35320 498254 35329
rect 487804 31136 487856 31142
rect 487804 31078 487856 31084
rect 486424 10396 486476 10402
rect 486424 10338 486476 10344
rect 482836 9036 482888 9042
rect 482836 8978 482888 8984
rect 481730 6216 481786 6225
rect 481730 6151 481786 6160
rect 480536 3868 480588 3874
rect 480536 3810 480588 3816
rect 479524 3800 479576 3806
rect 479524 3742 479576 3748
rect 479340 3392 479392 3398
rect 479340 3334 479392 3340
rect 479352 480 479380 3334
rect 480548 480 480576 3810
rect 481744 480 481772 6151
rect 482848 480 482876 8978
rect 485228 8968 485280 8974
rect 485228 8910 485280 8916
rect 484032 3732 484084 3738
rect 484032 3674 484084 3680
rect 484044 480 484072 3674
rect 485240 480 485268 8910
rect 486436 480 486464 10338
rect 487620 4004 487672 4010
rect 487620 3946 487672 3952
rect 487632 480 487660 3946
rect 487816 3534 487844 31078
rect 488540 24268 488592 24274
rect 488540 24210 488592 24216
rect 488552 16574 488580 24210
rect 488552 16546 488856 16574
rect 487804 3528 487856 3534
rect 487804 3470 487856 3476
rect 488828 480 488856 16546
rect 489932 3398 489960 35294
rect 494060 35284 494112 35290
rect 498198 35255 498254 35264
rect 494060 35226 494112 35232
rect 494072 16574 494100 35226
rect 496818 24304 496874 24313
rect 496818 24239 496874 24248
rect 496832 16574 496860 24239
rect 494072 16546 494744 16574
rect 496832 16546 497136 16574
rect 490012 15972 490064 15978
rect 490012 15914 490064 15920
rect 489920 3392 489972 3398
rect 489920 3334 489972 3340
rect 490024 3210 490052 15914
rect 493048 11892 493100 11898
rect 493048 11834 493100 11840
rect 492312 4956 492364 4962
rect 492312 4898 492364 4904
rect 490748 3392 490800 3398
rect 490748 3334 490800 3340
rect 489932 3182 490052 3210
rect 489932 480 489960 3182
rect 476918 354 477030 480
rect 476500 326 477030 354
rect 476918 -960 477030 326
rect 478114 -960 478226 480
rect 479310 -960 479422 480
rect 480506 -960 480618 480
rect 481702 -960 481814 480
rect 482806 -960 482918 480
rect 484002 -960 484114 480
rect 485198 -960 485310 480
rect 486394 -960 486506 480
rect 487590 -960 487702 480
rect 488786 -960 488898 480
rect 489890 -960 490002 480
rect 490760 354 490788 3334
rect 492324 480 492352 4898
rect 491086 354 491198 480
rect 490760 326 491198 354
rect 491086 -960 491198 326
rect 492282 -960 492394 480
rect 493060 354 493088 11834
rect 494716 480 494744 16546
rect 495438 10296 495494 10305
rect 495438 10231 495494 10240
rect 493478 354 493590 480
rect 493060 326 493590 354
rect 493478 -960 493590 326
rect 494674 -960 494786 480
rect 495452 354 495480 10231
rect 497108 480 497136 16546
rect 498212 480 498240 35255
rect 498290 26888 498346 26897
rect 498290 26823 498346 26832
rect 498304 16574 498332 26823
rect 503720 22976 503772 22982
rect 503720 22918 503772 22924
rect 498304 16546 498976 16574
rect 495870 354 495982 480
rect 495452 326 495982 354
rect 495870 -960 495982 326
rect 497066 -960 497178 480
rect 498170 -960 498282 480
rect 498948 354 498976 16546
rect 500592 13184 500644 13190
rect 500592 13126 500644 13132
rect 500604 480 500632 13126
rect 502984 6248 503036 6254
rect 502984 6190 503036 6196
rect 501788 3596 501840 3602
rect 501788 3538 501840 3544
rect 501800 480 501828 3538
rect 502996 480 503024 6190
rect 499366 354 499478 480
rect 498948 326 499478 354
rect 499366 -960 499478 326
rect 500562 -960 500674 480
rect 501758 -960 501870 480
rect 502954 -960 503066 480
rect 503732 354 503760 22918
rect 505112 16574 505140 38014
rect 507860 38004 507912 38010
rect 507860 37946 507912 37952
rect 506480 22908 506532 22914
rect 506480 22850 506532 22856
rect 505112 16546 505416 16574
rect 505388 480 505416 16546
rect 506492 480 506520 22850
rect 507872 16574 507900 37946
rect 539600 37936 539652 37942
rect 539600 37878 539652 37884
rect 514758 33960 514814 33969
rect 514758 33895 514814 33904
rect 512000 32496 512052 32502
rect 512000 32438 512052 32444
rect 507872 16546 508912 16574
rect 507216 15904 507268 15910
rect 507216 15846 507268 15852
rect 504150 354 504262 480
rect 503732 326 504262 354
rect 504150 -960 504262 326
rect 505346 -960 505458 480
rect 506450 -960 506562 480
rect 507228 354 507256 15846
rect 508884 480 508912 16546
rect 510068 7676 510120 7682
rect 510068 7618 510120 7624
rect 510080 480 510108 7618
rect 511264 3936 511316 3942
rect 511264 3878 511316 3884
rect 511276 480 511304 3878
rect 507646 354 507758 480
rect 507228 326 507758 354
rect 507646 -960 507758 326
rect 508842 -960 508954 480
rect 510038 -960 510150 480
rect 511234 -960 511346 480
rect 512012 354 512040 32438
rect 513378 28384 513434 28393
rect 513378 28319 513434 28328
rect 512430 354 512542 480
rect 512012 326 512542 354
rect 513392 354 513420 28319
rect 514772 3602 514800 33895
rect 532698 33824 532754 33833
rect 532698 33759 532754 33768
rect 529940 31068 529992 31074
rect 529940 31010 529992 31016
rect 516138 28248 516194 28257
rect 516138 28183 516194 28192
rect 514850 17232 514906 17241
rect 514850 17167 514906 17176
rect 514760 3596 514812 3602
rect 514760 3538 514812 3544
rect 514864 3482 514892 17167
rect 516152 16574 516180 28183
rect 517520 22840 517572 22846
rect 517520 22782 517572 22788
rect 517532 16574 517560 22782
rect 520280 21480 520332 21486
rect 520280 21422 520332 21428
rect 516152 16546 517192 16574
rect 517532 16546 517928 16574
rect 515588 3596 515640 3602
rect 515588 3538 515640 3544
rect 514772 3454 514892 3482
rect 514772 480 514800 3454
rect 513534 354 513646 480
rect 513392 326 513646 354
rect 512430 -960 512542 326
rect 513534 -960 513646 326
rect 514730 -960 514842 480
rect 515600 354 515628 3538
rect 517164 480 517192 16546
rect 515926 354 516038 480
rect 515600 326 516038 354
rect 515926 -960 516038 326
rect 517122 -960 517234 480
rect 517900 354 517928 16546
rect 519542 3496 519598 3505
rect 519542 3431 519598 3440
rect 519556 480 519584 3431
rect 518318 354 518430 480
rect 517900 326 518430 354
rect 518318 -960 518430 326
rect 519514 -960 519626 480
rect 520292 354 520320 21422
rect 521660 17604 521712 17610
rect 521660 17546 521712 17552
rect 520710 354 520822 480
rect 520292 326 520822 354
rect 521672 354 521700 17546
rect 524420 17536 524472 17542
rect 524420 17478 524472 17484
rect 524432 16574 524460 17478
rect 528560 17468 528612 17474
rect 528560 17410 528612 17416
rect 524432 16546 525472 16574
rect 523776 11824 523828 11830
rect 523776 11766 523828 11772
rect 523040 3664 523092 3670
rect 523040 3606 523092 3612
rect 523052 480 523080 3606
rect 521814 354 521926 480
rect 521672 326 521926 354
rect 520710 -960 520822 326
rect 521814 -960 521926 326
rect 523010 -960 523122 480
rect 523788 354 523816 11766
rect 525444 480 525472 16546
rect 527824 11756 527876 11762
rect 527824 11698 527876 11704
rect 526628 3800 526680 3806
rect 526628 3742 526680 3748
rect 526640 480 526668 3742
rect 527836 480 527864 11698
rect 524206 354 524318 480
rect 523788 326 524318 354
rect 524206 -960 524318 326
rect 525402 -960 525514 480
rect 526598 -960 526710 480
rect 527794 -960 527906 480
rect 528572 354 528600 17410
rect 528990 354 529102 480
rect 528572 326 529102 354
rect 529952 354 529980 31010
rect 531318 30968 531374 30977
rect 531318 30903 531374 30912
rect 531332 3602 531360 30903
rect 532712 16574 532740 33759
rect 538220 29776 538272 29782
rect 538220 29718 538272 29724
rect 536840 18624 536892 18630
rect 536840 18566 536892 18572
rect 535460 17400 535512 17406
rect 535460 17342 535512 17348
rect 535472 16574 535500 17342
rect 536852 16574 536880 18566
rect 532712 16546 533752 16574
rect 535472 16546 536144 16574
rect 536852 16546 537248 16574
rect 531410 11928 531466 11937
rect 531410 11863 531466 11872
rect 531320 3596 531372 3602
rect 531320 3538 531372 3544
rect 531424 3482 531452 11863
rect 532148 3596 532200 3602
rect 532148 3538 532200 3544
rect 531332 3454 531452 3482
rect 531332 480 531360 3454
rect 530094 354 530206 480
rect 529952 326 530206 354
rect 528990 -960 529102 326
rect 530094 -960 530206 326
rect 531290 -960 531402 480
rect 532160 354 532188 3538
rect 533724 480 533752 16546
rect 534446 11792 534502 11801
rect 534446 11727 534502 11736
rect 532486 354 532598 480
rect 532160 326 532598 354
rect 532486 -960 532598 326
rect 533682 -960 533794 480
rect 534460 354 534488 11727
rect 536116 480 536144 16546
rect 537220 480 537248 16546
rect 534878 354 534990 480
rect 534460 326 534990 354
rect 534878 -960 534990 326
rect 536074 -960 536186 480
rect 537178 -960 537290 480
rect 538232 354 538260 29718
rect 539612 3602 539640 37878
rect 543740 36916 543792 36922
rect 543740 36858 543792 36864
rect 540980 21412 541032 21418
rect 540980 21354 541032 21360
rect 539692 17332 539744 17338
rect 539692 17274 539744 17280
rect 539600 3596 539652 3602
rect 539600 3538 539652 3544
rect 539704 3482 539732 17274
rect 540992 16574 541020 21354
rect 543752 16574 543780 36858
rect 547880 36848 547932 36854
rect 547880 36790 547932 36796
rect 545120 25560 545172 25566
rect 545120 25502 545172 25508
rect 545132 16574 545160 25502
rect 546500 17264 546552 17270
rect 546500 17206 546552 17212
rect 540992 16546 542032 16574
rect 543752 16546 544424 16574
rect 545132 16546 545528 16574
rect 540428 3596 540480 3602
rect 540428 3538 540480 3544
rect 539612 3454 539732 3482
rect 539612 480 539640 3454
rect 538374 354 538486 480
rect 538232 326 538486 354
rect 538374 -960 538486 326
rect 539570 -960 539682 480
rect 540440 354 540468 3538
rect 542004 480 542032 16546
rect 542728 14476 542780 14482
rect 542728 14418 542780 14424
rect 540766 354 540878 480
rect 540440 326 540878 354
rect 540766 -960 540878 326
rect 541962 -960 542074 480
rect 542740 354 542768 14418
rect 544396 480 544424 16546
rect 545500 480 545528 16546
rect 543158 354 543270 480
rect 542740 326 543270 354
rect 543158 -960 543270 326
rect 544354 -960 544466 480
rect 545458 -960 545570 480
rect 546512 354 546540 17206
rect 547892 480 547920 36790
rect 554780 36780 554832 36786
rect 554780 36722 554832 36728
rect 549258 35184 549314 35193
rect 549258 35119 549314 35128
rect 549272 16574 549300 35119
rect 550638 32600 550694 32609
rect 550638 32535 550694 32544
rect 550652 16574 550680 32535
rect 552018 32464 552074 32473
rect 552018 32399 552074 32408
rect 552032 16574 552060 32399
rect 549272 16546 550312 16574
rect 550652 16546 551048 16574
rect 552032 16546 552704 16574
rect 549074 8936 549130 8945
rect 549074 8871 549130 8880
rect 549088 480 549116 8871
rect 550284 480 550312 16546
rect 546654 354 546766 480
rect 546512 326 546766 354
rect 546654 -960 546766 326
rect 547850 -960 547962 480
rect 549046 -960 549158 480
rect 550242 -960 550354 480
rect 551020 354 551048 16546
rect 552676 480 552704 16546
rect 553768 6180 553820 6186
rect 553768 6122 553820 6128
rect 553780 480 553808 6122
rect 551438 354 551550 480
rect 551020 326 551550 354
rect 551438 -960 551550 326
rect 552634 -960 552746 480
rect 553738 -960 553850 480
rect 554792 354 554820 36722
rect 557540 36712 557592 36718
rect 557540 36654 557592 36660
rect 556252 24200 556304 24206
rect 556252 24142 556304 24148
rect 556264 16574 556292 24142
rect 557552 16574 557580 36654
rect 580356 36644 580408 36650
rect 580356 36586 580408 36592
rect 580264 36576 580316 36582
rect 580264 36518 580316 36524
rect 561680 35216 561732 35222
rect 561680 35158 561732 35164
rect 558920 28280 558972 28286
rect 558920 28222 558972 28228
rect 558932 16574 558960 28222
rect 560300 26988 560352 26994
rect 560300 26930 560352 26936
rect 560312 16574 560340 26930
rect 561692 16574 561720 35158
rect 564440 33788 564492 33794
rect 564440 33730 564492 33736
rect 563060 24132 563112 24138
rect 563060 24074 563112 24080
rect 556264 16546 556936 16574
rect 557552 16546 558592 16574
rect 558932 16546 559328 16574
rect 560312 16546 560432 16574
rect 561692 16546 562088 16574
rect 556160 3528 556212 3534
rect 556160 3470 556212 3476
rect 556172 480 556200 3470
rect 554934 354 555046 480
rect 554792 326 555046 354
rect 554934 -960 555046 326
rect 556130 -960 556242 480
rect 556908 354 556936 16546
rect 558564 480 558592 16546
rect 557326 354 557438 480
rect 556908 326 557438 354
rect 557326 -960 557438 326
rect 558522 -960 558634 480
rect 559300 354 559328 16546
rect 559718 354 559830 480
rect 559300 326 559830 354
rect 560404 354 560432 16546
rect 562060 480 562088 16546
rect 560822 354 560934 480
rect 560404 326 560934 354
rect 559718 -960 559830 326
rect 560822 -960 560934 326
rect 562018 -960 562130 480
rect 563072 354 563100 24074
rect 564452 480 564480 33730
rect 576860 32428 576912 32434
rect 576860 32370 576912 32376
rect 572720 29708 572772 29714
rect 572720 29650 572772 29656
rect 569958 25664 570014 25673
rect 569958 25599 570014 25608
rect 568578 24168 568634 24177
rect 568578 24103 568634 24112
rect 564532 22772 564584 22778
rect 564532 22714 564584 22720
rect 564544 16574 564572 22714
rect 568592 16574 568620 24103
rect 569972 16574 570000 25599
rect 564544 16546 565216 16574
rect 568592 16546 568712 16574
rect 569972 16546 570368 16574
rect 563214 354 563326 480
rect 563072 326 563326 354
rect 563214 -960 563326 326
rect 564410 -960 564522 480
rect 565188 354 565216 16546
rect 567566 11656 567622 11665
rect 567566 11591 567622 11600
rect 566830 4856 566886 4865
rect 566830 4791 566886 4800
rect 566844 480 566872 4791
rect 565606 354 565718 480
rect 565188 326 565718 354
rect 565606 -960 565718 326
rect 566802 -960 566914 480
rect 567580 354 567608 11591
rect 567998 354 568110 480
rect 567580 326 568110 354
rect 568684 354 568712 16546
rect 570340 480 570368 16546
rect 571524 7608 571576 7614
rect 571524 7550 571576 7556
rect 571536 480 571564 7550
rect 572732 3534 572760 29650
rect 572812 26920 572864 26926
rect 572812 26862 572864 26868
rect 572720 3528 572772 3534
rect 572720 3470 572772 3476
rect 572824 3346 572852 26862
rect 576872 16574 576900 32370
rect 579620 29640 579672 29646
rect 579620 29582 579672 29588
rect 576872 16546 576992 16574
rect 575112 10328 575164 10334
rect 575112 10270 575164 10276
rect 573548 3528 573600 3534
rect 573548 3470 573600 3476
rect 572732 3318 572852 3346
rect 572732 480 572760 3318
rect 569102 354 569214 480
rect 568684 326 569214 354
rect 567998 -960 568110 326
rect 569102 -960 569214 326
rect 570298 -960 570410 480
rect 571494 -960 571606 480
rect 572690 -960 572802 480
rect 573560 354 573588 3470
rect 575124 480 575152 10270
rect 576308 4820 576360 4826
rect 576308 4762 576360 4768
rect 576320 480 576348 4762
rect 573886 354 573998 480
rect 573560 326 573998 354
rect 573886 -960 573998 326
rect 575082 -960 575194 480
rect 576278 -960 576390 480
rect 576964 354 576992 16546
rect 578608 13116 578660 13122
rect 578608 13058 578660 13064
rect 578620 480 578648 13058
rect 577382 354 577494 480
rect 576964 326 577494 354
rect 577382 -960 577494 326
rect 578578 -960 578690 480
rect 579632 354 579660 29582
rect 580276 19825 580304 36518
rect 580368 33153 580396 36586
rect 580354 33144 580410 33153
rect 580354 33079 580410 33088
rect 580998 25528 581054 25537
rect 580998 25463 581054 25472
rect 580262 19816 580318 19825
rect 580262 19751 580318 19760
rect 580172 6860 580224 6866
rect 580172 6802 580224 6808
rect 580184 6633 580212 6802
rect 580170 6624 580226 6633
rect 580170 6559 580226 6568
rect 581012 480 581040 25463
rect 581090 21312 581146 21321
rect 581090 21247 581146 21256
rect 581104 16574 581132 21247
rect 581104 16546 581776 16574
rect 579774 354 579886 480
rect 579632 326 579886 354
rect 579774 -960 579886 326
rect 580970 -960 581082 480
rect 581748 354 581776 16546
rect 583392 3460 583444 3466
rect 583392 3402 583444 3408
rect 583404 480 583432 3402
rect 582166 354 582278 480
rect 581748 326 582278 354
rect 582166 -960 582278 326
rect 583362 -960 583474 480
<< via2 >>
rect 3422 684256 3478 684312
rect 3514 671200 3570 671256
rect 3422 658144 3478 658200
rect 3422 632068 3424 632088
rect 3424 632068 3476 632088
rect 3476 632068 3478 632088
rect 3422 632032 3478 632068
rect 3146 619112 3202 619168
rect 3238 606056 3294 606112
rect 3330 579944 3386 580000
rect 3422 566888 3478 566944
rect 3422 553832 3478 553888
rect 2962 527856 3018 527912
rect 3330 423544 3386 423600
rect 3330 410488 3386 410544
rect 3330 397468 3332 397488
rect 3332 397468 3384 397488
rect 3384 397468 3386 397488
rect 3330 397432 3386 397468
rect 3330 371320 3386 371376
rect 2962 358400 3018 358456
rect 3054 345344 3110 345400
rect 3514 514820 3570 514856
rect 3514 514800 3516 514820
rect 3516 514800 3568 514820
rect 3568 514800 3570 514820
rect 3514 501744 3570 501800
rect 3606 475632 3662 475688
rect 3698 462576 3754 462632
rect 3790 449520 3846 449576
rect 3422 319232 3478 319288
rect 3238 306176 3294 306232
rect 3422 293120 3478 293176
rect 3054 267144 3110 267200
rect 3330 214920 3386 214976
rect 3238 201864 3294 201920
rect 3330 162832 3386 162888
rect 3514 254088 3570 254144
rect 3514 241032 3570 241088
rect 3606 188808 3662 188864
rect 3422 149776 3478 149832
rect 3422 136720 3478 136776
rect 111890 591640 111946 591696
rect 111798 590960 111854 591016
rect 111890 590280 111946 590336
rect 111798 589600 111854 589656
rect 111798 588920 111854 588976
rect 112258 588240 112314 588296
rect 111798 587560 111854 587616
rect 111798 586200 111854 586256
rect 112718 586880 112774 586936
rect 111982 585520 112038 585576
rect 111890 584840 111946 584896
rect 111798 584160 111854 584216
rect 111798 583480 111854 583536
rect 111890 582800 111946 582856
rect 111798 582120 111854 582176
rect 111982 581440 112038 581496
rect 111890 580760 111946 580816
rect 111798 580080 111854 580136
rect 111890 579400 111946 579456
rect 111798 578720 111854 578776
rect 111798 578040 111854 578096
rect 112442 577360 112498 577416
rect 111890 576680 111946 576736
rect 111798 576000 111854 576056
rect 111890 575320 111946 575376
rect 111798 574640 111854 574696
rect 111890 573960 111946 574016
rect 111798 573280 111854 573336
rect 111890 572600 111946 572656
rect 111798 571920 111854 571976
rect 111982 571240 112038 571296
rect 111798 570560 111854 570616
rect 111890 569880 111946 569936
rect 111798 569200 111854 569256
rect 111982 568520 112038 568576
rect 111798 567196 111800 567216
rect 111800 567196 111852 567216
rect 111852 567196 111854 567216
rect 111798 567160 111854 567196
rect 111890 566480 111946 566536
rect 111798 565800 111854 565856
rect 111890 565120 111946 565176
rect 111798 564476 111800 564496
rect 111800 564476 111852 564496
rect 111852 564476 111854 564496
rect 111798 564440 111854 564476
rect 111798 563100 111854 563136
rect 111798 563080 111800 563100
rect 111800 563080 111852 563100
rect 111852 563080 111854 563100
rect 112350 567840 112406 567896
rect 112626 562400 112682 562456
rect 111798 561740 111854 561776
rect 111798 561720 111800 561740
rect 111800 561720 111852 561740
rect 111852 561720 111854 561740
rect 112442 561040 112498 561096
rect 111798 560360 111854 560416
rect 111890 559680 111946 559736
rect 111798 559020 111854 559056
rect 111798 559000 111800 559020
rect 111800 559000 111852 559020
rect 111852 559000 111854 559020
rect 111890 558320 111946 558376
rect 111798 557660 111854 557696
rect 111798 557640 111800 557660
rect 111800 557640 111852 557660
rect 111852 557640 111854 557660
rect 111798 556960 111854 557016
rect 111982 556280 112038 556336
rect 111890 555600 111946 555656
rect 111798 554940 111854 554976
rect 111798 554920 111800 554940
rect 111800 554920 111852 554940
rect 111852 554920 111854 554940
rect 112074 554240 112130 554296
rect 111798 553560 111854 553616
rect 111890 552880 111946 552936
rect 111798 552200 111854 552256
rect 111890 551520 111946 551576
rect 111798 550840 111854 550896
rect 111890 550160 111946 550216
rect 111798 549480 111854 549536
rect 111890 548800 111946 548856
rect 111798 548140 111854 548176
rect 111798 548120 111800 548140
rect 111800 548120 111852 548140
rect 111852 548120 111854 548140
rect 111798 546760 111854 546816
rect 111890 546080 111946 546136
rect 111798 545400 111854 545456
rect 111798 544040 111854 544096
rect 111890 543360 111946 543416
rect 111798 542680 111854 542736
rect 111798 542000 111854 542056
rect 112350 540640 112406 540696
rect 111798 539960 111854 540016
rect 111890 539280 111946 539336
rect 111798 538600 111854 538656
rect 111890 537920 111946 537976
rect 111798 537240 111854 537296
rect 111890 536560 111946 536616
rect 111798 535880 111854 535936
rect 111798 535200 111854 535256
rect 111890 534520 111946 534576
rect 112258 532480 112314 532536
rect 112994 563760 113050 563816
rect 112810 547440 112866 547496
rect 112718 533840 112774 533896
rect 112626 530440 112682 530496
rect 112350 529760 112406 529816
rect 111798 528400 111854 528456
rect 112258 527720 112314 527776
rect 112350 527040 112406 527096
rect 112074 525680 112130 525736
rect 111890 524320 111946 524376
rect 111798 523640 111854 523696
rect 111890 522960 111946 523016
rect 111798 522280 111854 522336
rect 111890 521600 111946 521656
rect 111798 520920 111854 520976
rect 111798 520240 111854 520296
rect 112350 519560 112406 519616
rect 112258 518880 112314 518936
rect 111798 517540 111854 517576
rect 111798 517520 111800 517540
rect 111800 517520 111852 517540
rect 111852 517520 111854 517540
rect 111890 516840 111946 516896
rect 111798 516180 111854 516216
rect 111798 516160 111800 516180
rect 111800 516160 111852 516180
rect 111852 516160 111854 516180
rect 111890 515480 111946 515536
rect 111798 514836 111800 514856
rect 111800 514836 111852 514856
rect 111852 514836 111854 514856
rect 111798 514800 111854 514836
rect 111890 514120 111946 514176
rect 111798 513460 111854 513496
rect 111798 513440 111800 513460
rect 111800 513440 111852 513460
rect 111852 513440 111854 513460
rect 111982 512760 112038 512816
rect 111798 512080 111854 512136
rect 111890 511400 111946 511456
rect 111798 510720 111854 510776
rect 111798 509360 111854 509416
rect 111890 508680 111946 508736
rect 111798 508000 111854 508056
rect 111798 507320 111854 507376
rect 111890 506640 111946 506696
rect 111798 505960 111854 506016
rect 112350 505280 112406 505336
rect 111890 504600 111946 504656
rect 111798 503940 111854 503976
rect 111798 503920 111800 503940
rect 111800 503920 111852 503940
rect 111852 503920 111854 503940
rect 111890 503240 111946 503296
rect 111798 502560 111854 502616
rect 111798 501880 111854 501936
rect 111890 501200 111946 501256
rect 111798 499840 111854 499896
rect 111982 500520 112038 500576
rect 111982 499160 112038 499216
rect 111798 498480 111854 498536
rect 111890 497800 111946 497856
rect 111798 497120 111854 497176
rect 111890 496440 111946 496496
rect 111798 495780 111854 495816
rect 111798 495760 111800 495780
rect 111800 495760 111852 495780
rect 111852 495760 111854 495780
rect 111798 495100 111854 495136
rect 111798 495080 111800 495100
rect 111800 495080 111852 495100
rect 111852 495080 111854 495100
rect 111798 494400 111854 494456
rect 111798 493720 111854 493776
rect 111890 492360 111946 492416
rect 111798 491680 111854 491736
rect 111890 491000 111946 491056
rect 111798 490320 111854 490376
rect 111890 489640 111946 489696
rect 111798 488960 111854 489016
rect 111890 488280 111946 488336
rect 111798 487600 111854 487656
rect 111890 486920 111946 486976
rect 111798 486240 111854 486296
rect 111798 484880 111854 484936
rect 111890 484200 111946 484256
rect 111798 483520 111854 483576
rect 111890 482840 111946 482896
rect 111798 482160 111854 482216
rect 111890 481480 111946 481536
rect 111798 480800 111854 480856
rect 111890 480120 111946 480176
rect 111798 479440 111854 479496
rect 111890 478760 111946 478816
rect 111798 478080 111854 478136
rect 111798 476720 111854 476776
rect 111890 476040 111946 476096
rect 111798 475360 111854 475416
rect 111798 474680 111854 474736
rect 111890 474000 111946 474056
rect 111798 473320 111854 473376
rect 111890 472640 111946 472696
rect 111798 471960 111854 472016
rect 111890 471280 111946 471336
rect 111798 470620 111854 470656
rect 111798 470600 111800 470620
rect 111800 470600 111852 470620
rect 111852 470600 111854 470620
rect 111798 469920 111854 469976
rect 111798 469260 111854 469296
rect 111798 469240 111800 469260
rect 111800 469240 111852 469260
rect 111852 469240 111854 469260
rect 111890 468560 111946 468616
rect 111798 467916 111800 467936
rect 111800 467916 111852 467936
rect 111852 467916 111854 467936
rect 111798 467880 111854 467916
rect 111890 467200 111946 467256
rect 111798 466540 111854 466576
rect 111798 466520 111800 466540
rect 111800 466520 111852 466540
rect 111852 466520 111854 466540
rect 111890 465840 111946 465896
rect 111798 465160 111854 465216
rect 111890 464480 111946 464536
rect 111798 463820 111854 463856
rect 111798 463800 111800 463820
rect 111800 463800 111852 463820
rect 111852 463800 111854 463820
rect 111890 463120 111946 463176
rect 111798 462460 111854 462496
rect 111798 462440 111800 462460
rect 111800 462440 111852 462460
rect 111852 462440 111854 462460
rect 111890 461760 111946 461816
rect 111798 461080 111854 461136
rect 111798 460400 111854 460456
rect 112350 459720 112406 459776
rect 111890 459040 111946 459096
rect 111798 458360 111854 458416
rect 112258 457680 112314 457736
rect 111798 457000 111854 457056
rect 111890 456320 111946 456376
rect 111798 455640 111854 455696
rect 111798 454960 111854 455016
rect 111798 454280 111854 454336
rect 111890 453600 111946 453656
rect 111798 452920 111854 452976
rect 111890 452240 111946 452296
rect 111798 451560 111854 451616
rect 111890 450880 111946 450936
rect 111798 450200 111854 450256
rect 111890 449520 111946 449576
rect 111798 448840 111854 448896
rect 111798 448160 111854 448216
rect 112718 525000 112774 525056
rect 112902 544720 112958 544776
rect 112810 518200 112866 518256
rect 112902 510040 112958 510096
rect 113086 541320 113142 541376
rect 113086 533160 113142 533216
rect 113086 531800 113142 531856
rect 113086 531120 113142 531176
rect 113086 529080 113142 529136
rect 113086 526360 113142 526416
rect 113086 493040 113142 493096
rect 112994 485560 113050 485616
rect 113086 477400 113142 477456
rect 111798 314200 111854 314256
rect 111798 313112 111854 313168
rect 111890 312704 111946 312760
rect 111798 311772 111854 311808
rect 111798 311752 111800 311772
rect 111800 311752 111852 311772
rect 111852 311752 111854 311772
rect 111890 311344 111946 311400
rect 111798 310428 111800 310448
rect 111800 310428 111852 310448
rect 111852 310428 111854 310448
rect 111798 310392 111854 310428
rect 111890 309984 111946 310040
rect 111798 309068 111800 309088
rect 111800 309068 111852 309088
rect 111852 309068 111854 309088
rect 111798 309032 111854 309068
rect 111890 308624 111946 308680
rect 111798 307708 111800 307728
rect 111800 307708 111852 307728
rect 111852 307708 111854 307728
rect 111798 307672 111854 307708
rect 111798 307264 111854 307320
rect 111798 306332 111854 306368
rect 111798 306312 111800 306332
rect 111800 306312 111852 306332
rect 111852 306312 111854 306332
rect 111890 305904 111946 305960
rect 111798 304852 111800 304872
rect 111800 304852 111852 304872
rect 111852 304852 111854 304872
rect 111798 304816 111854 304852
rect 111890 304544 111946 304600
rect 111798 303492 111800 303512
rect 111800 303492 111852 303512
rect 111852 303492 111854 303512
rect 111798 303456 111854 303492
rect 111890 303184 111946 303240
rect 111798 302132 111800 302152
rect 111800 302132 111852 302152
rect 111852 302132 111854 302152
rect 111798 302096 111854 302132
rect 111890 301824 111946 301880
rect 111890 300756 111946 300792
rect 111890 300736 111892 300756
rect 111892 300736 111944 300756
rect 111944 300736 111946 300756
rect 111798 300328 111854 300384
rect 111982 299920 112038 299976
rect 111798 298968 111854 299024
rect 111798 298424 111854 298480
rect 111798 297608 111854 297664
rect 111890 297200 111946 297256
rect 111798 296384 111854 296440
rect 111890 295840 111946 295896
rect 111798 294888 111854 294944
rect 111890 294480 111946 294536
rect 111798 293664 111854 293720
rect 111890 293120 111946 293176
rect 111798 292168 111854 292224
rect 111890 291760 111946 291816
rect 111798 290808 111854 290864
rect 111890 290400 111946 290456
rect 111798 289448 111854 289504
rect 111890 289040 111946 289096
rect 111798 288088 111854 288144
rect 111890 287680 111946 287736
rect 111798 286728 111854 286784
rect 111890 286320 111946 286376
rect 111798 285368 111854 285424
rect 111890 284960 111946 285016
rect 111798 284008 111854 284064
rect 111890 283600 111946 283656
rect 112074 282784 112130 282840
rect 111798 282240 111854 282296
rect 111798 281288 111854 281344
rect 111890 280880 111946 280936
rect 111798 279928 111854 279984
rect 111890 279520 111946 279576
rect 111798 278432 111854 278488
rect 111890 278160 111946 278216
rect 111798 277208 111854 277264
rect 111890 276800 111946 276856
rect 111798 275848 111854 275904
rect 111890 275440 111946 275496
rect 111798 274352 111854 274408
rect 111890 274080 111946 274136
rect 111798 273028 111800 273048
rect 111800 273028 111852 273048
rect 111852 273028 111854 273048
rect 111798 272992 111854 273028
rect 111890 272720 111946 272776
rect 111798 271632 111854 271688
rect 111890 271360 111946 271416
rect 111798 270272 111854 270328
rect 111890 270000 111946 270056
rect 111798 268948 111800 268968
rect 111800 268948 111852 268968
rect 111852 268948 111854 268968
rect 111798 268912 111854 268948
rect 111890 268640 111946 268696
rect 111798 267552 111854 267608
rect 111890 267144 111946 267200
rect 111798 266228 111800 266248
rect 111800 266228 111852 266248
rect 111852 266228 111854 266248
rect 111798 266192 111854 266228
rect 111890 265920 111946 265976
rect 111798 264852 111854 264888
rect 111798 264832 111800 264852
rect 111800 264832 111852 264852
rect 111852 264832 111854 264852
rect 111890 264424 111946 264480
rect 111798 263492 111854 263528
rect 111798 263472 111800 263492
rect 111800 263472 111852 263492
rect 111852 263472 111854 263492
rect 111890 263064 111946 263120
rect 112166 262112 112222 262168
rect 111798 261704 111854 261760
rect 111798 260788 111800 260808
rect 111800 260788 111852 260808
rect 111852 260788 111854 260808
rect 111798 260752 111854 260788
rect 111890 260344 111946 260400
rect 111798 259292 111800 259312
rect 111800 259292 111852 259312
rect 111852 259292 111854 259312
rect 111798 259256 111854 259292
rect 111890 258984 111946 259040
rect 111798 257932 111800 257952
rect 111800 257932 111852 257952
rect 111852 257932 111854 257952
rect 111798 257896 111854 257932
rect 111890 257624 111946 257680
rect 111798 256264 111854 256320
rect 111798 254904 111854 254960
rect 111798 253852 111800 253872
rect 111800 253852 111852 253872
rect 111852 253852 111854 253872
rect 111798 253816 111854 253852
rect 111890 253544 111946 253600
rect 111798 253000 111854 253056
rect 111798 252184 111854 252240
rect 112258 251640 112314 251696
rect 111798 250824 111854 250880
rect 111890 250280 111946 250336
rect 111798 249464 111854 249520
rect 111798 247968 111854 248024
rect 111890 247560 111946 247616
rect 111798 246608 111854 246664
rect 111890 246200 111946 246256
rect 111798 245248 111854 245304
rect 111890 244840 111946 244896
rect 111798 243888 111854 243944
rect 111798 242528 111854 242584
rect 112350 243480 112406 243536
rect 111982 242120 112038 242176
rect 111890 241440 111946 241496
rect 111798 240760 111854 240816
rect 111798 239808 111854 239864
rect 111890 239400 111946 239456
rect 111798 238448 111854 238504
rect 111890 238040 111946 238096
rect 111798 237088 111854 237144
rect 112350 236680 112406 236736
rect 111798 235728 111854 235784
rect 111890 235320 111946 235376
rect 111798 234368 111854 234424
rect 111890 233960 111946 234016
rect 111798 233144 111854 233200
rect 111798 232464 111854 232520
rect 111798 231240 111854 231296
rect 111798 230288 111854 230344
rect 111890 229880 111946 229936
rect 111798 228928 111854 228984
rect 111890 228520 111946 228576
rect 111798 227568 111854 227624
rect 111890 227160 111946 227216
rect 112350 226208 112406 226264
rect 111798 225664 111854 225720
rect 111798 224712 111854 224768
rect 111890 224440 111946 224496
rect 111798 223352 111854 223408
rect 111890 223080 111946 223136
rect 111798 221992 111854 222048
rect 111890 221584 111946 221640
rect 111798 220632 111854 220688
rect 111890 220224 111946 220280
rect 111798 217948 111800 217968
rect 111800 217948 111852 217968
rect 111852 217948 111854 217968
rect 111798 217912 111854 217948
rect 111890 217640 111946 217696
rect 111798 216144 111854 216200
rect 111798 215228 111800 215248
rect 111800 215228 111852 215248
rect 111852 215228 111854 215248
rect 111798 215192 111854 215228
rect 111890 214784 111946 214840
rect 111798 213868 111800 213888
rect 111800 213868 111852 213888
rect 111852 213868 111854 213888
rect 111798 213832 111854 213868
rect 111890 213424 111946 213480
rect 111798 212492 111854 212528
rect 111798 212472 111800 212492
rect 111800 212472 111852 212492
rect 111852 212472 111854 212492
rect 111890 212064 111946 212120
rect 111798 211132 111854 211168
rect 111798 211112 111800 211132
rect 111800 211112 111852 211132
rect 111852 211112 111854 211132
rect 111890 210704 111946 210760
rect 111798 209616 111854 209672
rect 111798 208256 111854 208312
rect 111798 206932 111800 206952
rect 111800 206932 111852 206952
rect 111852 206932 111854 206952
rect 111798 206896 111854 206932
rect 111890 206624 111946 206680
rect 111982 206080 112038 206136
rect 111798 204992 111854 205048
rect 111890 204720 111946 204776
rect 111798 203632 111854 203688
rect 111890 203360 111946 203416
rect 111798 202544 111854 202600
rect 111890 202000 111946 202056
rect 111798 201048 111854 201104
rect 112994 261024 113050 261080
rect 112994 260480 113050 260536
rect 113086 256536 113142 256592
rect 112994 255176 113050 255232
rect 112810 248920 112866 248976
rect 112902 231784 112958 231840
rect 112626 219272 112682 219328
rect 112810 219000 112866 219056
rect 112902 216552 112958 216608
rect 112442 209344 112498 209400
rect 112350 208120 112406 208176
rect 112074 200640 112130 200696
rect 111798 199688 111854 199744
rect 111890 199280 111946 199336
rect 111798 198328 111854 198384
rect 112258 197240 112314 197296
rect 111798 196560 111854 196616
rect 111798 195608 111854 195664
rect 111890 195200 111946 195256
rect 111798 194248 111854 194304
rect 111890 193704 111946 193760
rect 111798 192888 111854 192944
rect 111890 192480 111946 192536
rect 111798 191528 111854 191584
rect 111798 190848 111854 190904
rect 111798 190168 111854 190224
rect 111890 189760 111946 189816
rect 111798 188808 111854 188864
rect 111890 188400 111946 188456
rect 111798 187448 111854 187504
rect 111890 187040 111946 187096
rect 111798 185680 111854 185736
rect 111798 184592 111854 184648
rect 111890 184320 111946 184376
rect 111798 182960 111854 183016
rect 111798 182008 111854 182064
rect 111798 181464 111854 181520
rect 111798 180512 111854 180568
rect 111890 180240 111946 180296
rect 111798 179152 111854 179208
rect 111890 178880 111946 178936
rect 111798 176432 111854 176488
rect 111890 176160 111946 176216
rect 111982 175208 112038 175264
rect 112902 197920 112958 197976
rect 112534 183504 112590 183560
rect 112902 186224 112958 186280
rect 112718 177928 112774 177984
rect 112810 177520 112866 177576
rect 112442 174800 112498 174856
rect 111798 173712 111854 173768
rect 111890 173304 111946 173360
rect 111798 172080 111854 172136
rect 111798 171012 111854 171048
rect 111798 170992 111800 171012
rect 111800 170992 111852 171012
rect 111852 170992 111854 171012
rect 111890 170584 111946 170640
rect 3422 110608 3478 110664
rect 3422 97552 3478 97608
rect 3422 84632 3478 84688
rect 3514 71576 3570 71632
rect 3606 58520 3662 58576
rect 3698 45464 3754 45520
rect 3790 32408 3846 32464
rect 135258 120808 135314 120864
rect 135442 118224 135498 118280
rect 135258 86844 135260 86864
rect 135260 86844 135312 86864
rect 135312 86844 135314 86864
rect 135258 86808 135314 86844
rect 135810 84768 135866 84824
rect 135350 71612 135352 71632
rect 135352 71612 135404 71632
rect 135404 71612 135406 71632
rect 135350 71576 135406 71612
rect 135718 68856 135774 68912
rect 135626 61512 135682 61568
rect 135258 56380 135260 56400
rect 135260 56380 135312 56400
rect 135312 56380 135314 56400
rect 135258 56344 135314 56380
rect 136546 130464 136602 130520
rect 136546 127880 136602 127936
rect 136546 125432 136602 125488
rect 136178 123528 136234 123584
rect 136546 115504 136602 115560
rect 136546 112784 136602 112840
rect 136546 110200 136602 110256
rect 136546 107480 136602 107536
rect 136546 104796 136548 104816
rect 136548 104796 136600 104816
rect 136600 104796 136602 104816
rect 136546 104760 136602 104796
rect 136178 102856 136234 102912
rect 136178 100136 136234 100192
rect 136546 95104 136602 95160
rect 136086 92420 136088 92440
rect 136088 92420 136140 92440
rect 136140 92420 136142 92440
rect 136086 92384 136142 92420
rect 136546 89528 136602 89584
rect 136546 82220 136548 82240
rect 136548 82220 136600 82240
rect 136600 82220 136602 82240
rect 136546 82184 136602 82220
rect 136086 79600 136142 79656
rect 136546 77052 136548 77072
rect 136548 77052 136600 77072
rect 136600 77052 136602 77072
rect 136546 77016 136602 77052
rect 136546 73772 136602 73808
rect 136546 73752 136548 73772
rect 136548 73752 136600 73772
rect 136600 73752 136602 73772
rect 136086 66172 136088 66192
rect 136088 66172 136140 66192
rect 136140 66172 136142 66192
rect 136086 66136 136142 66172
rect 136546 64132 136548 64152
rect 136548 64132 136600 64152
rect 136600 64132 136602 64152
rect 136546 64096 136602 64132
rect 136546 58964 136548 58984
rect 136548 58964 136600 58984
rect 136600 58964 136602 58984
rect 136546 58928 136602 58964
rect 136546 53488 136602 53544
rect 136730 97688 136786 97744
rect 135350 50940 135352 50960
rect 135352 50940 135404 50960
rect 135404 50940 135406 50960
rect 135350 50904 135406 50940
rect 134614 48320 134670 48376
rect 22742 24792 22798 24848
rect 18602 24112 18658 24168
rect 1398 21256 1454 21312
rect 3422 19352 3478 19408
rect 3606 11600 3662 11656
rect 3422 6432 3478 6488
rect 19338 22616 19394 22672
rect 20718 18536 20774 18592
rect 23018 8880 23074 8936
rect 36726 10240 36782 10296
rect 38382 6160 38438 6216
rect 41878 15816 41934 15872
rect 40682 6296 40738 6352
rect 56046 4800 56102 4856
rect 75918 17176 75974 17232
rect 74998 12960 75054 13016
rect 73802 4936 73858 4992
rect 93858 21392 93914 21448
rect 77298 14456 77354 14512
rect 91558 14592 91614 14648
rect 94686 13096 94742 13152
rect 131118 18808 131174 18864
rect 129738 18672 129794 18728
rect 109314 9016 109370 9072
rect 112810 9152 112866 9208
rect 111614 5072 111670 5128
rect 127070 17312 127126 17368
rect 133326 47504 133382 47560
rect 136546 47640 136602 47696
rect 137282 46280 137338 46336
rect 134798 46144 134854 46200
rect 135626 45500 135628 45520
rect 135628 45500 135680 45520
rect 135680 45500 135682 45520
rect 135626 45464 135682 45500
rect 135902 44784 135958 44840
rect 135442 29416 135498 29472
rect 136546 43460 136548 43480
rect 136548 43460 136600 43480
rect 136600 43460 136602 43480
rect 136546 43424 136602 43460
rect 136086 40840 136142 40896
rect 136546 37848 136602 37904
rect 136546 35400 136602 35456
rect 136546 32988 136548 33008
rect 136548 32988 136600 33008
rect 136600 32988 136602 33008
rect 136546 32952 136602 32988
rect 136546 27512 136602 27568
rect 140042 49272 140098 49328
rect 142894 48456 142950 48512
rect 146298 44920 146354 44976
rect 144918 43424 144974 43480
rect 147678 37848 147734 37904
rect 153842 390768 153898 390824
rect 153934 382880 153990 382936
rect 154026 378528 154082 378584
rect 154578 406852 154580 406872
rect 154580 406852 154632 406872
rect 154632 406852 154634 406872
rect 154578 406816 154634 406852
rect 154946 407360 155002 407416
rect 154946 406544 155002 406600
rect 154854 406272 154910 406328
rect 154762 406000 154818 406056
rect 154670 405728 154726 405784
rect 154578 405476 154634 405512
rect 154578 405456 154580 405476
rect 154580 405456 154632 405476
rect 154632 405456 154634 405476
rect 154762 405184 154818 405240
rect 154946 404912 155002 404968
rect 154854 404640 154910 404696
rect 154670 404096 154726 404152
rect 154762 403824 154818 403880
rect 154946 403552 155002 403608
rect 154854 403280 154910 403336
rect 155222 403008 155278 403064
rect 154670 402756 154726 402792
rect 154670 402736 154672 402756
rect 154672 402736 154724 402756
rect 154724 402736 154726 402756
rect 154854 402464 154910 402520
rect 154762 402192 154818 402248
rect 154946 401648 155002 401704
rect 155222 401920 155278 401976
rect 154854 401104 154910 401160
rect 154946 400832 155002 400888
rect 155130 401376 155186 401432
rect 155038 400288 155094 400344
rect 154946 400016 155002 400072
rect 154854 399744 154910 399800
rect 155038 399472 155094 399528
rect 154762 399200 154818 399256
rect 155222 400560 155278 400616
rect 155130 398928 155186 398984
rect 154578 398384 154634 398440
rect 154946 398656 155002 398712
rect 154854 398112 154910 398168
rect 154670 397568 154726 397624
rect 155038 397840 155094 397896
rect 154946 397296 155002 397352
rect 155038 397024 155094 397080
rect 154854 396752 154910 396808
rect 154762 396480 154818 396536
rect 155130 396208 155186 396264
rect 154670 395700 154672 395720
rect 154672 395700 154724 395720
rect 154724 395700 154726 395720
rect 154670 395664 154726 395700
rect 154946 395936 155002 395992
rect 154854 395392 154910 395448
rect 154762 395120 154818 395176
rect 154670 394596 154726 394632
rect 154670 394576 154672 394596
rect 154672 394576 154724 394596
rect 154724 394576 154726 394596
rect 154578 394304 154634 394360
rect 154762 394032 154818 394088
rect 155038 394848 155094 394904
rect 154946 393760 155002 393816
rect 154854 393488 154910 393544
rect 154946 393236 155002 393272
rect 154946 393216 154948 393236
rect 154948 393216 155000 393236
rect 155000 393216 155002 393236
rect 155038 392944 155094 393000
rect 154946 392672 155002 392728
rect 154854 392400 154910 392456
rect 154762 392128 154818 392184
rect 154946 391876 155002 391912
rect 154946 391856 154948 391876
rect 154948 391856 155000 391876
rect 155000 391856 155002 391876
rect 154670 391584 154726 391640
rect 154762 391312 154818 391368
rect 154946 391040 155002 391096
rect 154946 390496 155002 390552
rect 154946 389952 155002 390008
rect 154854 389680 154910 389736
rect 154578 389408 154634 389464
rect 155222 390224 155278 390280
rect 155038 389136 155094 389192
rect 154670 388864 154726 388920
rect 154762 388592 154818 388648
rect 154946 388320 155002 388376
rect 154854 388048 154910 388104
rect 155222 387776 155278 387832
rect 154946 387504 155002 387560
rect 154854 387232 154910 387288
rect 155038 386960 155094 387016
rect 154762 386688 154818 386744
rect 155130 386416 155186 386472
rect 154670 385872 154726 385928
rect 154946 386164 155002 386200
rect 154946 386144 154948 386164
rect 154948 386144 155000 386164
rect 155000 386144 155002 386164
rect 154854 385328 154910 385384
rect 155038 385056 155094 385112
rect 154946 384820 154948 384840
rect 154948 384820 155000 384840
rect 155000 384820 155002 384840
rect 154946 384784 155002 384820
rect 155038 384512 155094 384568
rect 155130 384240 155186 384296
rect 154854 383968 154910 384024
rect 154670 383696 154726 383752
rect 155314 385600 155370 385656
rect 154946 383460 154948 383480
rect 154948 383460 155000 383480
rect 155000 383460 155002 383480
rect 154946 383424 155002 383460
rect 154854 383152 154910 383208
rect 154946 382608 155002 382664
rect 154670 382336 154726 382392
rect 154946 382064 155002 382120
rect 154578 381792 154634 381848
rect 154854 381520 154910 381576
rect 154946 381248 155002 381304
rect 154946 380704 155002 380760
rect 154946 380432 155002 380488
rect 154854 380160 154910 380216
rect 154762 379888 154818 379944
rect 155038 379616 155094 379672
rect 154946 379364 155002 379400
rect 154946 379344 154948 379364
rect 154948 379344 155000 379364
rect 155000 379344 155002 379364
rect 154854 379072 154910 379128
rect 154946 378800 155002 378856
rect 155038 378256 155094 378312
rect 154946 377984 155002 378040
rect 154762 377168 154818 377224
rect 154946 377712 155002 377768
rect 155038 377440 155094 377496
rect 154854 376896 154910 376952
rect 154946 376660 154948 376680
rect 154948 376660 155000 376680
rect 155000 376660 155002 376680
rect 154946 376624 155002 376660
rect 154946 376352 155002 376408
rect 154854 376080 154910 376136
rect 155038 375808 155094 375864
rect 154670 375536 154726 375592
rect 154946 375284 155002 375320
rect 154946 375264 154948 375284
rect 154948 375264 155000 375284
rect 155000 375264 155002 375284
rect 154854 374992 154910 375048
rect 154578 374720 154634 374776
rect 154578 373904 154634 373960
rect 154946 373632 155002 373688
rect 154854 373360 154910 373416
rect 154762 373088 154818 373144
rect 154670 372816 154726 372872
rect 154946 372544 155002 372600
rect 154762 372272 154818 372328
rect 154946 372000 155002 372056
rect 154854 371456 154910 371512
rect 154946 370912 155002 370968
rect 154854 370640 154910 370696
rect 154762 370368 154818 370424
rect 154670 370096 154726 370152
rect 154670 368736 154726 368792
rect 154946 369552 155002 369608
rect 154854 369280 154910 369336
rect 154762 368464 154818 368520
rect 154578 368192 154634 368248
rect 154762 367376 154818 367432
rect 154946 367920 155002 367976
rect 154854 367104 154910 367160
rect 154946 366832 155002 366888
rect 154670 366288 154726 366344
rect 154854 366016 154910 366072
rect 154670 365492 154726 365528
rect 154670 365472 154672 365492
rect 154672 365472 154724 365492
rect 154724 365472 154726 365492
rect 154762 364928 154818 364984
rect 154946 365200 155002 365256
rect 154854 364656 154910 364712
rect 155130 374448 155186 374504
rect 155130 371728 155186 371784
rect 155130 371184 155186 371240
rect 155498 380976 155554 381032
rect 155682 407088 155738 407144
rect 155774 404368 155830 404424
rect 155406 374176 155462 374232
rect 155314 369824 155370 369880
rect 155130 369008 155186 369064
rect 155130 366560 155186 366616
rect 155130 364384 155186 364440
rect 154762 363840 154818 363896
rect 154946 364132 155002 364168
rect 154946 364112 154948 364132
rect 154948 364112 155000 364132
rect 155000 364112 155002 364132
rect 154854 363568 154910 363624
rect 155038 363296 155094 363352
rect 154946 362752 155002 362808
rect 154854 362208 154910 362264
rect 155038 361936 155094 361992
rect 154578 361664 154634 361720
rect 154578 361120 154634 361176
rect 154946 361392 155002 361448
rect 154854 360848 154910 360904
rect 154762 360576 154818 360632
rect 155038 360304 155094 360360
rect 154946 360052 155002 360088
rect 154946 360032 154948 360052
rect 154948 360032 155000 360052
rect 155000 360032 155002 360052
rect 154578 359488 154634 359544
rect 154854 359216 154910 359272
rect 155038 359760 155094 359816
rect 154946 358944 155002 359000
rect 154578 358672 154634 358728
rect 155222 363024 155278 363080
rect 155130 358400 155186 358456
rect 154946 357856 155002 357912
rect 154762 357584 154818 357640
rect 154946 357312 155002 357368
rect 155038 357040 155094 357096
rect 154946 356768 155002 356824
rect 154854 356496 154910 356552
rect 154762 356224 154818 356280
rect 154578 355988 154580 356008
rect 154580 355988 154632 356008
rect 154632 355988 154634 356008
rect 154578 355952 154634 355988
rect 154946 355680 155002 355736
rect 154854 355408 154910 355464
rect 155038 355136 155094 355192
rect 154578 354612 154634 354648
rect 154578 354592 154580 354612
rect 154580 354592 154632 354612
rect 154632 354592 154634 354612
rect 154762 354048 154818 354104
rect 154946 354320 155002 354376
rect 154854 353504 154910 353560
rect 154854 353232 154910 353288
rect 154946 352960 155002 353016
rect 154762 352416 154818 352472
rect 155038 352688 155094 352744
rect 154854 352144 154910 352200
rect 154762 351328 154818 351384
rect 154946 351600 155002 351656
rect 154854 351056 154910 351112
rect 155498 367648 155554 367704
rect 155590 365744 155646 365800
rect 155406 362480 155462 362536
rect 155314 354864 155370 354920
rect 155590 358128 155646 358184
rect 155590 353776 155646 353832
rect 155406 351872 155462 351928
rect 155130 350784 155186 350840
rect 155038 350512 155094 350568
rect 154578 350240 154634 350296
rect 154946 349968 155002 350024
rect 154946 349696 155002 349752
rect 154854 349424 154910 349480
rect 155498 349152 155554 349208
rect 155038 348880 155094 348936
rect 154854 348608 154910 348664
rect 154762 348336 154818 348392
rect 154946 348064 155002 348120
rect 154946 347792 155002 347848
rect 154854 347248 154910 347304
rect 154578 346976 154634 347032
rect 155038 347520 155094 347576
rect 154946 346704 155002 346760
rect 154854 346432 154910 346488
rect 155038 346160 155094 346216
rect 154946 345888 155002 345944
rect 154854 345480 154910 345536
rect 154946 345092 155002 345128
rect 154946 345072 154948 345092
rect 154948 345072 155000 345092
rect 155000 345072 155002 345092
rect 155590 345344 155646 345400
rect 154578 343984 154634 344040
rect 154578 343712 154634 343768
rect 155038 344800 155094 344856
rect 154946 344528 155002 344584
rect 154854 344256 154910 344312
rect 155038 343440 155094 343496
rect 154854 342896 154910 342952
rect 154946 342372 155002 342408
rect 154946 342352 154948 342372
rect 154948 342352 155000 342372
rect 155000 342352 155002 342372
rect 154762 342080 154818 342136
rect 154946 341808 155002 341864
rect 154854 341264 154910 341320
rect 155038 341536 155094 341592
rect 155130 340992 155186 341048
rect 155038 340720 155094 340776
rect 154762 340448 154818 340504
rect 154946 340176 155002 340232
rect 154854 339904 154910 339960
rect 154946 339632 155002 339688
rect 154670 339360 154726 339416
rect 154854 339088 154910 339144
rect 155038 338816 155094 338872
rect 154946 338544 155002 338600
rect 154762 338000 154818 338056
rect 154578 337184 154634 337240
rect 154854 337728 154910 337784
rect 155038 337456 155094 337512
rect 154946 336912 155002 336968
rect 155222 338272 155278 338328
rect 154762 336640 154818 336696
rect 154670 336368 154726 336424
rect 155038 336096 155094 336152
rect 154854 335824 154910 335880
rect 154946 335552 155002 335608
rect 154762 334736 154818 334792
rect 155130 334464 155186 334520
rect 154946 334192 155002 334248
rect 154854 333920 154910 333976
rect 154762 333376 154818 333432
rect 154026 333104 154082 333160
rect 153934 323856 153990 323912
rect 153842 302640 153898 302696
rect 154578 332852 154634 332888
rect 154578 332832 154580 332852
rect 154580 332832 154632 332852
rect 154632 332832 154634 332852
rect 154946 333648 155002 333704
rect 154762 332560 154818 332616
rect 154946 332016 155002 332072
rect 154854 331472 154910 331528
rect 155038 331744 155094 331800
rect 154946 331200 155002 331256
rect 155038 330928 155094 330984
rect 154854 330384 154910 330440
rect 154946 330112 155002 330168
rect 155130 330656 155186 330712
rect 154578 329840 154634 329896
rect 154854 329568 154910 329624
rect 155130 329296 155186 329352
rect 155038 329024 155094 329080
rect 154946 328752 155002 328808
rect 154578 328516 154580 328536
rect 154580 328516 154632 328536
rect 154632 328516 154634 328536
rect 154578 328480 154634 328516
rect 155038 328208 155094 328264
rect 154670 327936 154726 327992
rect 154578 325796 154580 325816
rect 154580 325796 154632 325816
rect 154632 325796 154634 325816
rect 154578 325760 154634 325796
rect 154578 321680 154634 321736
rect 154854 327664 154910 327720
rect 154946 327392 155002 327448
rect 154762 327120 154818 327176
rect 154854 326848 154910 326904
rect 154762 326304 154818 326360
rect 154946 326576 155002 326632
rect 155038 326032 155094 326088
rect 155038 325488 155094 325544
rect 154762 325216 154818 325272
rect 154854 324944 154910 325000
rect 154946 324672 155002 324728
rect 154946 324400 155002 324456
rect 155038 324128 155094 324184
rect 154946 323584 155002 323640
rect 154854 323312 154910 323368
rect 154946 323076 154948 323096
rect 154948 323076 155000 323096
rect 155000 323076 155002 323096
rect 154946 323040 155002 323076
rect 155038 322768 155094 322824
rect 154762 322496 154818 322552
rect 154854 322224 154910 322280
rect 154946 321952 155002 322008
rect 155038 321408 155094 321464
rect 154762 321136 154818 321192
rect 154946 320864 155002 320920
rect 154854 320592 154910 320648
rect 154946 320320 155002 320376
rect 154854 320048 154910 320104
rect 154762 319776 154818 319832
rect 155038 319504 155094 319560
rect 154946 319232 155002 319288
rect 154670 318688 154726 318744
rect 154762 318416 154818 318472
rect 155038 318144 155094 318200
rect 154854 317872 154910 317928
rect 154946 317636 154948 317656
rect 154948 317636 155000 317656
rect 155000 317636 155002 317656
rect 154946 317600 155002 317636
rect 154762 317328 154818 317384
rect 154578 316784 154634 316840
rect 154854 317056 154910 317112
rect 155038 316512 155094 316568
rect 154946 316240 155002 316296
rect 155038 315968 155094 316024
rect 154854 315696 154910 315752
rect 154762 315424 154818 315480
rect 154946 315152 155002 315208
rect 154762 314608 154818 314664
rect 154578 313792 154634 313848
rect 154854 314336 154910 314392
rect 154946 313556 154948 313576
rect 154948 313556 155000 313576
rect 155000 313556 155002 313576
rect 154946 313520 155002 313556
rect 154946 313248 155002 313304
rect 154854 312976 154910 313032
rect 154762 312704 154818 312760
rect 154578 312432 154634 312488
rect 154946 312180 155002 312216
rect 154946 312160 154948 312180
rect 154948 312160 155000 312180
rect 155000 312160 155002 312180
rect 154578 311908 154634 311944
rect 154578 311888 154580 311908
rect 154580 311888 154632 311908
rect 154632 311888 154634 311908
rect 154762 311616 154818 311672
rect 154578 309712 154634 309768
rect 154578 308080 154634 308136
rect 154578 304000 154634 304056
rect 154854 311344 154910 311400
rect 155038 311072 155094 311128
rect 154946 310800 155002 310856
rect 154854 310528 154910 310584
rect 154854 310256 154910 310312
rect 154762 309984 154818 310040
rect 154946 309440 155002 309496
rect 154946 309188 155002 309224
rect 154946 309168 154948 309188
rect 154948 309168 155000 309188
rect 155000 309168 155002 309188
rect 155038 308896 155094 308952
rect 154762 308624 154818 308680
rect 154854 308352 154910 308408
rect 154946 307808 155002 307864
rect 155038 307536 155094 307592
rect 154762 307264 154818 307320
rect 154946 306992 155002 307048
rect 154854 306720 154910 306776
rect 154946 306468 155002 306504
rect 154946 306448 154948 306468
rect 154948 306448 155000 306468
rect 155000 306448 155002 306468
rect 154854 306176 154910 306232
rect 154762 305904 154818 305960
rect 154946 305360 155002 305416
rect 154854 304816 154910 304872
rect 154762 303728 154818 303784
rect 154946 304544 155002 304600
rect 154946 303456 155002 303512
rect 154854 302912 154910 302968
rect 154670 302404 154672 302424
rect 154672 302404 154724 302424
rect 154724 302404 154726 302424
rect 154670 302368 154726 302404
rect 155130 305088 155186 305144
rect 155130 303184 155186 303240
rect 154854 302096 154910 302152
rect 154762 301824 154818 301880
rect 154670 301552 154726 301608
rect 154578 301280 154634 301336
rect 154854 300464 154910 300520
rect 154762 300192 154818 300248
rect 154670 299920 154726 299976
rect 154578 299668 154634 299704
rect 154578 299648 154580 299668
rect 154580 299648 154632 299668
rect 154632 299648 154634 299668
rect 154762 299376 154818 299432
rect 154578 298832 154634 298888
rect 154670 298288 154726 298344
rect 154578 297472 154634 297528
rect 154946 299104 155002 299160
rect 154854 298560 154910 298616
rect 154946 298016 155002 298072
rect 154762 297744 154818 297800
rect 155038 297200 155094 297256
rect 154854 296656 154910 296712
rect 154762 296112 154818 296168
rect 154670 295840 154726 295896
rect 154578 295604 154580 295624
rect 154580 295604 154632 295624
rect 154632 295604 154634 295624
rect 154578 295568 154634 295604
rect 154946 296384 155002 296440
rect 154762 295024 154818 295080
rect 154670 294752 154726 294808
rect 154578 294208 154634 294264
rect 154854 294480 154910 294536
rect 154578 293972 154580 293992
rect 154580 293972 154632 293992
rect 154632 293972 154634 293992
rect 154578 293936 154634 293972
rect 154578 293664 154634 293720
rect 154670 293392 154726 293448
rect 154578 292596 154634 292632
rect 154578 292576 154580 292596
rect 154580 292576 154632 292596
rect 154632 292576 154634 292596
rect 155498 343168 155554 343224
rect 155682 342624 155738 342680
rect 155590 335280 155646 335336
rect 155866 335008 155922 335064
rect 155774 332288 155830 332344
rect 155498 318960 155554 319016
rect 155590 314880 155646 314936
rect 155682 314064 155738 314120
rect 155590 305632 155646 305688
rect 155314 300736 155370 300792
rect 155222 292848 155278 292904
rect 155498 304272 155554 304328
rect 155590 301008 155646 301064
rect 155498 296928 155554 296984
rect 155406 295296 155462 295352
rect 155314 292304 155370 292360
rect 152554 49136 152610 49192
rect 154946 129920 155002 129976
rect 154946 128016 155002 128072
rect 154946 126112 155002 126168
rect 154486 124208 154542 124264
rect 154946 122304 155002 122360
rect 154578 120400 154634 120456
rect 154578 118496 154634 118552
rect 154762 114688 154818 114744
rect 154946 112784 155002 112840
rect 154854 110880 154910 110936
rect 154578 105168 154634 105224
rect 154578 103264 154634 103320
rect 154946 101360 155002 101416
rect 154946 99456 155002 99512
rect 154854 97552 154910 97608
rect 154946 95648 155002 95704
rect 154578 93744 154634 93800
rect 154946 91840 155002 91896
rect 154946 89936 155002 89992
rect 154946 88032 155002 88088
rect 154946 86128 155002 86184
rect 154946 84244 155002 84280
rect 154946 84224 154948 84244
rect 154948 84224 155000 84244
rect 155000 84224 155002 84244
rect 154946 82320 155002 82376
rect 154762 80416 154818 80472
rect 154946 78512 155002 78568
rect 154946 76608 155002 76664
rect 154946 74704 155002 74760
rect 154578 72800 154634 72856
rect 154946 70896 155002 70952
rect 154578 69028 154580 69048
rect 154580 69028 154632 69048
rect 154632 69028 154634 69048
rect 154578 68992 154634 69028
rect 154946 67088 155002 67144
rect 154578 65184 154634 65240
rect 154578 63280 154634 63336
rect 154946 61376 155002 61432
rect 154946 59472 155002 59528
rect 154946 57568 155002 57624
rect 154946 55664 155002 55720
rect 154946 53760 155002 53816
rect 153934 48864 153990 48920
rect 155406 116592 155462 116648
rect 155498 108976 155554 109032
rect 155314 107072 155370 107128
rect 157982 52128 158038 52184
rect 158074 50088 158130 50144
rect 157890 49544 157946 49600
rect 149058 35128 149114 35184
rect 216678 52828 216734 52864
rect 216678 52808 216680 52828
rect 216680 52808 216732 52828
rect 216732 52808 216734 52828
rect 159914 51584 159970 51640
rect 159362 51040 159418 51096
rect 158258 49000 158314 49056
rect 160328 51856 160384 51912
rect 160190 51720 160246 51776
rect 160512 51822 160568 51878
rect 160972 51856 161028 51912
rect 160650 51584 160706 51640
rect 161156 51720 161212 51776
rect 161340 51890 161396 51946
rect 161386 51720 161442 51776
rect 161708 51856 161764 51912
rect 161984 51856 162040 51912
rect 160742 46008 160798 46064
rect 160742 24112 160798 24168
rect 161754 51584 161810 51640
rect 161386 48864 161442 48920
rect 161754 48864 161810 48920
rect 162444 51856 162500 51912
rect 162030 45872 162086 45928
rect 162306 51448 162362 51504
rect 162720 51856 162776 51912
rect 162996 51808 163052 51810
rect 162996 51756 162998 51808
rect 162998 51756 163050 51808
rect 163050 51756 163052 51808
rect 162996 51754 163052 51756
rect 162766 51448 162822 51504
rect 162858 51060 162914 51096
rect 162858 51040 162860 51060
rect 162860 51040 162912 51060
rect 162912 51040 162914 51060
rect 162950 48864 163006 48920
rect 163456 51856 163512 51912
rect 163640 51754 163696 51810
rect 163916 51856 163972 51912
rect 164100 51856 164156 51912
rect 164468 51856 164524 51912
rect 164054 51720 164110 51776
rect 164744 51856 164800 51912
rect 163134 48728 163190 48784
rect 163318 48728 163374 48784
rect 163502 51584 163558 51640
rect 163410 46824 163466 46880
rect 164422 48592 164478 48648
rect 164882 51720 164938 51776
rect 164698 51312 164754 51368
rect 165388 51890 165444 51946
rect 165572 51890 165628 51946
rect 165848 51890 165904 51946
rect 166124 51856 166180 51912
rect 166676 51890 166732 51946
rect 165296 51720 165352 51776
rect 165066 51584 165122 51640
rect 165250 51448 165306 51504
rect 165158 51312 165214 51368
rect 165434 51584 165490 51640
rect 166768 51720 166824 51776
rect 165802 51312 165858 51368
rect 165710 49408 165766 49464
rect 165894 49408 165950 49464
rect 167596 51890 167652 51946
rect 166952 51822 167008 51878
rect 167274 51720 167330 51776
rect 167412 51756 167414 51776
rect 167414 51756 167466 51776
rect 167466 51756 167468 51776
rect 167780 51890 167836 51946
rect 167964 51822 168020 51878
rect 167412 51720 167468 51756
rect 166722 51584 166778 51640
rect 166630 51448 166686 51504
rect 163686 6160 163742 6216
rect 166722 47368 166778 47424
rect 167090 47368 167146 47424
rect 167274 47640 167330 47696
rect 167182 46144 167238 46200
rect 167366 47504 167422 47560
rect 168608 51890 168664 51946
rect 168792 51856 168848 51912
rect 167734 51584 167790 51640
rect 167734 51448 167790 51504
rect 168976 51720 169032 51776
rect 168654 51584 168710 51640
rect 168562 48048 168618 48104
rect 167826 45736 167882 45792
rect 167182 4800 167238 4856
rect 168746 51448 168802 51504
rect 169712 51890 169768 51946
rect 169758 51448 169814 51504
rect 170172 51856 170228 51912
rect 170080 51720 170136 51776
rect 170632 51856 170688 51912
rect 170126 51620 170128 51640
rect 170128 51620 170180 51640
rect 170180 51620 170182 51640
rect 170126 51584 170182 51620
rect 169666 50224 169722 50280
rect 169942 51312 169998 51368
rect 170126 51040 170182 51096
rect 170770 51720 170826 51776
rect 170310 48728 170366 48784
rect 170310 48592 170366 48648
rect 170586 51584 170642 51640
rect 170862 51448 170918 51504
rect 170770 50224 170826 50280
rect 171276 51856 171332 51912
rect 171046 50768 171102 50824
rect 171644 51856 171700 51912
rect 171230 51448 171286 51504
rect 171414 51312 171470 51368
rect 171598 51584 171654 51640
rect 171506 51176 171562 51232
rect 172104 51822 172160 51878
rect 172656 51822 172712 51878
rect 172334 51448 172390 51504
rect 172334 51312 172390 51368
rect 172518 51448 172574 51504
rect 172426 49408 172482 49464
rect 172150 48864 172206 48920
rect 173116 51856 173172 51912
rect 172794 51448 172850 51504
rect 172886 50496 172942 50552
rect 173070 51312 173126 51368
rect 173760 51856 173816 51912
rect 173944 51856 174000 51912
rect 173162 47504 173218 47560
rect 173852 51720 173908 51776
rect 174220 51720 174276 51776
rect 174404 51856 174460 51912
rect 174450 51720 174506 51776
rect 174634 51720 174690 51776
rect 174864 51856 174920 51912
rect 173806 51448 173862 51504
rect 174174 51312 174230 51368
rect 174358 50768 174414 50824
rect 173990 49952 174046 50008
rect 174266 49952 174322 50008
rect 173990 48184 174046 48240
rect 175278 51040 175334 51096
rect 174266 48048 174322 48104
rect 175646 51720 175702 51776
rect 176152 51890 176208 51946
rect 176106 51720 176162 51776
rect 176474 50088 176530 50144
rect 177026 49564 177082 49600
rect 177026 49544 177028 49564
rect 177028 49544 177080 49564
rect 177080 49544 177082 49564
rect 177118 49000 177174 49056
rect 176934 48592 176990 48648
rect 174542 46144 174598 46200
rect 177532 51890 177588 51946
rect 177302 49272 177358 49328
rect 177992 51856 178048 51912
rect 177762 51448 177818 51504
rect 177762 50088 177818 50144
rect 178636 51856 178692 51912
rect 178912 51856 178968 51912
rect 177762 49952 177818 50008
rect 177670 49136 177726 49192
rect 177578 48456 177634 48512
rect 177854 49272 177910 49328
rect 177946 49136 178002 49192
rect 177946 48900 177948 48920
rect 177948 48900 178000 48920
rect 178000 48900 178002 48920
rect 177946 48864 178002 48900
rect 178314 48320 178370 48376
rect 178958 51720 179014 51776
rect 179648 51856 179704 51912
rect 178866 51448 178922 51504
rect 178774 51040 178830 51096
rect 177670 24792 177726 24848
rect 179142 51196 179198 51232
rect 179142 51176 179144 51196
rect 179144 51176 179196 51196
rect 179196 51176 179198 51196
rect 180384 51856 180440 51912
rect 179970 47912 180026 47968
rect 180154 47912 180210 47968
rect 181028 51890 181084 51946
rect 181304 51890 181360 51946
rect 180430 47912 180486 47968
rect 180890 48456 180946 48512
rect 181258 48320 181314 48376
rect 181166 47912 181222 47968
rect 181074 44784 181130 44840
rect 182408 51890 182464 51946
rect 182960 51890 183016 51946
rect 182454 49680 182510 49736
rect 182362 49000 182418 49056
rect 182270 48728 182326 48784
rect 182178 47504 182234 47560
rect 182546 48456 182602 48512
rect 183604 51856 183660 51912
rect 184156 51856 184212 51912
rect 183926 49680 183982 49736
rect 184616 51856 184672 51912
rect 183650 46144 183706 46200
rect 185628 51856 185684 51912
rect 184478 48728 184534 48784
rect 184570 48456 184626 48512
rect 184754 48320 184810 48376
rect 186042 48456 186098 48512
rect 186134 48320 186190 48376
rect 187008 51856 187064 51912
rect 186502 50088 186558 50144
rect 187146 49000 187202 49056
rect 187238 48456 187294 48512
rect 187146 48320 187202 48376
rect 187606 48728 187662 48784
rect 187514 48592 187570 48648
rect 187422 48320 187478 48376
rect 188848 51856 188904 51912
rect 188894 48592 188950 48648
rect 188986 48320 189042 48376
rect 189262 49952 189318 50008
rect 189722 48320 189778 48376
rect 189814 45464 189870 45520
rect 190090 44376 190146 44432
rect 190550 3984 190606 4040
rect 191378 49952 191434 50008
rect 191470 49816 191526 49872
rect 190734 3848 190790 3904
rect 191746 50088 191802 50144
rect 191654 49952 191710 50008
rect 192528 51890 192584 51946
rect 192896 51856 192952 51912
rect 193356 51856 193412 51912
rect 193540 51890 193596 51946
rect 192942 48728 192998 48784
rect 193126 48592 193182 48648
rect 193034 48456 193090 48512
rect 193908 51856 193964 51912
rect 193586 47368 193642 47424
rect 193862 49952 193918 50008
rect 194828 51856 194884 51912
rect 195104 51856 195160 51912
rect 195472 51890 195528 51946
rect 195840 51890 195896 51946
rect 194230 50088 194286 50144
rect 194414 47504 194470 47560
rect 194322 47368 194378 47424
rect 194690 47504 194746 47560
rect 194874 47368 194930 47424
rect 195702 49680 195758 49736
rect 195610 47504 195666 47560
rect 196576 51856 196632 51912
rect 195886 47640 195942 47696
rect 195794 47368 195850 47424
rect 195610 47232 195666 47288
rect 196346 49680 196402 49736
rect 196070 21392 196126 21448
rect 197128 51856 197184 51912
rect 197266 48592 197322 48648
rect 198416 51856 198472 51912
rect 198600 51890 198656 51946
rect 198462 48864 198518 48920
rect 198554 48592 198610 48648
rect 199014 48320 199070 48376
rect 199842 48592 199898 48648
rect 199934 48456 199990 48512
rect 199750 48320 199806 48376
rect 200026 41384 200082 41440
rect 200026 35944 200082 36000
rect 201268 51856 201324 51912
rect 201820 51890 201876 51946
rect 201406 48320 201462 48376
rect 201498 46144 201554 46200
rect 202372 51856 202428 51912
rect 202050 49680 202106 49736
rect 201958 46688 202014 46744
rect 201866 46416 201922 46472
rect 201866 46144 201922 46200
rect 202510 48864 202566 48920
rect 202602 48592 202658 48648
rect 202786 48456 202842 48512
rect 202694 48320 202750 48376
rect 204120 51856 204176 51912
rect 204488 51856 204544 51912
rect 204166 50088 204222 50144
rect 203982 48864 204038 48920
rect 203798 48320 203854 48376
rect 205224 51890 205280 51946
rect 205408 51856 205464 51912
rect 204534 50088 204590 50144
rect 204902 49816 204958 49872
rect 205454 50088 205510 50144
rect 205362 48320 205418 48376
rect 206144 51890 206200 51946
rect 206328 51890 206384 51946
rect 206880 51890 206936 51946
rect 207064 51856 207120 51912
rect 206190 49952 206246 50008
rect 206466 48320 206522 48376
rect 207340 51720 207396 51776
rect 207616 51720 207672 51776
rect 206926 50088 206982 50144
rect 206834 49952 206890 50008
rect 207386 50088 207442 50144
rect 208168 51856 208224 51912
rect 207018 4800 207074 4856
rect 208076 51720 208132 51776
rect 208030 49816 208086 49872
rect 208306 50088 208362 50144
rect 208306 48592 208362 48648
rect 208996 51856 209052 51912
rect 208950 51720 209006 51776
rect 209272 51856 209328 51912
rect 209640 51890 209696 51946
rect 209548 51720 209604 51776
rect 209134 48900 209136 48920
rect 209136 48900 209188 48920
rect 209188 48900 209190 48920
rect 209134 48864 209190 48900
rect 210284 51856 210340 51912
rect 209318 50088 209374 50144
rect 209594 50088 209650 50144
rect 209594 49680 209650 49736
rect 209778 49952 209834 50008
rect 209870 49680 209926 49736
rect 209778 49000 209834 49056
rect 209778 48728 209834 48784
rect 210054 48864 210110 48920
rect 210560 51856 210616 51912
rect 210928 51856 210984 51912
rect 210330 48728 210386 48784
rect 211112 51890 211168 51946
rect 210790 48728 210846 48784
rect 211066 50088 211122 50144
rect 211664 51720 211720 51776
rect 211342 50088 211398 50144
rect 210422 17176 210478 17232
rect 211250 45736 211306 45792
rect 212308 51890 212364 51946
rect 212492 51856 212548 51912
rect 212216 51720 212272 51776
rect 212262 48728 212318 48784
rect 211802 17720 211858 17776
rect 213320 51856 213376 51912
rect 213366 51720 213422 51776
rect 213872 51856 213928 51912
rect 213688 51756 213690 51776
rect 213690 51756 213742 51776
rect 213742 51756 213744 51776
rect 213688 51720 213744 51756
rect 213826 51720 213882 51776
rect 213642 49952 213698 50008
rect 213826 48864 213882 48920
rect 214194 49680 214250 49736
rect 214792 51890 214848 51946
rect 214700 51720 214756 51776
rect 214194 48320 214250 48376
rect 214562 47912 214618 47968
rect 215022 48864 215078 48920
rect 214838 48320 214894 48376
rect 215528 51890 215584 51946
rect 215206 48728 215262 48784
rect 215114 47912 215170 47968
rect 215758 48728 215814 48784
rect 216402 49816 216458 49872
rect 217322 47504 217378 47560
rect 219714 413072 219770 413128
rect 219990 413480 220046 413536
rect 219806 412664 219862 412720
rect 219898 411440 219954 411496
rect 219806 410624 219862 410680
rect 220082 411884 220084 411904
rect 220084 411884 220136 411904
rect 220136 411884 220138 411904
rect 220082 411848 220138 411884
rect 220082 410216 220138 410272
rect 219990 409400 220046 409456
rect 220082 408992 220138 409048
rect 219898 408584 219954 408640
rect 219898 407768 219954 407824
rect 220082 407360 220138 407416
rect 219898 406136 219954 406192
rect 220082 405728 220138 405784
rect 219898 404912 219954 404968
rect 220082 404504 220138 404560
rect 220082 403688 220138 403744
rect 219990 403280 220046 403336
rect 219806 402872 219862 402928
rect 219714 402464 219770 402520
rect 220174 401648 220230 401704
rect 220082 401276 220084 401296
rect 220084 401276 220136 401296
rect 220136 401276 220138 401296
rect 220082 401240 220138 401276
rect 220174 400424 220230 400480
rect 219990 400016 220046 400072
rect 220082 399200 220138 399256
rect 220174 398792 220230 398848
rect 220082 397976 220138 398032
rect 220174 397568 220230 397624
rect 220174 396344 220230 396400
rect 219898 395936 219954 395992
rect 220082 395528 220138 395584
rect 220174 395120 220230 395176
rect 219990 393896 220046 393952
rect 220174 393488 220230 393544
rect 220266 392672 220322 392728
rect 220174 392264 220230 392320
rect 219898 389816 219954 389872
rect 220082 388184 220138 388240
rect 220266 391040 220322 391096
rect 220450 390632 220506 390688
rect 220358 389408 220414 389464
rect 220450 388592 220506 388648
rect 220174 387776 220230 387832
rect 220266 386960 220322 387016
rect 220450 386552 220506 386608
rect 220174 385736 220230 385792
rect 220450 385328 220506 385384
rect 220358 384920 220414 384976
rect 220266 384104 220322 384160
rect 220082 383288 220138 383344
rect 219714 380024 219770 380080
rect 219438 374720 219494 374776
rect 219990 375944 220046 376000
rect 219990 375536 220046 375592
rect 219898 373496 219954 373552
rect 218702 52128 218758 52184
rect 219990 371456 220046 371512
rect 219714 368600 219770 368656
rect 219898 367376 219954 367432
rect 219622 365744 219678 365800
rect 219990 365336 220046 365392
rect 219714 364520 219770 364576
rect 219898 360440 219954 360496
rect 219714 358808 219770 358864
rect 219438 358400 219494 358456
rect 219990 357584 220046 357640
rect 219898 356768 219954 356824
rect 219806 354728 219862 354784
rect 219898 351872 219954 351928
rect 219990 351056 220046 351112
rect 219898 350648 219954 350704
rect 219898 349424 219954 349480
rect 219898 343712 219954 343768
rect 219806 341672 219862 341728
rect 219898 340484 219900 340504
rect 219900 340484 219952 340504
rect 219952 340484 219954 340504
rect 219898 340448 219954 340484
rect 219530 339632 219586 339688
rect 219898 338000 219954 338056
rect 219990 334736 220046 334792
rect 219806 333124 219862 333160
rect 219806 333104 219808 333124
rect 219808 333104 219860 333124
rect 219860 333104 219862 333124
rect 219898 332288 219954 332344
rect 219898 331492 219954 331528
rect 219898 331472 219900 331492
rect 219900 331472 219952 331492
rect 219952 331472 219954 331492
rect 219714 330656 219770 330712
rect 219530 329044 219586 329080
rect 219530 329024 219532 329044
rect 219532 329024 219584 329044
rect 219584 329024 219586 329044
rect 219530 326984 219586 327040
rect 219898 324944 219954 325000
rect 219714 323332 219770 323368
rect 219714 323312 219716 323332
rect 219716 323312 219768 323332
rect 219768 323312 219770 323332
rect 218794 48456 218850 48512
rect 219990 318436 220046 318472
rect 219990 318416 219992 318436
rect 219992 318416 220044 318436
rect 220044 318416 220046 318436
rect 219990 315560 220046 315616
rect 219898 313112 219954 313168
rect 219714 309032 219770 309088
rect 219898 308624 219954 308680
rect 219898 302912 219954 302968
rect 219990 301280 220046 301336
rect 219990 298832 220046 298888
rect 219898 295976 219954 296032
rect 219898 294752 219954 294808
rect 219898 292304 219954 292360
rect 219530 288224 219586 288280
rect 219898 287000 219954 287056
rect 219898 286592 219954 286648
rect 220450 383696 220506 383752
rect 220450 382880 220506 382936
rect 220542 382472 220598 382528
rect 220726 413888 220782 413944
rect 220726 412256 220782 412312
rect 220726 411032 220782 411088
rect 220726 409808 220782 409864
rect 220726 408176 220782 408232
rect 220726 406988 220728 407008
rect 220728 406988 220780 407008
rect 220780 406988 220782 407008
rect 220726 406952 220782 406988
rect 220726 406544 220782 406600
rect 220726 405356 220728 405376
rect 220728 405356 220780 405376
rect 220780 405356 220782 405376
rect 220726 405320 220782 405356
rect 220726 404096 220782 404152
rect 220726 402056 220782 402112
rect 220726 400832 220782 400888
rect 220726 399608 220782 399664
rect 220726 398384 220782 398440
rect 220726 397160 220782 397216
rect 220726 396752 220782 396808
rect 220726 394712 220782 394768
rect 220726 394304 220782 394360
rect 220726 393080 220782 393136
rect 220726 391876 220782 391912
rect 220726 391856 220728 391876
rect 220728 391856 220780 391876
rect 220780 391856 220782 391876
rect 220726 391484 220728 391504
rect 220728 391484 220780 391504
rect 220780 391484 220782 391504
rect 220726 391448 220782 391484
rect 220726 390224 220782 390280
rect 220726 389000 220782 389056
rect 220726 387368 220782 387424
rect 220726 386144 220782 386200
rect 220726 384512 220782 384568
rect 220726 382064 220782 382120
rect 220634 381656 220690 381712
rect 220542 381248 220598 381304
rect 220726 380840 220782 380896
rect 220726 380468 220728 380488
rect 220728 380468 220780 380488
rect 220780 380468 220782 380488
rect 220726 380432 220782 380468
rect 220634 379616 220690 379672
rect 220542 378800 220598 378856
rect 220726 379208 220782 379264
rect 220634 378392 220690 378448
rect 220726 378020 220728 378040
rect 220728 378020 220780 378040
rect 220780 378020 220782 378040
rect 220726 377984 220782 378020
rect 220634 377576 220690 377632
rect 220542 377168 220598 377224
rect 220450 376760 220506 376816
rect 220726 376352 220782 376408
rect 220726 375128 220782 375184
rect 220634 374312 220690 374368
rect 220542 373904 220598 373960
rect 220634 373088 220690 373144
rect 220726 372680 220782 372736
rect 220358 372308 220360 372328
rect 220360 372308 220412 372328
rect 220412 372308 220414 372328
rect 220358 372272 220414 372308
rect 220450 371864 220506 371920
rect 220634 371068 220690 371104
rect 220634 371048 220636 371068
rect 220636 371048 220688 371068
rect 220688 371048 220690 371068
rect 220726 370640 220782 370696
rect 220542 370232 220598 370288
rect 220542 369824 220598 369880
rect 220634 369416 220690 369472
rect 220634 369008 220690 369064
rect 220726 368192 220782 368248
rect 220542 367784 220598 367840
rect 220726 366988 220782 367024
rect 220726 366968 220728 366988
rect 220728 366968 220780 366988
rect 220780 366968 220782 366988
rect 220542 366560 220598 366616
rect 220634 366152 220690 366208
rect 220634 364928 220690 364984
rect 220542 364148 220544 364168
rect 220544 364148 220596 364168
rect 220596 364148 220598 364168
rect 220542 364112 220598 364148
rect 220726 363704 220782 363760
rect 220634 363296 220690 363352
rect 220726 362888 220782 362944
rect 220450 362108 220452 362128
rect 220452 362108 220504 362128
rect 220504 362108 220506 362128
rect 220450 362072 220506 362108
rect 220634 362480 220690 362536
rect 220542 361664 220598 361720
rect 220450 360884 220452 360904
rect 220452 360884 220504 360904
rect 220504 360884 220506 360904
rect 220450 360848 220506 360884
rect 220726 361256 220782 361312
rect 220634 360032 220690 360088
rect 220726 359624 220782 359680
rect 220726 359252 220728 359272
rect 220728 359252 220780 359272
rect 220780 359252 220782 359272
rect 220726 359216 220782 359252
rect 220634 357992 220690 358048
rect 220634 357212 220636 357232
rect 220636 357212 220688 357232
rect 220688 357212 220690 357232
rect 220634 357176 220690 357212
rect 220726 356360 220782 356416
rect 220726 355988 220728 356008
rect 220728 355988 220780 356008
rect 220780 355988 220782 356008
rect 220726 355952 220782 355988
rect 220726 355544 220782 355600
rect 220542 355136 220598 355192
rect 220634 354356 220636 354376
rect 220636 354356 220688 354376
rect 220688 354356 220690 354376
rect 220634 354320 220690 354356
rect 220542 353504 220598 353560
rect 220450 352724 220452 352744
rect 220452 352724 220504 352744
rect 220504 352724 220506 352744
rect 220450 352688 220506 352724
rect 220450 352280 220506 352336
rect 220358 350240 220414 350296
rect 220542 349832 220598 349888
rect 220726 353912 220782 353968
rect 220726 353096 220782 353152
rect 220726 351464 220782 351520
rect 220542 349036 220598 349072
rect 220542 349016 220544 349036
rect 220544 349016 220596 349036
rect 220596 349016 220598 349036
rect 220450 347792 220506 347848
rect 220450 346976 220506 347032
rect 220358 344936 220414 344992
rect 220450 342524 220452 342544
rect 220452 342524 220504 342544
rect 220504 342524 220506 342544
rect 220450 342488 220506 342524
rect 220726 348608 220782 348664
rect 220634 348200 220690 348256
rect 220726 347384 220782 347440
rect 220634 346568 220690 346624
rect 220726 346160 220782 346216
rect 220726 345752 220782 345808
rect 220634 345344 220690 345400
rect 220726 344528 220782 344584
rect 220634 344120 220690 344176
rect 220634 343340 220636 343360
rect 220636 343340 220688 343360
rect 220688 343340 220690 343360
rect 220634 343304 220690 343340
rect 220726 342896 220782 342952
rect 220726 342116 220728 342136
rect 220728 342116 220780 342136
rect 220780 342116 220782 342136
rect 220726 342080 220782 342116
rect 220542 341264 220598 341320
rect 220266 340856 220322 340912
rect 220174 340040 220230 340096
rect 220726 339224 220782 339280
rect 220634 338816 220690 338872
rect 220450 338408 220506 338464
rect 220634 337592 220690 337648
rect 220542 336776 220598 336832
rect 220726 337184 220782 337240
rect 220634 336368 220690 336424
rect 220542 335960 220598 336016
rect 220726 335572 220782 335608
rect 220726 335552 220728 335572
rect 220728 335552 220780 335572
rect 220780 335552 220782 335572
rect 220174 335144 220230 335200
rect 220358 334328 220414 334384
rect 220450 333920 220506 333976
rect 220634 333512 220690 333568
rect 220726 332696 220782 332752
rect 220542 331880 220598 331936
rect 220542 331064 220598 331120
rect 220726 330248 220782 330304
rect 220634 329840 220690 329896
rect 220542 329432 220598 329488
rect 220726 328616 220782 328672
rect 220266 328208 220322 328264
rect 220266 327800 220322 327856
rect 220726 327392 220782 327448
rect 220634 326576 220690 326632
rect 220358 326168 220414 326224
rect 220726 325780 220782 325816
rect 220726 325760 220728 325780
rect 220728 325760 220780 325780
rect 220780 325760 220782 325780
rect 220266 325352 220322 325408
rect 220726 324572 220728 324592
rect 220728 324572 220780 324592
rect 220780 324572 220782 324592
rect 220726 324536 220782 324572
rect 220266 324128 220322 324184
rect 220266 321272 220322 321328
rect 220266 320456 220322 320512
rect 220634 323720 220690 323776
rect 220726 322904 220782 322960
rect 220542 322496 220598 322552
rect 220634 322088 220690 322144
rect 220726 321700 220782 321736
rect 220726 321680 220728 321700
rect 220728 321680 220780 321700
rect 220780 321680 220782 321700
rect 220726 320864 220782 320920
rect 220450 320048 220506 320104
rect 220450 319640 220506 319696
rect 220358 319232 220414 319288
rect 220726 318824 220782 318880
rect 220634 318008 220690 318064
rect 220726 317600 220782 317656
rect 220726 317192 220782 317248
rect 220634 316784 220690 316840
rect 220450 316376 220506 316432
rect 220634 315968 220690 316024
rect 220542 314780 220544 314800
rect 220544 314780 220596 314800
rect 220596 314780 220598 314800
rect 220542 314744 220598 314780
rect 220726 315152 220782 315208
rect 220634 314336 220690 314392
rect 220450 313928 220506 313984
rect 220726 313520 220782 313576
rect 220450 312704 220506 312760
rect 220450 312296 220506 312352
rect 220726 311924 220728 311944
rect 220728 311924 220780 311944
rect 220780 311924 220782 311944
rect 220726 311888 220782 311924
rect 220634 311480 220690 311536
rect 220542 310684 220598 310720
rect 220542 310664 220544 310684
rect 220544 310664 220596 310684
rect 220596 310664 220598 310684
rect 220726 311072 220782 311128
rect 220726 310256 220782 310312
rect 220542 309848 220598 309904
rect 220634 309460 220690 309496
rect 220634 309440 220636 309460
rect 220636 309440 220688 309460
rect 220688 309440 220690 309460
rect 220634 308216 220690 308272
rect 220726 307808 220782 307864
rect 220542 307400 220598 307456
rect 220634 306992 220690 307048
rect 220726 306584 220782 306640
rect 220542 306176 220598 306232
rect 220634 305768 220690 305824
rect 220726 305380 220782 305416
rect 220726 305360 220728 305380
rect 220728 305360 220780 305380
rect 220780 305360 220782 305380
rect 220726 304952 220782 305008
rect 220450 304544 220506 304600
rect 220634 304136 220690 304192
rect 220726 303748 220782 303784
rect 220726 303728 220728 303748
rect 220728 303728 220780 303748
rect 220780 303728 220782 303748
rect 220542 303320 220598 303376
rect 220726 302504 220782 302560
rect 220634 302096 220690 302152
rect 220542 301688 220598 301744
rect 220726 300872 220782 300928
rect 220634 300056 220690 300112
rect 220726 299648 220782 299704
rect 220542 299240 220598 299296
rect 220726 298424 220782 298480
rect 220634 298016 220690 298072
rect 220358 296792 220414 296848
rect 220266 295160 220322 295216
rect 220266 290264 220322 290320
rect 220726 297628 220782 297664
rect 220726 297608 220728 297628
rect 220728 297608 220780 297628
rect 220780 297608 220782 297628
rect 220726 297200 220782 297256
rect 220634 296384 220690 296440
rect 220726 295568 220782 295624
rect 220726 294344 220782 294400
rect 220450 293936 220506 293992
rect 220634 293528 220690 293584
rect 220542 292732 220598 292768
rect 220542 292712 220544 292732
rect 220544 292712 220596 292732
rect 220596 292712 220598 292732
rect 220726 293120 220782 293176
rect 220634 291896 220690 291952
rect 220726 291488 220782 291544
rect 220726 291080 220782 291136
rect 220634 290672 220690 290728
rect 220726 289876 220782 289912
rect 220726 289856 220728 289876
rect 220728 289856 220780 289876
rect 220780 289856 220782 289876
rect 220542 289448 220598 289504
rect 220634 289040 220690 289096
rect 220726 288632 220782 288688
rect 220634 287816 220690 287872
rect 220726 287428 220782 287464
rect 220726 287408 220728 287428
rect 220728 287408 220780 287428
rect 220780 287408 220782 287428
rect 220634 286184 220690 286240
rect 220726 285776 220782 285832
rect 219162 49136 219218 49192
rect 218978 48320 219034 48376
rect 221554 51584 221610 51640
rect 221462 50224 221518 50280
rect 221646 49408 221702 49464
rect 226982 49272 227038 49328
rect 232502 51448 232558 51504
rect 234066 50496 234122 50552
rect 233882 50360 233938 50416
rect 229926 49544 229982 49600
rect 229742 48728 229798 48784
rect 231858 46280 231914 46336
rect 230478 42064 230534 42120
rect 240782 51176 240838 51232
rect 239402 50632 239458 50688
rect 240966 51312 241022 51368
rect 233422 6024 233478 6080
rect 246302 700304 246358 700360
rect 246302 48184 246358 48240
rect 243542 48048 243598 48104
rect 251270 645768 251326 645824
rect 251178 644544 251234 644600
rect 251178 643320 251234 643376
rect 251178 642096 251234 642152
rect 251178 640872 251234 640928
rect 251178 639648 251234 639704
rect 251178 638424 251234 638480
rect 250442 637200 250498 637256
rect 251178 635976 251234 636032
rect 251270 634752 251326 634808
rect 251178 633528 251234 633584
rect 251178 632304 251234 632360
rect 251178 631080 251234 631136
rect 251178 629856 251234 629912
rect 251178 628632 251234 628688
rect 251178 627408 251234 627464
rect 251178 626184 251234 626240
rect 251270 624960 251326 625016
rect 251178 623772 251180 623792
rect 251180 623772 251232 623792
rect 251232 623772 251234 623792
rect 251178 623736 251234 623772
rect 251178 622512 251234 622568
rect 251178 621288 251234 621344
rect 251178 620064 251234 620120
rect 251178 618840 251234 618896
rect 251178 617616 251234 617672
rect 251178 616392 251234 616448
rect 251178 615168 251234 615224
rect 251270 613944 251326 614000
rect 251178 612756 251180 612776
rect 251180 612756 251232 612776
rect 251232 612756 251234 612776
rect 251178 612720 251234 612756
rect 251178 611496 251234 611552
rect 251178 610272 251234 610328
rect 251178 609048 251234 609104
rect 251178 607824 251234 607880
rect 250534 606600 250590 606656
rect 251178 605376 251234 605432
rect 251178 604152 251234 604208
rect 251270 601724 251326 601760
rect 251270 601704 251272 601724
rect 251272 601704 251324 601724
rect 251324 601704 251326 601724
rect 251178 600480 251234 600536
rect 251178 599256 251234 599312
rect 251178 598032 251234 598088
rect 251178 595584 251234 595640
rect 251178 594360 251234 594416
rect 251178 593136 251234 593192
rect 251270 591912 251326 591968
rect 251178 590724 251180 590744
rect 251180 590724 251232 590744
rect 251232 590724 251234 590744
rect 251178 590688 251234 590724
rect 251178 589464 251234 589520
rect 251178 588240 251234 588296
rect 250626 587016 250682 587072
rect 251178 585792 251234 585848
rect 251178 584568 251234 584624
rect 251178 583344 251234 583400
rect 251178 582120 251234 582176
rect 251178 580896 251234 580952
rect 251270 579708 251272 579728
rect 251272 579708 251324 579728
rect 251324 579708 251326 579728
rect 251270 579672 251326 579708
rect 251178 578448 251234 578504
rect 251270 577224 251326 577280
rect 251178 576000 251234 576056
rect 251178 574776 251234 574832
rect 251178 573552 251234 573608
rect 251178 572328 251234 572384
rect 251178 571104 251234 571160
rect 251270 569880 251326 569936
rect 251178 568656 251234 568712
rect 251178 567432 251234 567488
rect 251178 566208 251234 566264
rect 251178 564984 251234 565040
rect 251178 563760 251234 563816
rect 251178 562536 251234 562592
rect 251178 561312 251234 561368
rect 251178 560088 251234 560144
rect 251270 558864 251326 558920
rect 251178 557660 251234 557696
rect 251178 557640 251180 557660
rect 251180 557640 251232 557660
rect 251232 557640 251234 557660
rect 251178 556416 251234 556472
rect 251178 555192 251234 555248
rect 251178 553968 251234 554024
rect 251178 552744 251234 552800
rect 251178 551520 251234 551576
rect 251178 550296 251234 550352
rect 251270 549072 251326 549128
rect 251178 547884 251180 547904
rect 251180 547884 251232 547904
rect 251232 547884 251234 547904
rect 251178 547848 251234 547884
rect 251178 546624 251234 546680
rect 251178 545400 251234 545456
rect 251178 544176 251234 544232
rect 250718 542952 250774 543008
rect 251178 541728 251234 541784
rect 251178 540504 251234 540560
rect 251178 539280 251234 539336
rect 251178 538056 251234 538112
rect 251178 535608 251234 535664
rect 251178 534384 251234 534440
rect 251178 496168 251234 496224
rect 251178 494944 251234 495000
rect 251178 493720 251234 493776
rect 251178 492496 251234 492552
rect 250810 491272 250866 491328
rect 251178 490048 251234 490104
rect 251178 488824 251234 488880
rect 251178 487600 251234 487656
rect 251178 486376 251234 486432
rect 251178 485152 251234 485208
rect 251178 483928 251234 483984
rect 251178 482704 251234 482760
rect 251178 481480 251234 481536
rect 251178 479032 251234 479088
rect 251178 477808 251234 477864
rect 251178 476584 251234 476640
rect 251178 475360 251234 475416
rect 251178 474136 251234 474192
rect 251178 472912 251234 472968
rect 251178 471688 251234 471744
rect 251270 470464 251326 470520
rect 251178 469276 251180 469296
rect 251180 469276 251232 469296
rect 251232 469276 251234 469296
rect 251178 469240 251234 469276
rect 251178 466792 251234 466848
rect 251638 465568 251694 465624
rect 251178 464344 251234 464400
rect 251178 463120 251234 463176
rect 251178 460672 251234 460728
rect 251178 459448 251234 459504
rect 251178 457000 251234 457056
rect 251178 455776 251234 455832
rect 251178 454552 251234 454608
rect 251730 453328 251786 453384
rect 251178 452104 251234 452160
rect 251178 450880 251234 450936
rect 251178 449656 251234 449712
rect 251178 447208 251234 447264
rect 251178 445984 251234 446040
rect 251178 444760 251234 444816
rect 250902 443536 250958 443592
rect 251178 442312 251234 442368
rect 251178 441088 251234 441144
rect 251178 439864 251234 439920
rect 251178 438640 251234 438696
rect 251270 437416 251326 437472
rect 251178 436212 251234 436248
rect 251178 436192 251180 436212
rect 251180 436192 251232 436212
rect 251232 436192 251234 436212
rect 251178 434968 251234 435024
rect 251178 433744 251234 433800
rect 251178 432520 251234 432576
rect 251178 431296 251234 431352
rect 251178 430072 251234 430128
rect 251178 428848 251234 428904
rect 251270 427624 251326 427680
rect 251178 426436 251180 426456
rect 251180 426436 251232 426456
rect 251232 426436 251234 426456
rect 251178 426400 251234 426436
rect 251178 425176 251234 425232
rect 251178 423952 251234 424008
rect 250994 422728 251050 422784
rect 251178 421504 251234 421560
rect 251178 420280 251234 420336
rect 251178 419056 251234 419112
rect 251178 417832 251234 417888
rect 251270 416608 251326 416664
rect 251178 415420 251180 415440
rect 251180 415420 251232 415440
rect 251232 415420 251234 415440
rect 251178 415384 251234 415420
rect 251178 414160 251234 414216
rect 251178 412936 251234 412992
rect 251178 411712 251234 411768
rect 251178 410488 251234 410544
rect 251178 409264 251234 409320
rect 251178 408040 251234 408096
rect 251638 406816 251694 406872
rect 251178 405592 251234 405648
rect 251086 403144 251142 403200
rect 251178 401920 251234 401976
rect 251730 404368 251786 404424
rect 251178 399472 251234 399528
rect 251178 398248 251234 398304
rect 251178 397024 251234 397080
rect 251178 395800 251234 395856
rect 251638 394576 251694 394632
rect 251178 393372 251234 393408
rect 251178 393352 251180 393372
rect 251180 393352 251232 393372
rect 251232 393352 251234 393372
rect 251178 392128 251234 392184
rect 251178 390904 251234 390960
rect 251178 389680 251234 389736
rect 251454 388456 251510 388512
rect 251730 387232 251786 387288
rect 251454 386008 251510 386064
rect 251178 384784 251234 384840
rect 251178 383560 251234 383616
rect 249246 50904 249302 50960
rect 249062 50768 249118 50824
rect 251914 602928 251970 602984
rect 252098 596808 252154 596864
rect 252006 533160 252062 533216
rect 251914 400696 251970 400752
rect 252190 536832 252246 536888
rect 252374 480256 252430 480312
rect 252190 468016 252246 468072
rect 252098 458224 252154 458280
rect 252466 461896 252522 461952
rect 252374 448432 252430 448488
rect 559654 700304 559710 700360
rect 580170 697176 580226 697232
rect 580170 683848 580226 683904
rect 580538 644000 580594 644056
rect 580262 630808 580318 630864
rect 580170 617480 580226 617536
rect 253294 51040 253350 51096
rect 247038 43424 247094 43480
rect 251270 6840 251326 6896
rect 256698 310528 256754 310584
rect 256698 308488 256754 308544
rect 256790 306448 256846 306504
rect 256698 302368 256754 302424
rect 256698 300328 256754 300384
rect 256698 298288 256754 298344
rect 256698 296248 256754 296304
rect 256698 294208 256754 294264
rect 256698 292168 256754 292224
rect 256698 290128 256754 290184
rect 256698 288088 256754 288144
rect 257342 286048 257398 286104
rect 256698 281968 256754 282024
rect 256698 279928 256754 279984
rect 256698 277888 256754 277944
rect 256698 275848 256754 275904
rect 256698 273808 256754 273864
rect 256698 269728 256754 269784
rect 256698 265648 256754 265704
rect 256698 263608 256754 263664
rect 256698 261568 256754 261624
rect 256698 259528 256754 259584
rect 256698 257488 256754 257544
rect 256698 255448 256754 255504
rect 256698 253408 256754 253464
rect 256698 251368 256754 251424
rect 256698 249328 256754 249384
rect 256698 247288 256754 247344
rect 256698 245248 256754 245304
rect 256698 243208 256754 243264
rect 256698 241168 256754 241224
rect 256698 239128 256754 239184
rect 256698 237088 256754 237144
rect 257710 304408 257766 304464
rect 257618 284008 257674 284064
rect 257434 271768 257490 271824
rect 257802 267688 257858 267744
rect 257342 235048 257398 235104
rect 256698 233008 256754 233064
rect 256330 230968 256386 231024
rect 256698 228964 256700 228984
rect 256700 228964 256752 228984
rect 256752 228964 256754 228984
rect 256698 228928 256754 228964
rect 256698 226888 256754 226944
rect 256698 224884 256700 224904
rect 256700 224884 256752 224904
rect 256752 224884 256754 224904
rect 256698 224848 256754 224884
rect 256698 222808 256754 222864
rect 256698 220788 256754 220824
rect 256698 220768 256700 220788
rect 256700 220768 256752 220788
rect 256752 220768 256754 220788
rect 256698 218728 256754 218784
rect 256698 216688 256754 216744
rect 256698 214648 256754 214704
rect 256698 212608 256754 212664
rect 256698 210568 256754 210624
rect 256238 208528 256294 208584
rect 256698 206488 256754 206544
rect 256698 204448 256754 204504
rect 256698 202408 256754 202464
rect 256698 200368 256754 200424
rect 256698 198328 256754 198384
rect 256698 196288 256754 196344
rect 256698 194248 256754 194304
rect 256698 192208 256754 192264
rect 256698 190168 256754 190224
rect 256698 188128 256754 188184
rect 256698 186088 256754 186144
rect 256698 184048 256754 184104
rect 256698 182008 256754 182064
rect 256698 179968 256754 180024
rect 256698 177964 256700 177984
rect 256700 177964 256752 177984
rect 256752 177964 256754 177984
rect 256698 177928 256754 177964
rect 256698 175888 256754 175944
rect 256698 171808 256754 171864
rect 256698 169768 256754 169824
rect 256698 167728 256754 167784
rect 256698 165688 256754 165744
rect 256698 163648 256754 163704
rect 256698 161608 256754 161664
rect 256698 159568 256754 159624
rect 256698 155488 256754 155544
rect 256698 153448 256754 153504
rect 256698 151408 256754 151464
rect 256698 149368 256754 149424
rect 256698 147328 256754 147384
rect 256698 145288 256754 145344
rect 256698 143248 256754 143304
rect 256698 141208 256754 141264
rect 256698 139168 256754 139224
rect 256698 135088 256754 135144
rect 256698 133048 256754 133104
rect 256146 131008 256202 131064
rect 256698 128968 256754 129024
rect 256698 126948 256754 126984
rect 256698 126928 256700 126948
rect 256700 126928 256752 126948
rect 256752 126928 256754 126948
rect 256698 124888 256754 124944
rect 256698 120808 256754 120864
rect 256698 118768 256754 118824
rect 256698 116728 256754 116784
rect 256698 114688 256754 114744
rect 256698 112648 256754 112704
rect 256698 110608 256754 110664
rect 256698 108568 256754 108624
rect 256698 106528 256754 106584
rect 256698 104488 256754 104544
rect 256698 102448 256754 102504
rect 256698 100408 256754 100464
rect 256054 98368 256110 98424
rect 256698 96328 256754 96384
rect 256698 94288 256754 94344
rect 256698 92248 256754 92304
rect 256698 90208 256754 90264
rect 256698 88168 256754 88224
rect 256698 86128 256754 86184
rect 256698 84124 256700 84144
rect 256700 84124 256752 84144
rect 256752 84124 256754 84144
rect 256698 84088 256754 84124
rect 256698 82048 256754 82104
rect 256698 80028 256754 80064
rect 256698 80008 256700 80028
rect 256700 80008 256752 80028
rect 256752 80008 256754 80028
rect 256698 77968 256754 78024
rect 256698 75928 256754 75984
rect 256698 73888 256754 73944
rect 256698 71848 256754 71904
rect 256698 69808 256754 69864
rect 256698 67768 256754 67824
rect 256698 63688 256754 63744
rect 256698 61648 256754 61704
rect 256698 59608 256754 59664
rect 256698 57568 256754 57624
rect 256698 55528 256754 55584
rect 257802 173848 257858 173904
rect 257434 157528 257490 157584
rect 257526 137128 257582 137184
rect 257434 65728 257490 65784
rect 257342 53488 257398 53544
rect 256698 51448 256754 51504
rect 256698 49408 256754 49464
rect 260102 46144 260158 46200
rect 550086 41112 550142 41168
rect 266358 36488 266414 36544
rect 285678 35536 285734 35592
rect 260654 3984 260710 4040
rect 264978 13504 265034 13560
rect 264150 3848 264206 3904
rect 268382 13368 268438 13424
rect 267738 3712 267794 3768
rect 271142 14728 271198 14784
rect 278318 3576 278374 3632
rect 284298 24384 284354 24440
rect 283102 13232 283158 13288
rect 284390 17584 284446 17640
rect 318798 37848 318854 37904
rect 303618 34176 303674 34232
rect 300858 18536 300914 18592
rect 303158 6704 303214 6760
rect 320178 29824 320234 29880
rect 318062 13096 318118 13152
rect 322110 14592 322166 14648
rect 338118 29688 338174 29744
rect 336738 21800 336794 21856
rect 353298 21664 353354 21720
rect 355230 15952 355286 16008
rect 356334 6568 356390 6624
rect 357530 32680 357586 32736
rect 371238 31048 371294 31104
rect 370594 6432 370650 6488
rect 373998 28464 374054 28520
rect 374090 21528 374146 21584
rect 552662 41248 552718 41304
rect 580170 537784 580226 537840
rect 580170 524476 580226 524512
rect 580170 524456 580172 524476
rect 580172 524456 580224 524476
rect 580224 524456 580226 524476
rect 580170 511264 580226 511320
rect 580170 458088 580226 458144
rect 579802 378392 579858 378448
rect 579986 365064 580042 365120
rect 580170 351908 580172 351928
rect 580172 351908 580224 351928
rect 580224 351908 580226 351928
rect 580170 351872 580226 351908
rect 580170 325216 580226 325272
rect 580446 590960 580502 591016
rect 580354 577632 580410 577688
rect 580630 564304 580686 564360
rect 580538 484608 580594 484664
rect 580630 471416 580686 471472
rect 580722 431568 580778 431624
rect 580814 418240 580870 418296
rect 580906 404912 580962 404968
rect 580446 312024 580502 312080
rect 580262 298696 580318 298752
rect 580170 272176 580226 272232
rect 580170 258848 580226 258904
rect 579618 232328 579674 232384
rect 580170 219000 580226 219056
rect 580170 179152 580226 179208
rect 579986 152632 580042 152688
rect 580170 139304 580226 139360
rect 580170 112784 580226 112840
rect 580170 72936 580226 72992
rect 580078 59608 580134 59664
rect 580354 245520 580410 245576
rect 580446 205672 580502 205728
rect 580538 192480 580594 192536
rect 580630 165824 580686 165880
rect 580722 125976 580778 126032
rect 580814 99456 580870 99512
rect 580906 86128 580962 86184
rect 580814 46280 580870 46336
rect 580630 41928 580686 41984
rect 390558 35400 390614 35456
rect 392582 12960 392638 13016
rect 407118 34040 407174 34096
rect 423678 29552 423734 29608
rect 407210 20032 407266 20088
rect 410798 14456 410854 14512
rect 409602 6296 409658 6352
rect 445758 26968 445814 27024
rect 426438 21392 426494 21448
rect 423770 4936 423826 4992
rect 428462 15816 428518 15872
rect 442998 19896 443054 19952
rect 445022 9016 445078 9072
rect 462318 12008 462374 12064
rect 463698 17448 463754 17504
rect 468666 3304 468722 3360
rect 477498 17312 477554 17368
rect 481730 6160 481786 6216
rect 498198 35264 498254 35320
rect 496818 24248 496874 24304
rect 495438 10240 495494 10296
rect 498290 26832 498346 26888
rect 514758 33904 514814 33960
rect 513378 28328 513434 28384
rect 532698 33768 532754 33824
rect 516138 28192 516194 28248
rect 514850 17176 514906 17232
rect 519542 3440 519598 3496
rect 531318 30912 531374 30968
rect 531410 11872 531466 11928
rect 534446 11736 534502 11792
rect 549258 35128 549314 35184
rect 550638 32544 550694 32600
rect 552018 32408 552074 32464
rect 549074 8880 549130 8936
rect 569958 25608 570014 25664
rect 568578 24112 568634 24168
rect 567566 11600 567622 11656
rect 566830 4800 566886 4856
rect 580354 33088 580410 33144
rect 580998 25472 581054 25528
rect 580262 19760 580318 19816
rect 580170 6568 580226 6624
rect 581090 21256 581146 21312
<< metal3 >>
rect 246297 700362 246363 700365
rect 559649 700362 559715 700365
rect 246297 700360 559715 700362
rect 246297 700304 246302 700360
rect 246358 700304 559654 700360
rect 559710 700304 559715 700360
rect 246297 700302 559715 700304
rect 246297 700299 246363 700302
rect 559649 700299 559715 700302
rect -960 697220 480 697460
rect 580165 697234 580231 697237
rect 583520 697234 584960 697324
rect 580165 697232 584960 697234
rect 580165 697176 580170 697232
rect 580226 697176 584960 697232
rect 580165 697174 584960 697176
rect 580165 697171 580231 697174
rect 583520 697084 584960 697174
rect -960 684314 480 684404
rect 3417 684314 3483 684317
rect -960 684312 3483 684314
rect -960 684256 3422 684312
rect 3478 684256 3483 684312
rect -960 684254 3483 684256
rect -960 684164 480 684254
rect 3417 684251 3483 684254
rect 580165 683906 580231 683909
rect 583520 683906 584960 683996
rect 580165 683904 584960 683906
rect 580165 683848 580170 683904
rect 580226 683848 584960 683904
rect 580165 683846 584960 683848
rect 580165 683843 580231 683846
rect 583520 683756 584960 683846
rect -960 671258 480 671348
rect 3509 671258 3575 671261
rect -960 671256 3575 671258
rect -960 671200 3514 671256
rect 3570 671200 3575 671256
rect -960 671198 3575 671200
rect -960 671108 480 671198
rect 3509 671195 3575 671198
rect 251766 670652 251772 670716
rect 251836 670714 251842 670716
rect 583520 670714 584960 670804
rect 251836 670654 584960 670714
rect 251836 670652 251842 670654
rect 583520 670564 584960 670654
rect -960 658202 480 658292
rect 3417 658202 3483 658205
rect -960 658200 3483 658202
rect -960 658144 3422 658200
rect 3478 658144 3483 658200
rect -960 658142 3483 658144
rect -960 658052 480 658142
rect 3417 658139 3483 658142
rect 583520 657236 584960 657476
rect 251265 645826 251331 645829
rect 251265 645824 253644 645826
rect 251265 645768 251270 645824
rect 251326 645768 253644 645824
rect 251265 645766 253644 645768
rect 251265 645763 251331 645766
rect -960 644996 480 645236
rect 251173 644602 251239 644605
rect 251173 644600 253644 644602
rect 251173 644544 251178 644600
rect 251234 644544 253644 644600
rect 251173 644542 253644 644544
rect 251173 644539 251239 644542
rect 580533 644058 580599 644061
rect 583520 644058 584960 644148
rect 580533 644056 584960 644058
rect 580533 644000 580538 644056
rect 580594 644000 584960 644056
rect 580533 643998 584960 644000
rect 580533 643995 580599 643998
rect 583520 643908 584960 643998
rect 251173 643378 251239 643381
rect 251173 643376 253644 643378
rect 251173 643320 251178 643376
rect 251234 643320 253644 643376
rect 251173 643318 253644 643320
rect 251173 643315 251239 643318
rect 251173 642154 251239 642157
rect 251173 642152 253644 642154
rect 251173 642096 251178 642152
rect 251234 642096 253644 642152
rect 251173 642094 253644 642096
rect 251173 642091 251239 642094
rect 251173 640930 251239 640933
rect 251173 640928 253644 640930
rect 251173 640872 251178 640928
rect 251234 640872 253644 640928
rect 251173 640870 253644 640872
rect 251173 640867 251239 640870
rect 251173 639706 251239 639709
rect 251173 639704 253644 639706
rect 251173 639648 251178 639704
rect 251234 639648 253644 639704
rect 251173 639646 253644 639648
rect 251173 639643 251239 639646
rect 251173 638482 251239 638485
rect 251173 638480 253644 638482
rect 251173 638424 251178 638480
rect 251234 638424 253644 638480
rect 251173 638422 253644 638424
rect 251173 638419 251239 638422
rect 250437 637258 250503 637261
rect 250437 637256 253644 637258
rect 250437 637200 250442 637256
rect 250498 637200 253644 637256
rect 250437 637198 253644 637200
rect 250437 637195 250503 637198
rect 251173 636034 251239 636037
rect 251173 636032 253644 636034
rect 251173 635976 251178 636032
rect 251234 635976 253644 636032
rect 251173 635974 253644 635976
rect 251173 635971 251239 635974
rect 251265 634810 251331 634813
rect 251265 634808 253644 634810
rect 251265 634752 251270 634808
rect 251326 634752 253644 634808
rect 251265 634750 253644 634752
rect 251265 634747 251331 634750
rect 251173 633586 251239 633589
rect 251173 633584 253644 633586
rect 251173 633528 251178 633584
rect 251234 633528 253644 633584
rect 251173 633526 253644 633528
rect 251173 633523 251239 633526
rect 251173 632362 251239 632365
rect 251173 632360 253644 632362
rect 251173 632304 251178 632360
rect 251234 632304 253644 632360
rect 251173 632302 253644 632304
rect 251173 632299 251239 632302
rect -960 632090 480 632180
rect 3417 632090 3483 632093
rect -960 632088 3483 632090
rect -960 632032 3422 632088
rect 3478 632032 3483 632088
rect -960 632030 3483 632032
rect -960 631940 480 632030
rect 3417 632027 3483 632030
rect 251173 631138 251239 631141
rect 251173 631136 253644 631138
rect 251173 631080 251178 631136
rect 251234 631080 253644 631136
rect 251173 631078 253644 631080
rect 251173 631075 251239 631078
rect 580257 630866 580323 630869
rect 583520 630866 584960 630956
rect 580257 630864 584960 630866
rect 580257 630808 580262 630864
rect 580318 630808 584960 630864
rect 580257 630806 584960 630808
rect 580257 630803 580323 630806
rect 583520 630716 584960 630806
rect 251173 629914 251239 629917
rect 251173 629912 253644 629914
rect 251173 629856 251178 629912
rect 251234 629856 253644 629912
rect 251173 629854 253644 629856
rect 251173 629851 251239 629854
rect 251173 628690 251239 628693
rect 251173 628688 253644 628690
rect 251173 628632 251178 628688
rect 251234 628632 253644 628688
rect 251173 628630 253644 628632
rect 251173 628627 251239 628630
rect 251173 627466 251239 627469
rect 251173 627464 253644 627466
rect 251173 627408 251178 627464
rect 251234 627408 253644 627464
rect 251173 627406 253644 627408
rect 251173 627403 251239 627406
rect 251173 626242 251239 626245
rect 251173 626240 253644 626242
rect 251173 626184 251178 626240
rect 251234 626184 253644 626240
rect 251173 626182 253644 626184
rect 251173 626179 251239 626182
rect 251265 625018 251331 625021
rect 251265 625016 253644 625018
rect 251265 624960 251270 625016
rect 251326 624960 253644 625016
rect 251265 624958 253644 624960
rect 251265 624955 251331 624958
rect 251173 623794 251239 623797
rect 251173 623792 253644 623794
rect 251173 623736 251178 623792
rect 251234 623736 253644 623792
rect 251173 623734 253644 623736
rect 251173 623731 251239 623734
rect 251173 622570 251239 622573
rect 251173 622568 253644 622570
rect 251173 622512 251178 622568
rect 251234 622512 253644 622568
rect 251173 622510 253644 622512
rect 251173 622507 251239 622510
rect 251173 621346 251239 621349
rect 251173 621344 253644 621346
rect 251173 621288 251178 621344
rect 251234 621288 253644 621344
rect 251173 621286 253644 621288
rect 251173 621283 251239 621286
rect 251173 620122 251239 620125
rect 251173 620120 253644 620122
rect 251173 620064 251178 620120
rect 251234 620064 253644 620120
rect 251173 620062 253644 620064
rect 251173 620059 251239 620062
rect -960 619170 480 619260
rect 3141 619170 3207 619173
rect -960 619168 3207 619170
rect -960 619112 3146 619168
rect 3202 619112 3207 619168
rect -960 619110 3207 619112
rect -960 619020 480 619110
rect 3141 619107 3207 619110
rect 251173 618898 251239 618901
rect 251173 618896 253644 618898
rect 251173 618840 251178 618896
rect 251234 618840 253644 618896
rect 251173 618838 253644 618840
rect 251173 618835 251239 618838
rect 251173 617674 251239 617677
rect 251173 617672 253644 617674
rect 251173 617616 251178 617672
rect 251234 617616 253644 617672
rect 251173 617614 253644 617616
rect 251173 617611 251239 617614
rect 580165 617538 580231 617541
rect 583520 617538 584960 617628
rect 580165 617536 584960 617538
rect 580165 617480 580170 617536
rect 580226 617480 584960 617536
rect 580165 617478 584960 617480
rect 580165 617475 580231 617478
rect 583520 617388 584960 617478
rect 251173 616450 251239 616453
rect 251173 616448 253644 616450
rect 251173 616392 251178 616448
rect 251234 616392 253644 616448
rect 251173 616390 253644 616392
rect 251173 616387 251239 616390
rect 251173 615226 251239 615229
rect 251173 615224 253644 615226
rect 251173 615168 251178 615224
rect 251234 615168 253644 615224
rect 251173 615166 253644 615168
rect 251173 615163 251239 615166
rect 251265 614002 251331 614005
rect 251265 614000 253644 614002
rect 251265 613944 251270 614000
rect 251326 613944 253644 614000
rect 251265 613942 253644 613944
rect 251265 613939 251331 613942
rect 251173 612778 251239 612781
rect 251173 612776 253644 612778
rect 251173 612720 251178 612776
rect 251234 612720 253644 612776
rect 251173 612718 253644 612720
rect 251173 612715 251239 612718
rect 251173 611554 251239 611557
rect 251173 611552 253644 611554
rect 251173 611496 251178 611552
rect 251234 611496 253644 611552
rect 251173 611494 253644 611496
rect 251173 611491 251239 611494
rect 251173 610330 251239 610333
rect 251173 610328 253644 610330
rect 251173 610272 251178 610328
rect 251234 610272 253644 610328
rect 251173 610270 253644 610272
rect 251173 610267 251239 610270
rect 251173 609106 251239 609109
rect 251173 609104 253644 609106
rect 251173 609048 251178 609104
rect 251234 609048 253644 609104
rect 251173 609046 253644 609048
rect 251173 609043 251239 609046
rect 251173 607882 251239 607885
rect 251173 607880 253644 607882
rect 251173 607824 251178 607880
rect 251234 607824 253644 607880
rect 251173 607822 253644 607824
rect 251173 607819 251239 607822
rect 250529 606658 250595 606661
rect 250529 606656 253644 606658
rect 250529 606600 250534 606656
rect 250590 606600 253644 606656
rect 250529 606598 253644 606600
rect 250529 606595 250595 606598
rect -960 606114 480 606204
rect 3233 606114 3299 606117
rect -960 606112 3299 606114
rect -960 606056 3238 606112
rect 3294 606056 3299 606112
rect -960 606054 3299 606056
rect -960 605964 480 606054
rect 3233 606051 3299 606054
rect 251173 605434 251239 605437
rect 251173 605432 253644 605434
rect 251173 605376 251178 605432
rect 251234 605376 253644 605432
rect 251173 605374 253644 605376
rect 251173 605371 251239 605374
rect 251173 604210 251239 604213
rect 251173 604208 253644 604210
rect 251173 604152 251178 604208
rect 251234 604152 253644 604208
rect 251173 604150 253644 604152
rect 251173 604147 251239 604150
rect 583520 604060 584960 604300
rect 251909 602986 251975 602989
rect 251909 602984 253644 602986
rect 251909 602928 251914 602984
rect 251970 602928 253644 602984
rect 251909 602926 253644 602928
rect 251909 602923 251975 602926
rect 251265 601762 251331 601765
rect 251265 601760 253644 601762
rect 251265 601704 251270 601760
rect 251326 601704 253644 601760
rect 251265 601702 253644 601704
rect 251265 601699 251331 601702
rect 251173 600538 251239 600541
rect 251173 600536 253644 600538
rect 251173 600480 251178 600536
rect 251234 600480 253644 600536
rect 251173 600478 253644 600480
rect 251173 600475 251239 600478
rect 251173 599314 251239 599317
rect 251173 599312 253644 599314
rect 251173 599256 251178 599312
rect 251234 599256 253644 599312
rect 251173 599254 253644 599256
rect 251173 599251 251239 599254
rect 251173 598090 251239 598093
rect 251173 598088 253644 598090
rect 251173 598032 251178 598088
rect 251234 598032 253644 598088
rect 251173 598030 253644 598032
rect 251173 598027 251239 598030
rect 252093 596866 252159 596869
rect 252093 596864 253644 596866
rect 252093 596808 252098 596864
rect 252154 596808 253644 596864
rect 252093 596806 253644 596808
rect 252093 596803 252159 596806
rect 251173 595642 251239 595645
rect 251173 595640 253644 595642
rect 251173 595584 251178 595640
rect 251234 595584 253644 595640
rect 251173 595582 253644 595584
rect 251173 595579 251239 595582
rect 251173 594418 251239 594421
rect 251173 594416 253644 594418
rect 251173 594360 251178 594416
rect 251234 594360 253644 594416
rect 251173 594358 253644 594360
rect 251173 594355 251239 594358
rect 251173 593194 251239 593197
rect 251173 593192 253644 593194
rect -960 592908 480 593148
rect 251173 593136 251178 593192
rect 251234 593136 253644 593192
rect 251173 593134 253644 593136
rect 251173 593131 251239 593134
rect 251265 591970 251331 591973
rect 251265 591968 253644 591970
rect 251265 591912 251270 591968
rect 251326 591912 253644 591968
rect 251265 591910 253644 591912
rect 251265 591907 251331 591910
rect 111885 591698 111951 591701
rect 109940 591696 111951 591698
rect 109940 591640 111890 591696
rect 111946 591640 111951 591696
rect 109940 591638 111951 591640
rect 111885 591635 111951 591638
rect 111793 591018 111859 591021
rect 109940 591016 111859 591018
rect 109940 590960 111798 591016
rect 111854 590960 111859 591016
rect 109940 590958 111859 590960
rect 111793 590955 111859 590958
rect 580441 591018 580507 591021
rect 583520 591018 584960 591108
rect 580441 591016 584960 591018
rect 580441 590960 580446 591016
rect 580502 590960 584960 591016
rect 580441 590958 584960 590960
rect 580441 590955 580507 590958
rect 583520 590868 584960 590958
rect 251173 590746 251239 590749
rect 251173 590744 253644 590746
rect 251173 590688 251178 590744
rect 251234 590688 253644 590744
rect 251173 590686 253644 590688
rect 251173 590683 251239 590686
rect 111885 590338 111951 590341
rect 109940 590336 111951 590338
rect 109940 590280 111890 590336
rect 111946 590280 111951 590336
rect 109940 590278 111951 590280
rect 111885 590275 111951 590278
rect 111793 589658 111859 589661
rect 109940 589656 111859 589658
rect 109940 589600 111798 589656
rect 111854 589600 111859 589656
rect 109940 589598 111859 589600
rect 111793 589595 111859 589598
rect 251173 589522 251239 589525
rect 251173 589520 253644 589522
rect 251173 589464 251178 589520
rect 251234 589464 253644 589520
rect 251173 589462 253644 589464
rect 251173 589459 251239 589462
rect 111793 588978 111859 588981
rect 109940 588976 111859 588978
rect 109940 588920 111798 588976
rect 111854 588920 111859 588976
rect 109940 588918 111859 588920
rect 111793 588915 111859 588918
rect 112253 588298 112319 588301
rect 109940 588296 112319 588298
rect 109940 588240 112258 588296
rect 112314 588240 112319 588296
rect 109940 588238 112319 588240
rect 112253 588235 112319 588238
rect 251173 588298 251239 588301
rect 251173 588296 253644 588298
rect 251173 588240 251178 588296
rect 251234 588240 253644 588296
rect 251173 588238 253644 588240
rect 251173 588235 251239 588238
rect 111793 587618 111859 587621
rect 109940 587616 111859 587618
rect 109940 587560 111798 587616
rect 111854 587560 111859 587616
rect 109940 587558 111859 587560
rect 111793 587555 111859 587558
rect 250621 587074 250687 587077
rect 250621 587072 253644 587074
rect 250621 587016 250626 587072
rect 250682 587016 253644 587072
rect 250621 587014 253644 587016
rect 250621 587011 250687 587014
rect 112713 586938 112779 586941
rect 109940 586936 112779 586938
rect 109940 586880 112718 586936
rect 112774 586880 112779 586936
rect 109940 586878 112779 586880
rect 112713 586875 112779 586878
rect 111793 586258 111859 586261
rect 109940 586256 111859 586258
rect 109940 586200 111798 586256
rect 111854 586200 111859 586256
rect 109940 586198 111859 586200
rect 111793 586195 111859 586198
rect 251173 585850 251239 585853
rect 251173 585848 253644 585850
rect 251173 585792 251178 585848
rect 251234 585792 253644 585848
rect 251173 585790 253644 585792
rect 251173 585787 251239 585790
rect 111977 585578 112043 585581
rect 109940 585576 112043 585578
rect 109940 585520 111982 585576
rect 112038 585520 112043 585576
rect 109940 585518 112043 585520
rect 111977 585515 112043 585518
rect 111885 584898 111951 584901
rect 109940 584896 111951 584898
rect 109940 584840 111890 584896
rect 111946 584840 111951 584896
rect 109940 584838 111951 584840
rect 111885 584835 111951 584838
rect 251173 584626 251239 584629
rect 251173 584624 253644 584626
rect 251173 584568 251178 584624
rect 251234 584568 253644 584624
rect 251173 584566 253644 584568
rect 251173 584563 251239 584566
rect 111793 584218 111859 584221
rect 109940 584216 111859 584218
rect 109940 584160 111798 584216
rect 111854 584160 111859 584216
rect 109940 584158 111859 584160
rect 111793 584155 111859 584158
rect 111793 583538 111859 583541
rect 109940 583536 111859 583538
rect 109940 583480 111798 583536
rect 111854 583480 111859 583536
rect 109940 583478 111859 583480
rect 111793 583475 111859 583478
rect 251173 583402 251239 583405
rect 251173 583400 253644 583402
rect 251173 583344 251178 583400
rect 251234 583344 253644 583400
rect 251173 583342 253644 583344
rect 251173 583339 251239 583342
rect 111885 582858 111951 582861
rect 109940 582856 111951 582858
rect 109940 582800 111890 582856
rect 111946 582800 111951 582856
rect 109940 582798 111951 582800
rect 111885 582795 111951 582798
rect 111793 582178 111859 582181
rect 109940 582176 111859 582178
rect 109940 582120 111798 582176
rect 111854 582120 111859 582176
rect 109940 582118 111859 582120
rect 111793 582115 111859 582118
rect 251173 582178 251239 582181
rect 251173 582176 253644 582178
rect 251173 582120 251178 582176
rect 251234 582120 253644 582176
rect 251173 582118 253644 582120
rect 251173 582115 251239 582118
rect 111977 581498 112043 581501
rect 109940 581496 112043 581498
rect 109940 581440 111982 581496
rect 112038 581440 112043 581496
rect 109940 581438 112043 581440
rect 111977 581435 112043 581438
rect 251173 580954 251239 580957
rect 251173 580952 253644 580954
rect 251173 580896 251178 580952
rect 251234 580896 253644 580952
rect 251173 580894 253644 580896
rect 251173 580891 251239 580894
rect 111885 580818 111951 580821
rect 109940 580816 111951 580818
rect 109940 580760 111890 580816
rect 111946 580760 111951 580816
rect 109940 580758 111951 580760
rect 111885 580755 111951 580758
rect 111793 580138 111859 580141
rect 109940 580136 111859 580138
rect -960 580002 480 580092
rect 109940 580080 111798 580136
rect 111854 580080 111859 580136
rect 109940 580078 111859 580080
rect 111793 580075 111859 580078
rect 3325 580002 3391 580005
rect -960 580000 3391 580002
rect -960 579944 3330 580000
rect 3386 579944 3391 580000
rect -960 579942 3391 579944
rect -960 579852 480 579942
rect 3325 579939 3391 579942
rect 251265 579730 251331 579733
rect 251265 579728 253644 579730
rect 251265 579672 251270 579728
rect 251326 579672 253644 579728
rect 251265 579670 253644 579672
rect 251265 579667 251331 579670
rect 111885 579458 111951 579461
rect 109940 579456 111951 579458
rect 109940 579400 111890 579456
rect 111946 579400 111951 579456
rect 109940 579398 111951 579400
rect 111885 579395 111951 579398
rect 111793 578778 111859 578781
rect 109940 578776 111859 578778
rect 109940 578720 111798 578776
rect 111854 578720 111859 578776
rect 109940 578718 111859 578720
rect 111793 578715 111859 578718
rect 251173 578506 251239 578509
rect 251173 578504 253644 578506
rect 251173 578448 251178 578504
rect 251234 578448 253644 578504
rect 251173 578446 253644 578448
rect 251173 578443 251239 578446
rect 111793 578098 111859 578101
rect 109940 578096 111859 578098
rect 109940 578040 111798 578096
rect 111854 578040 111859 578096
rect 109940 578038 111859 578040
rect 111793 578035 111859 578038
rect 580349 577690 580415 577693
rect 583520 577690 584960 577780
rect 580349 577688 584960 577690
rect 580349 577632 580354 577688
rect 580410 577632 584960 577688
rect 580349 577630 584960 577632
rect 580349 577627 580415 577630
rect 583520 577540 584960 577630
rect 112437 577418 112503 577421
rect 109940 577416 112503 577418
rect 109940 577360 112442 577416
rect 112498 577360 112503 577416
rect 109940 577358 112503 577360
rect 112437 577355 112503 577358
rect 251265 577282 251331 577285
rect 251265 577280 253644 577282
rect 251265 577224 251270 577280
rect 251326 577224 253644 577280
rect 251265 577222 253644 577224
rect 251265 577219 251331 577222
rect 111885 576738 111951 576741
rect 109940 576736 111951 576738
rect 109940 576680 111890 576736
rect 111946 576680 111951 576736
rect 109940 576678 111951 576680
rect 111885 576675 111951 576678
rect 111793 576058 111859 576061
rect 109940 576056 111859 576058
rect 109940 576000 111798 576056
rect 111854 576000 111859 576056
rect 109940 575998 111859 576000
rect 111793 575995 111859 575998
rect 251173 576058 251239 576061
rect 251173 576056 253644 576058
rect 251173 576000 251178 576056
rect 251234 576000 253644 576056
rect 251173 575998 253644 576000
rect 251173 575995 251239 575998
rect 111885 575378 111951 575381
rect 109940 575376 111951 575378
rect 109940 575320 111890 575376
rect 111946 575320 111951 575376
rect 109940 575318 111951 575320
rect 111885 575315 111951 575318
rect 251173 574834 251239 574837
rect 251173 574832 253644 574834
rect 251173 574776 251178 574832
rect 251234 574776 253644 574832
rect 251173 574774 253644 574776
rect 251173 574771 251239 574774
rect 111793 574698 111859 574701
rect 109940 574696 111859 574698
rect 109940 574640 111798 574696
rect 111854 574640 111859 574696
rect 109940 574638 111859 574640
rect 111793 574635 111859 574638
rect 111885 574018 111951 574021
rect 109940 574016 111951 574018
rect 109940 573960 111890 574016
rect 111946 573960 111951 574016
rect 109940 573958 111951 573960
rect 111885 573955 111951 573958
rect 251173 573610 251239 573613
rect 251173 573608 253644 573610
rect 251173 573552 251178 573608
rect 251234 573552 253644 573608
rect 251173 573550 253644 573552
rect 251173 573547 251239 573550
rect 111793 573338 111859 573341
rect 109940 573336 111859 573338
rect 109940 573280 111798 573336
rect 111854 573280 111859 573336
rect 109940 573278 111859 573280
rect 111793 573275 111859 573278
rect 111885 572658 111951 572661
rect 109940 572656 111951 572658
rect 109940 572600 111890 572656
rect 111946 572600 111951 572656
rect 109940 572598 111951 572600
rect 111885 572595 111951 572598
rect 251173 572386 251239 572389
rect 251173 572384 253644 572386
rect 251173 572328 251178 572384
rect 251234 572328 253644 572384
rect 251173 572326 253644 572328
rect 251173 572323 251239 572326
rect 111793 571978 111859 571981
rect 109940 571976 111859 571978
rect 109940 571920 111798 571976
rect 111854 571920 111859 571976
rect 109940 571918 111859 571920
rect 111793 571915 111859 571918
rect 111977 571298 112043 571301
rect 109940 571296 112043 571298
rect 109940 571240 111982 571296
rect 112038 571240 112043 571296
rect 109940 571238 112043 571240
rect 111977 571235 112043 571238
rect 251173 571162 251239 571165
rect 251173 571160 253644 571162
rect 251173 571104 251178 571160
rect 251234 571104 253644 571160
rect 251173 571102 253644 571104
rect 251173 571099 251239 571102
rect 111793 570618 111859 570621
rect 109940 570616 111859 570618
rect 109940 570560 111798 570616
rect 111854 570560 111859 570616
rect 109940 570558 111859 570560
rect 111793 570555 111859 570558
rect 111885 569938 111951 569941
rect 109940 569936 111951 569938
rect 109940 569880 111890 569936
rect 111946 569880 111951 569936
rect 109940 569878 111951 569880
rect 111885 569875 111951 569878
rect 251265 569938 251331 569941
rect 251265 569936 253644 569938
rect 251265 569880 251270 569936
rect 251326 569880 253644 569936
rect 251265 569878 253644 569880
rect 251265 569875 251331 569878
rect 111793 569258 111859 569261
rect 109940 569256 111859 569258
rect 109940 569200 111798 569256
rect 111854 569200 111859 569256
rect 109940 569198 111859 569200
rect 111793 569195 111859 569198
rect 251173 568714 251239 568717
rect 251173 568712 253644 568714
rect 251173 568656 251178 568712
rect 251234 568656 253644 568712
rect 251173 568654 253644 568656
rect 251173 568651 251239 568654
rect 111977 568578 112043 568581
rect 109940 568576 112043 568578
rect 109940 568520 111982 568576
rect 112038 568520 112043 568576
rect 109940 568518 112043 568520
rect 111977 568515 112043 568518
rect 112345 567898 112411 567901
rect 109940 567896 112411 567898
rect 109940 567840 112350 567896
rect 112406 567840 112411 567896
rect 109940 567838 112411 567840
rect 112345 567835 112411 567838
rect 251173 567490 251239 567493
rect 251173 567488 253644 567490
rect 251173 567432 251178 567488
rect 251234 567432 253644 567488
rect 251173 567430 253644 567432
rect 251173 567427 251239 567430
rect 111793 567218 111859 567221
rect 109940 567216 111859 567218
rect 109940 567160 111798 567216
rect 111854 567160 111859 567216
rect 109940 567158 111859 567160
rect 111793 567155 111859 567158
rect -960 566946 480 567036
rect 3417 566946 3483 566949
rect -960 566944 3483 566946
rect -960 566888 3422 566944
rect 3478 566888 3483 566944
rect -960 566886 3483 566888
rect -960 566796 480 566886
rect 3417 566883 3483 566886
rect 111885 566538 111951 566541
rect 109940 566536 111951 566538
rect 109940 566480 111890 566536
rect 111946 566480 111951 566536
rect 109940 566478 111951 566480
rect 111885 566475 111951 566478
rect 251173 566266 251239 566269
rect 251173 566264 253644 566266
rect 251173 566208 251178 566264
rect 251234 566208 253644 566264
rect 251173 566206 253644 566208
rect 251173 566203 251239 566206
rect 111793 565858 111859 565861
rect 109940 565856 111859 565858
rect 109940 565800 111798 565856
rect 111854 565800 111859 565856
rect 109940 565798 111859 565800
rect 111793 565795 111859 565798
rect 111885 565178 111951 565181
rect 109940 565176 111951 565178
rect 109940 565120 111890 565176
rect 111946 565120 111951 565176
rect 109940 565118 111951 565120
rect 111885 565115 111951 565118
rect 251173 565042 251239 565045
rect 251173 565040 253644 565042
rect 251173 564984 251178 565040
rect 251234 564984 253644 565040
rect 251173 564982 253644 564984
rect 251173 564979 251239 564982
rect 111793 564498 111859 564501
rect 109940 564496 111859 564498
rect 109940 564440 111798 564496
rect 111854 564440 111859 564496
rect 109940 564438 111859 564440
rect 111793 564435 111859 564438
rect 580625 564362 580691 564365
rect 583520 564362 584960 564452
rect 580625 564360 584960 564362
rect 580625 564304 580630 564360
rect 580686 564304 584960 564360
rect 580625 564302 584960 564304
rect 580625 564299 580691 564302
rect 583520 564212 584960 564302
rect 112989 563818 113055 563821
rect 109940 563816 113055 563818
rect 109940 563760 112994 563816
rect 113050 563760 113055 563816
rect 109940 563758 113055 563760
rect 112989 563755 113055 563758
rect 251173 563818 251239 563821
rect 251173 563816 253644 563818
rect 251173 563760 251178 563816
rect 251234 563760 253644 563816
rect 251173 563758 253644 563760
rect 251173 563755 251239 563758
rect 111793 563138 111859 563141
rect 109940 563136 111859 563138
rect 109940 563080 111798 563136
rect 111854 563080 111859 563136
rect 109940 563078 111859 563080
rect 111793 563075 111859 563078
rect 251173 562594 251239 562597
rect 251173 562592 253644 562594
rect 251173 562536 251178 562592
rect 251234 562536 253644 562592
rect 251173 562534 253644 562536
rect 251173 562531 251239 562534
rect 112621 562458 112687 562461
rect 109940 562456 112687 562458
rect 109940 562400 112626 562456
rect 112682 562400 112687 562456
rect 109940 562398 112687 562400
rect 112621 562395 112687 562398
rect 111793 561778 111859 561781
rect 109940 561776 111859 561778
rect 109940 561720 111798 561776
rect 111854 561720 111859 561776
rect 109940 561718 111859 561720
rect 111793 561715 111859 561718
rect 251173 561370 251239 561373
rect 251173 561368 253644 561370
rect 251173 561312 251178 561368
rect 251234 561312 253644 561368
rect 251173 561310 253644 561312
rect 251173 561307 251239 561310
rect 112437 561098 112503 561101
rect 109940 561096 112503 561098
rect 109940 561040 112442 561096
rect 112498 561040 112503 561096
rect 109940 561038 112503 561040
rect 112437 561035 112503 561038
rect 111793 560418 111859 560421
rect 109940 560416 111859 560418
rect 109940 560360 111798 560416
rect 111854 560360 111859 560416
rect 109940 560358 111859 560360
rect 111793 560355 111859 560358
rect 251173 560146 251239 560149
rect 251173 560144 253644 560146
rect 251173 560088 251178 560144
rect 251234 560088 253644 560144
rect 251173 560086 253644 560088
rect 251173 560083 251239 560086
rect 111885 559738 111951 559741
rect 109940 559736 111951 559738
rect 109940 559680 111890 559736
rect 111946 559680 111951 559736
rect 109940 559678 111951 559680
rect 111885 559675 111951 559678
rect 111793 559058 111859 559061
rect 109940 559056 111859 559058
rect 109940 559000 111798 559056
rect 111854 559000 111859 559056
rect 109940 558998 111859 559000
rect 111793 558995 111859 558998
rect 251265 558922 251331 558925
rect 251265 558920 253644 558922
rect 251265 558864 251270 558920
rect 251326 558864 253644 558920
rect 251265 558862 253644 558864
rect 251265 558859 251331 558862
rect 111885 558378 111951 558381
rect 109940 558376 111951 558378
rect 109940 558320 111890 558376
rect 111946 558320 111951 558376
rect 109940 558318 111951 558320
rect 111885 558315 111951 558318
rect 111793 557698 111859 557701
rect 109940 557696 111859 557698
rect 109940 557640 111798 557696
rect 111854 557640 111859 557696
rect 109940 557638 111859 557640
rect 111793 557635 111859 557638
rect 251173 557698 251239 557701
rect 251173 557696 253644 557698
rect 251173 557640 251178 557696
rect 251234 557640 253644 557696
rect 251173 557638 253644 557640
rect 251173 557635 251239 557638
rect 111793 557018 111859 557021
rect 109940 557016 111859 557018
rect 109940 556960 111798 557016
rect 111854 556960 111859 557016
rect 109940 556958 111859 556960
rect 111793 556955 111859 556958
rect 251173 556474 251239 556477
rect 251173 556472 253644 556474
rect 251173 556416 251178 556472
rect 251234 556416 253644 556472
rect 251173 556414 253644 556416
rect 251173 556411 251239 556414
rect 111977 556338 112043 556341
rect 109940 556336 112043 556338
rect 109940 556280 111982 556336
rect 112038 556280 112043 556336
rect 109940 556278 112043 556280
rect 111977 556275 112043 556278
rect 111885 555658 111951 555661
rect 109940 555656 111951 555658
rect 109940 555600 111890 555656
rect 111946 555600 111951 555656
rect 109940 555598 111951 555600
rect 111885 555595 111951 555598
rect 251173 555250 251239 555253
rect 251173 555248 253644 555250
rect 251173 555192 251178 555248
rect 251234 555192 253644 555248
rect 251173 555190 253644 555192
rect 251173 555187 251239 555190
rect 111793 554978 111859 554981
rect 109940 554976 111859 554978
rect 109940 554920 111798 554976
rect 111854 554920 111859 554976
rect 109940 554918 111859 554920
rect 111793 554915 111859 554918
rect 112069 554298 112135 554301
rect 109940 554296 112135 554298
rect 109940 554240 112074 554296
rect 112130 554240 112135 554296
rect 109940 554238 112135 554240
rect 112069 554235 112135 554238
rect 251173 554026 251239 554029
rect 251173 554024 253644 554026
rect -960 553890 480 553980
rect 251173 553968 251178 554024
rect 251234 553968 253644 554024
rect 251173 553966 253644 553968
rect 251173 553963 251239 553966
rect 3417 553890 3483 553893
rect -960 553888 3483 553890
rect -960 553832 3422 553888
rect 3478 553832 3483 553888
rect -960 553830 3483 553832
rect -960 553740 480 553830
rect 3417 553827 3483 553830
rect 111793 553618 111859 553621
rect 109940 553616 111859 553618
rect 109940 553560 111798 553616
rect 111854 553560 111859 553616
rect 109940 553558 111859 553560
rect 111793 553555 111859 553558
rect 111885 552938 111951 552941
rect 109940 552936 111951 552938
rect 109940 552880 111890 552936
rect 111946 552880 111951 552936
rect 109940 552878 111951 552880
rect 111885 552875 111951 552878
rect 251173 552802 251239 552805
rect 251173 552800 253644 552802
rect 251173 552744 251178 552800
rect 251234 552744 253644 552800
rect 251173 552742 253644 552744
rect 251173 552739 251239 552742
rect 111793 552258 111859 552261
rect 109940 552256 111859 552258
rect 109940 552200 111798 552256
rect 111854 552200 111859 552256
rect 109940 552198 111859 552200
rect 111793 552195 111859 552198
rect 111885 551578 111951 551581
rect 109940 551576 111951 551578
rect 109940 551520 111890 551576
rect 111946 551520 111951 551576
rect 109940 551518 111951 551520
rect 111885 551515 111951 551518
rect 251173 551578 251239 551581
rect 251173 551576 253644 551578
rect 251173 551520 251178 551576
rect 251234 551520 253644 551576
rect 251173 551518 253644 551520
rect 251173 551515 251239 551518
rect 583520 551020 584960 551260
rect 111793 550898 111859 550901
rect 109940 550896 111859 550898
rect 109940 550840 111798 550896
rect 111854 550840 111859 550896
rect 109940 550838 111859 550840
rect 111793 550835 111859 550838
rect 251173 550354 251239 550357
rect 251173 550352 253644 550354
rect 251173 550296 251178 550352
rect 251234 550296 253644 550352
rect 251173 550294 253644 550296
rect 251173 550291 251239 550294
rect 111885 550218 111951 550221
rect 109940 550216 111951 550218
rect 109940 550160 111890 550216
rect 111946 550160 111951 550216
rect 109940 550158 111951 550160
rect 111885 550155 111951 550158
rect 111793 549538 111859 549541
rect 109940 549536 111859 549538
rect 109940 549480 111798 549536
rect 111854 549480 111859 549536
rect 109940 549478 111859 549480
rect 111793 549475 111859 549478
rect 251265 549130 251331 549133
rect 251265 549128 253644 549130
rect 251265 549072 251270 549128
rect 251326 549072 253644 549128
rect 251265 549070 253644 549072
rect 251265 549067 251331 549070
rect 111885 548858 111951 548861
rect 109940 548856 111951 548858
rect 109940 548800 111890 548856
rect 111946 548800 111951 548856
rect 109940 548798 111951 548800
rect 111885 548795 111951 548798
rect 111793 548178 111859 548181
rect 109940 548176 111859 548178
rect 109940 548120 111798 548176
rect 111854 548120 111859 548176
rect 109940 548118 111859 548120
rect 111793 548115 111859 548118
rect 251173 547906 251239 547909
rect 251173 547904 253644 547906
rect 251173 547848 251178 547904
rect 251234 547848 253644 547904
rect 251173 547846 253644 547848
rect 251173 547843 251239 547846
rect 112805 547498 112871 547501
rect 109940 547496 112871 547498
rect 109940 547440 112810 547496
rect 112866 547440 112871 547496
rect 109940 547438 112871 547440
rect 112805 547435 112871 547438
rect 111793 546818 111859 546821
rect 109940 546816 111859 546818
rect 109940 546760 111798 546816
rect 111854 546760 111859 546816
rect 109940 546758 111859 546760
rect 111793 546755 111859 546758
rect 251173 546682 251239 546685
rect 251173 546680 253644 546682
rect 251173 546624 251178 546680
rect 251234 546624 253644 546680
rect 251173 546622 253644 546624
rect 251173 546619 251239 546622
rect 111885 546138 111951 546141
rect 109940 546136 111951 546138
rect 109940 546080 111890 546136
rect 111946 546080 111951 546136
rect 109940 546078 111951 546080
rect 111885 546075 111951 546078
rect 111793 545458 111859 545461
rect 109940 545456 111859 545458
rect 109940 545400 111798 545456
rect 111854 545400 111859 545456
rect 109940 545398 111859 545400
rect 111793 545395 111859 545398
rect 251173 545458 251239 545461
rect 251173 545456 253644 545458
rect 251173 545400 251178 545456
rect 251234 545400 253644 545456
rect 251173 545398 253644 545400
rect 251173 545395 251239 545398
rect 112897 544778 112963 544781
rect 109940 544776 112963 544778
rect 109940 544720 112902 544776
rect 112958 544720 112963 544776
rect 109940 544718 112963 544720
rect 112897 544715 112963 544718
rect 251173 544234 251239 544237
rect 251173 544232 253644 544234
rect 251173 544176 251178 544232
rect 251234 544176 253644 544232
rect 251173 544174 253644 544176
rect 251173 544171 251239 544174
rect 111793 544098 111859 544101
rect 109940 544096 111859 544098
rect 109940 544040 111798 544096
rect 111854 544040 111859 544096
rect 109940 544038 111859 544040
rect 111793 544035 111859 544038
rect 111885 543418 111951 543421
rect 109940 543416 111951 543418
rect 109940 543360 111890 543416
rect 111946 543360 111951 543416
rect 109940 543358 111951 543360
rect 111885 543355 111951 543358
rect 250713 543010 250779 543013
rect 250713 543008 253644 543010
rect 250713 542952 250718 543008
rect 250774 542952 253644 543008
rect 250713 542950 253644 542952
rect 250713 542947 250779 542950
rect 111793 542738 111859 542741
rect 109940 542736 111859 542738
rect 109940 542680 111798 542736
rect 111854 542680 111859 542736
rect 109940 542678 111859 542680
rect 111793 542675 111859 542678
rect 111793 542058 111859 542061
rect 109940 542056 111859 542058
rect 109940 542000 111798 542056
rect 111854 542000 111859 542056
rect 109940 541998 111859 542000
rect 111793 541995 111859 541998
rect 251173 541786 251239 541789
rect 251173 541784 253644 541786
rect 251173 541728 251178 541784
rect 251234 541728 253644 541784
rect 251173 541726 253644 541728
rect 251173 541723 251239 541726
rect 113081 541378 113147 541381
rect 109940 541376 113147 541378
rect 109940 541320 113086 541376
rect 113142 541320 113147 541376
rect 109940 541318 113147 541320
rect 113081 541315 113147 541318
rect -960 540684 480 540924
rect 112345 540698 112411 540701
rect 109940 540696 112411 540698
rect 109940 540640 112350 540696
rect 112406 540640 112411 540696
rect 109940 540638 112411 540640
rect 112345 540635 112411 540638
rect 251173 540562 251239 540565
rect 251173 540560 253644 540562
rect 251173 540504 251178 540560
rect 251234 540504 253644 540560
rect 251173 540502 253644 540504
rect 251173 540499 251239 540502
rect 111793 540018 111859 540021
rect 109940 540016 111859 540018
rect 109940 539960 111798 540016
rect 111854 539960 111859 540016
rect 109940 539958 111859 539960
rect 111793 539955 111859 539958
rect 111885 539338 111951 539341
rect 109940 539336 111951 539338
rect 109940 539280 111890 539336
rect 111946 539280 111951 539336
rect 109940 539278 111951 539280
rect 111885 539275 111951 539278
rect 251173 539338 251239 539341
rect 251173 539336 253644 539338
rect 251173 539280 251178 539336
rect 251234 539280 253644 539336
rect 251173 539278 253644 539280
rect 251173 539275 251239 539278
rect 111793 538658 111859 538661
rect 109940 538656 111859 538658
rect 109940 538600 111798 538656
rect 111854 538600 111859 538656
rect 109940 538598 111859 538600
rect 111793 538595 111859 538598
rect 251173 538114 251239 538117
rect 251173 538112 253644 538114
rect 251173 538056 251178 538112
rect 251234 538056 253644 538112
rect 251173 538054 253644 538056
rect 251173 538051 251239 538054
rect 111885 537978 111951 537981
rect 109940 537976 111951 537978
rect 109940 537920 111890 537976
rect 111946 537920 111951 537976
rect 109940 537918 111951 537920
rect 111885 537915 111951 537918
rect 580165 537842 580231 537845
rect 583520 537842 584960 537932
rect 580165 537840 584960 537842
rect 580165 537784 580170 537840
rect 580226 537784 584960 537840
rect 580165 537782 584960 537784
rect 580165 537779 580231 537782
rect 583520 537692 584960 537782
rect 111793 537298 111859 537301
rect 109940 537296 111859 537298
rect 109940 537240 111798 537296
rect 111854 537240 111859 537296
rect 109940 537238 111859 537240
rect 111793 537235 111859 537238
rect 252185 536890 252251 536893
rect 252185 536888 253644 536890
rect 252185 536832 252190 536888
rect 252246 536832 253644 536888
rect 252185 536830 253644 536832
rect 252185 536827 252251 536830
rect 111885 536618 111951 536621
rect 109940 536616 111951 536618
rect 109940 536560 111890 536616
rect 111946 536560 111951 536616
rect 109940 536558 111951 536560
rect 111885 536555 111951 536558
rect 111793 535938 111859 535941
rect 109940 535936 111859 535938
rect 109940 535880 111798 535936
rect 111854 535880 111859 535936
rect 109940 535878 111859 535880
rect 111793 535875 111859 535878
rect 251173 535666 251239 535669
rect 251173 535664 253644 535666
rect 251173 535608 251178 535664
rect 251234 535608 253644 535664
rect 251173 535606 253644 535608
rect 251173 535603 251239 535606
rect 111793 535258 111859 535261
rect 109940 535256 111859 535258
rect 109940 535200 111798 535256
rect 111854 535200 111859 535256
rect 109940 535198 111859 535200
rect 111793 535195 111859 535198
rect 111885 534578 111951 534581
rect 109940 534576 111951 534578
rect 109940 534520 111890 534576
rect 111946 534520 111951 534576
rect 109940 534518 111951 534520
rect 111885 534515 111951 534518
rect 251173 534442 251239 534445
rect 251173 534440 253644 534442
rect 251173 534384 251178 534440
rect 251234 534384 253644 534440
rect 251173 534382 253644 534384
rect 251173 534379 251239 534382
rect 112713 533898 112779 533901
rect 109940 533896 112779 533898
rect 109940 533840 112718 533896
rect 112774 533840 112779 533896
rect 109940 533838 112779 533840
rect 112713 533835 112779 533838
rect 113081 533218 113147 533221
rect 109940 533216 113147 533218
rect 109940 533160 113086 533216
rect 113142 533160 113147 533216
rect 109940 533158 113147 533160
rect 113081 533155 113147 533158
rect 252001 533218 252067 533221
rect 252001 533216 253644 533218
rect 252001 533160 252006 533216
rect 252062 533160 253644 533216
rect 252001 533158 253644 533160
rect 252001 533155 252067 533158
rect 112253 532538 112319 532541
rect 109940 532536 112319 532538
rect 109940 532480 112258 532536
rect 112314 532480 112319 532536
rect 109940 532478 112319 532480
rect 112253 532475 112319 532478
rect 113081 531858 113147 531861
rect 109940 531856 113147 531858
rect 109940 531800 113086 531856
rect 113142 531800 113147 531856
rect 109940 531798 113147 531800
rect 113081 531795 113147 531798
rect 113081 531178 113147 531181
rect 109940 531176 113147 531178
rect 109940 531120 113086 531176
rect 113142 531120 113147 531176
rect 109940 531118 113147 531120
rect 113081 531115 113147 531118
rect 112621 530498 112687 530501
rect 109940 530496 112687 530498
rect 109940 530440 112626 530496
rect 112682 530440 112687 530496
rect 109940 530438 112687 530440
rect 112621 530435 112687 530438
rect 112345 529818 112411 529821
rect 109940 529816 112411 529818
rect 109940 529760 112350 529816
rect 112406 529760 112411 529816
rect 109940 529758 112411 529760
rect 112345 529755 112411 529758
rect 113081 529138 113147 529141
rect 109940 529136 113147 529138
rect 109940 529080 113086 529136
rect 113142 529080 113147 529136
rect 109940 529078 113147 529080
rect 113081 529075 113147 529078
rect 111793 528458 111859 528461
rect 109940 528456 111859 528458
rect 109940 528400 111798 528456
rect 111854 528400 111859 528456
rect 109940 528398 111859 528400
rect 111793 528395 111859 528398
rect -960 527914 480 528004
rect 2957 527914 3023 527917
rect -960 527912 3023 527914
rect -960 527856 2962 527912
rect 3018 527856 3023 527912
rect -960 527854 3023 527856
rect -960 527764 480 527854
rect 2957 527851 3023 527854
rect 112253 527778 112319 527781
rect 109940 527776 112319 527778
rect 109940 527720 112258 527776
rect 112314 527720 112319 527776
rect 109940 527718 112319 527720
rect 112253 527715 112319 527718
rect 112345 527098 112411 527101
rect 109940 527096 112411 527098
rect 109940 527040 112350 527096
rect 112406 527040 112411 527096
rect 109940 527038 112411 527040
rect 112345 527035 112411 527038
rect 113081 526418 113147 526421
rect 109940 526416 113147 526418
rect 109940 526360 113086 526416
rect 113142 526360 113147 526416
rect 109940 526358 113147 526360
rect 113081 526355 113147 526358
rect 112069 525738 112135 525741
rect 109940 525736 112135 525738
rect 109940 525680 112074 525736
rect 112130 525680 112135 525736
rect 109940 525678 112135 525680
rect 112069 525675 112135 525678
rect 112713 525058 112779 525061
rect 109940 525056 112779 525058
rect 109940 525000 112718 525056
rect 112774 525000 112779 525056
rect 109940 524998 112779 525000
rect 112713 524995 112779 524998
rect 580165 524514 580231 524517
rect 583520 524514 584960 524604
rect 580165 524512 584960 524514
rect 580165 524456 580170 524512
rect 580226 524456 584960 524512
rect 580165 524454 584960 524456
rect 580165 524451 580231 524454
rect 111885 524378 111951 524381
rect 109940 524376 111951 524378
rect 109940 524320 111890 524376
rect 111946 524320 111951 524376
rect 583520 524364 584960 524454
rect 109940 524318 111951 524320
rect 111885 524315 111951 524318
rect 111793 523698 111859 523701
rect 109940 523696 111859 523698
rect 109940 523640 111798 523696
rect 111854 523640 111859 523696
rect 109940 523638 111859 523640
rect 111793 523635 111859 523638
rect 111885 523018 111951 523021
rect 109940 523016 111951 523018
rect 109940 522960 111890 523016
rect 111946 522960 111951 523016
rect 109940 522958 111951 522960
rect 111885 522955 111951 522958
rect 111793 522338 111859 522341
rect 109940 522336 111859 522338
rect 109940 522280 111798 522336
rect 111854 522280 111859 522336
rect 109940 522278 111859 522280
rect 111793 522275 111859 522278
rect 111885 521658 111951 521661
rect 109940 521656 111951 521658
rect 109940 521600 111890 521656
rect 111946 521600 111951 521656
rect 109940 521598 111951 521600
rect 111885 521595 111951 521598
rect 111793 520978 111859 520981
rect 109940 520976 111859 520978
rect 109940 520920 111798 520976
rect 111854 520920 111859 520976
rect 109940 520918 111859 520920
rect 111793 520915 111859 520918
rect 111793 520298 111859 520301
rect 109940 520296 111859 520298
rect 109940 520240 111798 520296
rect 111854 520240 111859 520296
rect 109940 520238 111859 520240
rect 111793 520235 111859 520238
rect 112345 519618 112411 519621
rect 109940 519616 112411 519618
rect 109940 519560 112350 519616
rect 112406 519560 112411 519616
rect 109940 519558 112411 519560
rect 112345 519555 112411 519558
rect 112253 518938 112319 518941
rect 109940 518936 112319 518938
rect 109940 518880 112258 518936
rect 112314 518880 112319 518936
rect 109940 518878 112319 518880
rect 112253 518875 112319 518878
rect 112805 518258 112871 518261
rect 109940 518256 112871 518258
rect 109940 518200 112810 518256
rect 112866 518200 112871 518256
rect 109940 518198 112871 518200
rect 112805 518195 112871 518198
rect 111793 517578 111859 517581
rect 109940 517576 111859 517578
rect 109940 517520 111798 517576
rect 111854 517520 111859 517576
rect 109940 517518 111859 517520
rect 111793 517515 111859 517518
rect 111885 516898 111951 516901
rect 109940 516896 111951 516898
rect 109940 516840 111890 516896
rect 111946 516840 111951 516896
rect 109940 516838 111951 516840
rect 111885 516835 111951 516838
rect 111793 516218 111859 516221
rect 109940 516216 111859 516218
rect 109940 516160 111798 516216
rect 111854 516160 111859 516216
rect 109940 516158 111859 516160
rect 111793 516155 111859 516158
rect 111885 515538 111951 515541
rect 109940 515536 111951 515538
rect 109940 515480 111890 515536
rect 111946 515480 111951 515536
rect 109940 515478 111951 515480
rect 111885 515475 111951 515478
rect -960 514858 480 514948
rect 3509 514858 3575 514861
rect 111793 514858 111859 514861
rect -960 514856 3575 514858
rect -960 514800 3514 514856
rect 3570 514800 3575 514856
rect -960 514798 3575 514800
rect 109940 514856 111859 514858
rect 109940 514800 111798 514856
rect 111854 514800 111859 514856
rect 109940 514798 111859 514800
rect -960 514708 480 514798
rect 3509 514795 3575 514798
rect 111793 514795 111859 514798
rect 111885 514178 111951 514181
rect 109940 514176 111951 514178
rect 109940 514120 111890 514176
rect 111946 514120 111951 514176
rect 109940 514118 111951 514120
rect 111885 514115 111951 514118
rect 111793 513498 111859 513501
rect 109940 513496 111859 513498
rect 109940 513440 111798 513496
rect 111854 513440 111859 513496
rect 109940 513438 111859 513440
rect 111793 513435 111859 513438
rect 111977 512818 112043 512821
rect 109940 512816 112043 512818
rect 109940 512760 111982 512816
rect 112038 512760 112043 512816
rect 109940 512758 112043 512760
rect 111977 512755 112043 512758
rect 111793 512138 111859 512141
rect 109940 512136 111859 512138
rect 109940 512080 111798 512136
rect 111854 512080 111859 512136
rect 109940 512078 111859 512080
rect 111793 512075 111859 512078
rect 111885 511458 111951 511461
rect 109940 511456 111951 511458
rect 109940 511400 111890 511456
rect 111946 511400 111951 511456
rect 109940 511398 111951 511400
rect 111885 511395 111951 511398
rect 580165 511322 580231 511325
rect 583520 511322 584960 511412
rect 580165 511320 584960 511322
rect 580165 511264 580170 511320
rect 580226 511264 584960 511320
rect 580165 511262 584960 511264
rect 580165 511259 580231 511262
rect 583520 511172 584960 511262
rect 111793 510778 111859 510781
rect 109940 510776 111859 510778
rect 109940 510720 111798 510776
rect 111854 510720 111859 510776
rect 109940 510718 111859 510720
rect 111793 510715 111859 510718
rect 112897 510098 112963 510101
rect 109940 510096 112963 510098
rect 109940 510040 112902 510096
rect 112958 510040 112963 510096
rect 109940 510038 112963 510040
rect 112897 510035 112963 510038
rect 111793 509418 111859 509421
rect 109940 509416 111859 509418
rect 109940 509360 111798 509416
rect 111854 509360 111859 509416
rect 109940 509358 111859 509360
rect 111793 509355 111859 509358
rect 111885 508738 111951 508741
rect 109940 508736 111951 508738
rect 109940 508680 111890 508736
rect 111946 508680 111951 508736
rect 109940 508678 111951 508680
rect 111885 508675 111951 508678
rect 111793 508058 111859 508061
rect 109940 508056 111859 508058
rect 109940 508000 111798 508056
rect 111854 508000 111859 508056
rect 109940 507998 111859 508000
rect 111793 507995 111859 507998
rect 111793 507378 111859 507381
rect 109940 507376 111859 507378
rect 109940 507320 111798 507376
rect 111854 507320 111859 507376
rect 109940 507318 111859 507320
rect 111793 507315 111859 507318
rect 111885 506698 111951 506701
rect 109940 506696 111951 506698
rect 109940 506640 111890 506696
rect 111946 506640 111951 506696
rect 109940 506638 111951 506640
rect 111885 506635 111951 506638
rect 111793 506018 111859 506021
rect 109940 506016 111859 506018
rect 109940 505960 111798 506016
rect 111854 505960 111859 506016
rect 109940 505958 111859 505960
rect 111793 505955 111859 505958
rect 112345 505338 112411 505341
rect 109940 505336 112411 505338
rect 109940 505280 112350 505336
rect 112406 505280 112411 505336
rect 109940 505278 112411 505280
rect 112345 505275 112411 505278
rect 111885 504658 111951 504661
rect 109940 504656 111951 504658
rect 109940 504600 111890 504656
rect 111946 504600 111951 504656
rect 109940 504598 111951 504600
rect 111885 504595 111951 504598
rect 111793 503978 111859 503981
rect 109940 503976 111859 503978
rect 109940 503920 111798 503976
rect 111854 503920 111859 503976
rect 109940 503918 111859 503920
rect 111793 503915 111859 503918
rect 111885 503298 111951 503301
rect 109940 503296 111951 503298
rect 109940 503240 111890 503296
rect 111946 503240 111951 503296
rect 109940 503238 111951 503240
rect 111885 503235 111951 503238
rect 111793 502618 111859 502621
rect 109940 502616 111859 502618
rect 109940 502560 111798 502616
rect 111854 502560 111859 502616
rect 109940 502558 111859 502560
rect 111793 502555 111859 502558
rect 111793 501938 111859 501941
rect 109940 501936 111859 501938
rect -960 501802 480 501892
rect 109940 501880 111798 501936
rect 111854 501880 111859 501936
rect 109940 501878 111859 501880
rect 111793 501875 111859 501878
rect 3509 501802 3575 501805
rect -960 501800 3575 501802
rect -960 501744 3514 501800
rect 3570 501744 3575 501800
rect -960 501742 3575 501744
rect -960 501652 480 501742
rect 3509 501739 3575 501742
rect 111885 501258 111951 501261
rect 109940 501256 111951 501258
rect 109940 501200 111890 501256
rect 111946 501200 111951 501256
rect 109940 501198 111951 501200
rect 111885 501195 111951 501198
rect 111977 500578 112043 500581
rect 109940 500576 112043 500578
rect 109940 500520 111982 500576
rect 112038 500520 112043 500576
rect 109940 500518 112043 500520
rect 111977 500515 112043 500518
rect 111793 499898 111859 499901
rect 109940 499896 111859 499898
rect 109940 499840 111798 499896
rect 111854 499840 111859 499896
rect 109940 499838 111859 499840
rect 111793 499835 111859 499838
rect 111977 499218 112043 499221
rect 109940 499216 112043 499218
rect 109940 499160 111982 499216
rect 112038 499160 112043 499216
rect 109940 499158 112043 499160
rect 111977 499155 112043 499158
rect 111793 498538 111859 498541
rect 109940 498536 111859 498538
rect 109940 498480 111798 498536
rect 111854 498480 111859 498536
rect 109940 498478 111859 498480
rect 111793 498475 111859 498478
rect 111885 497858 111951 497861
rect 109940 497856 111951 497858
rect 109940 497800 111890 497856
rect 111946 497800 111951 497856
rect 583520 497844 584960 498084
rect 109940 497798 111951 497800
rect 111885 497795 111951 497798
rect 111793 497178 111859 497181
rect 109940 497176 111859 497178
rect 109940 497120 111798 497176
rect 111854 497120 111859 497176
rect 109940 497118 111859 497120
rect 111793 497115 111859 497118
rect 111885 496498 111951 496501
rect 109940 496496 111951 496498
rect 109940 496440 111890 496496
rect 111946 496440 111951 496496
rect 109940 496438 111951 496440
rect 111885 496435 111951 496438
rect 251173 496226 251239 496229
rect 251173 496224 253644 496226
rect 251173 496168 251178 496224
rect 251234 496168 253644 496224
rect 251173 496166 253644 496168
rect 251173 496163 251239 496166
rect 111793 495818 111859 495821
rect 109940 495816 111859 495818
rect 109940 495760 111798 495816
rect 111854 495760 111859 495816
rect 109940 495758 111859 495760
rect 111793 495755 111859 495758
rect 111793 495138 111859 495141
rect 109940 495136 111859 495138
rect 109940 495080 111798 495136
rect 111854 495080 111859 495136
rect 109940 495078 111859 495080
rect 111793 495075 111859 495078
rect 251173 495002 251239 495005
rect 251173 495000 253644 495002
rect 251173 494944 251178 495000
rect 251234 494944 253644 495000
rect 251173 494942 253644 494944
rect 251173 494939 251239 494942
rect 111793 494458 111859 494461
rect 109940 494456 111859 494458
rect 109940 494400 111798 494456
rect 111854 494400 111859 494456
rect 109940 494398 111859 494400
rect 111793 494395 111859 494398
rect 111793 493778 111859 493781
rect 109940 493776 111859 493778
rect 109940 493720 111798 493776
rect 111854 493720 111859 493776
rect 109940 493718 111859 493720
rect 111793 493715 111859 493718
rect 251173 493778 251239 493781
rect 251173 493776 253644 493778
rect 251173 493720 251178 493776
rect 251234 493720 253644 493776
rect 251173 493718 253644 493720
rect 251173 493715 251239 493718
rect 113081 493098 113147 493101
rect 109940 493096 113147 493098
rect 109940 493040 113086 493096
rect 113142 493040 113147 493096
rect 109940 493038 113147 493040
rect 113081 493035 113147 493038
rect 251173 492554 251239 492557
rect 251173 492552 253644 492554
rect 251173 492496 251178 492552
rect 251234 492496 253644 492552
rect 251173 492494 253644 492496
rect 251173 492491 251239 492494
rect 111885 492418 111951 492421
rect 109940 492416 111951 492418
rect 109940 492360 111890 492416
rect 111946 492360 111951 492416
rect 109940 492358 111951 492360
rect 111885 492355 111951 492358
rect 111793 491738 111859 491741
rect 109940 491736 111859 491738
rect 109940 491680 111798 491736
rect 111854 491680 111859 491736
rect 109940 491678 111859 491680
rect 111793 491675 111859 491678
rect 250805 491330 250871 491333
rect 250805 491328 253644 491330
rect 250805 491272 250810 491328
rect 250866 491272 253644 491328
rect 250805 491270 253644 491272
rect 250805 491267 250871 491270
rect 111885 491058 111951 491061
rect 109940 491056 111951 491058
rect 109940 491000 111890 491056
rect 111946 491000 111951 491056
rect 109940 490998 111951 491000
rect 111885 490995 111951 490998
rect 111793 490378 111859 490381
rect 109940 490376 111859 490378
rect 109940 490320 111798 490376
rect 111854 490320 111859 490376
rect 109940 490318 111859 490320
rect 111793 490315 111859 490318
rect 251173 490106 251239 490109
rect 251173 490104 253644 490106
rect 251173 490048 251178 490104
rect 251234 490048 253644 490104
rect 251173 490046 253644 490048
rect 251173 490043 251239 490046
rect 111885 489698 111951 489701
rect 109940 489696 111951 489698
rect 109940 489640 111890 489696
rect 111946 489640 111951 489696
rect 109940 489638 111951 489640
rect 111885 489635 111951 489638
rect 111793 489018 111859 489021
rect 109940 489016 111859 489018
rect 109940 488960 111798 489016
rect 111854 488960 111859 489016
rect 109940 488958 111859 488960
rect 111793 488955 111859 488958
rect 251173 488882 251239 488885
rect 251173 488880 253644 488882
rect -960 488596 480 488836
rect 251173 488824 251178 488880
rect 251234 488824 253644 488880
rect 251173 488822 253644 488824
rect 251173 488819 251239 488822
rect 111885 488338 111951 488341
rect 109940 488336 111951 488338
rect 109940 488280 111890 488336
rect 111946 488280 111951 488336
rect 109940 488278 111951 488280
rect 111885 488275 111951 488278
rect 111793 487658 111859 487661
rect 109940 487656 111859 487658
rect 109940 487600 111798 487656
rect 111854 487600 111859 487656
rect 109940 487598 111859 487600
rect 111793 487595 111859 487598
rect 251173 487658 251239 487661
rect 251173 487656 253644 487658
rect 251173 487600 251178 487656
rect 251234 487600 253644 487656
rect 251173 487598 253644 487600
rect 251173 487595 251239 487598
rect 111885 486978 111951 486981
rect 109940 486976 111951 486978
rect 109940 486920 111890 486976
rect 111946 486920 111951 486976
rect 109940 486918 111951 486920
rect 111885 486915 111951 486918
rect 251173 486434 251239 486437
rect 251173 486432 253644 486434
rect 251173 486376 251178 486432
rect 251234 486376 253644 486432
rect 251173 486374 253644 486376
rect 251173 486371 251239 486374
rect 111793 486298 111859 486301
rect 109940 486296 111859 486298
rect 109940 486240 111798 486296
rect 111854 486240 111859 486296
rect 109940 486238 111859 486240
rect 111793 486235 111859 486238
rect 112989 485618 113055 485621
rect 109940 485616 113055 485618
rect 109940 485560 112994 485616
rect 113050 485560 113055 485616
rect 109940 485558 113055 485560
rect 112989 485555 113055 485558
rect 251173 485210 251239 485213
rect 251173 485208 253644 485210
rect 251173 485152 251178 485208
rect 251234 485152 253644 485208
rect 251173 485150 253644 485152
rect 251173 485147 251239 485150
rect 111793 484938 111859 484941
rect 109940 484936 111859 484938
rect 109940 484880 111798 484936
rect 111854 484880 111859 484936
rect 109940 484878 111859 484880
rect 111793 484875 111859 484878
rect 580533 484666 580599 484669
rect 583520 484666 584960 484756
rect 580533 484664 584960 484666
rect 580533 484608 580538 484664
rect 580594 484608 584960 484664
rect 580533 484606 584960 484608
rect 580533 484603 580599 484606
rect 583520 484516 584960 484606
rect 111885 484258 111951 484261
rect 109940 484256 111951 484258
rect 109940 484200 111890 484256
rect 111946 484200 111951 484256
rect 109940 484198 111951 484200
rect 111885 484195 111951 484198
rect 251173 483986 251239 483989
rect 251173 483984 253644 483986
rect 251173 483928 251178 483984
rect 251234 483928 253644 483984
rect 251173 483926 253644 483928
rect 251173 483923 251239 483926
rect 111793 483578 111859 483581
rect 109940 483576 111859 483578
rect 109940 483520 111798 483576
rect 111854 483520 111859 483576
rect 109940 483518 111859 483520
rect 111793 483515 111859 483518
rect 111885 482898 111951 482901
rect 109940 482896 111951 482898
rect 109940 482840 111890 482896
rect 111946 482840 111951 482896
rect 109940 482838 111951 482840
rect 111885 482835 111951 482838
rect 251173 482762 251239 482765
rect 251173 482760 253644 482762
rect 251173 482704 251178 482760
rect 251234 482704 253644 482760
rect 251173 482702 253644 482704
rect 251173 482699 251239 482702
rect 111793 482218 111859 482221
rect 109940 482216 111859 482218
rect 109940 482160 111798 482216
rect 111854 482160 111859 482216
rect 109940 482158 111859 482160
rect 111793 482155 111859 482158
rect 111885 481538 111951 481541
rect 109940 481536 111951 481538
rect 109940 481480 111890 481536
rect 111946 481480 111951 481536
rect 109940 481478 111951 481480
rect 111885 481475 111951 481478
rect 251173 481538 251239 481541
rect 251173 481536 253644 481538
rect 251173 481480 251178 481536
rect 251234 481480 253644 481536
rect 251173 481478 253644 481480
rect 251173 481475 251239 481478
rect 111793 480858 111859 480861
rect 109940 480856 111859 480858
rect 109940 480800 111798 480856
rect 111854 480800 111859 480856
rect 109940 480798 111859 480800
rect 111793 480795 111859 480798
rect 252369 480314 252435 480317
rect 252369 480312 253644 480314
rect 252369 480256 252374 480312
rect 252430 480256 253644 480312
rect 252369 480254 253644 480256
rect 252369 480251 252435 480254
rect 111885 480178 111951 480181
rect 109940 480176 111951 480178
rect 109940 480120 111890 480176
rect 111946 480120 111951 480176
rect 109940 480118 111951 480120
rect 111885 480115 111951 480118
rect 111793 479498 111859 479501
rect 109940 479496 111859 479498
rect 109940 479440 111798 479496
rect 111854 479440 111859 479496
rect 109940 479438 111859 479440
rect 111793 479435 111859 479438
rect 251173 479090 251239 479093
rect 251173 479088 253644 479090
rect 251173 479032 251178 479088
rect 251234 479032 253644 479088
rect 251173 479030 253644 479032
rect 251173 479027 251239 479030
rect 111885 478818 111951 478821
rect 109940 478816 111951 478818
rect 109940 478760 111890 478816
rect 111946 478760 111951 478816
rect 109940 478758 111951 478760
rect 111885 478755 111951 478758
rect 111793 478138 111859 478141
rect 109940 478136 111859 478138
rect 109940 478080 111798 478136
rect 111854 478080 111859 478136
rect 109940 478078 111859 478080
rect 111793 478075 111859 478078
rect 251173 477866 251239 477869
rect 251173 477864 253644 477866
rect 251173 477808 251178 477864
rect 251234 477808 253644 477864
rect 251173 477806 253644 477808
rect 251173 477803 251239 477806
rect 113081 477458 113147 477461
rect 109940 477456 113147 477458
rect 109940 477400 113086 477456
rect 113142 477400 113147 477456
rect 109940 477398 113147 477400
rect 113081 477395 113147 477398
rect 111793 476778 111859 476781
rect 109940 476776 111859 476778
rect 109940 476720 111798 476776
rect 111854 476720 111859 476776
rect 109940 476718 111859 476720
rect 111793 476715 111859 476718
rect 251173 476642 251239 476645
rect 251173 476640 253644 476642
rect 251173 476584 251178 476640
rect 251234 476584 253644 476640
rect 251173 476582 253644 476584
rect 251173 476579 251239 476582
rect 111885 476098 111951 476101
rect 109940 476096 111951 476098
rect 109940 476040 111890 476096
rect 111946 476040 111951 476096
rect 109940 476038 111951 476040
rect 111885 476035 111951 476038
rect -960 475690 480 475780
rect 3601 475690 3667 475693
rect -960 475688 3667 475690
rect -960 475632 3606 475688
rect 3662 475632 3667 475688
rect -960 475630 3667 475632
rect -960 475540 480 475630
rect 3601 475627 3667 475630
rect 111793 475418 111859 475421
rect 109940 475416 111859 475418
rect 109940 475360 111798 475416
rect 111854 475360 111859 475416
rect 109940 475358 111859 475360
rect 111793 475355 111859 475358
rect 251173 475418 251239 475421
rect 251173 475416 253644 475418
rect 251173 475360 251178 475416
rect 251234 475360 253644 475416
rect 251173 475358 253644 475360
rect 251173 475355 251239 475358
rect 111793 474738 111859 474741
rect 109940 474736 111859 474738
rect 109940 474680 111798 474736
rect 111854 474680 111859 474736
rect 109940 474678 111859 474680
rect 111793 474675 111859 474678
rect 251173 474194 251239 474197
rect 251173 474192 253644 474194
rect 251173 474136 251178 474192
rect 251234 474136 253644 474192
rect 251173 474134 253644 474136
rect 251173 474131 251239 474134
rect 111885 474058 111951 474061
rect 109940 474056 111951 474058
rect 109940 474000 111890 474056
rect 111946 474000 111951 474056
rect 109940 473998 111951 474000
rect 111885 473995 111951 473998
rect 111793 473378 111859 473381
rect 109940 473376 111859 473378
rect 109940 473320 111798 473376
rect 111854 473320 111859 473376
rect 109940 473318 111859 473320
rect 111793 473315 111859 473318
rect 251173 472970 251239 472973
rect 251173 472968 253644 472970
rect 251173 472912 251178 472968
rect 251234 472912 253644 472968
rect 251173 472910 253644 472912
rect 251173 472907 251239 472910
rect 111885 472698 111951 472701
rect 109940 472696 111951 472698
rect 109940 472640 111890 472696
rect 111946 472640 111951 472696
rect 109940 472638 111951 472640
rect 111885 472635 111951 472638
rect 111793 472018 111859 472021
rect 109940 472016 111859 472018
rect 109940 471960 111798 472016
rect 111854 471960 111859 472016
rect 109940 471958 111859 471960
rect 111793 471955 111859 471958
rect 251173 471746 251239 471749
rect 251173 471744 253644 471746
rect 251173 471688 251178 471744
rect 251234 471688 253644 471744
rect 251173 471686 253644 471688
rect 251173 471683 251239 471686
rect 580625 471474 580691 471477
rect 583520 471474 584960 471564
rect 580625 471472 584960 471474
rect 580625 471416 580630 471472
rect 580686 471416 584960 471472
rect 580625 471414 584960 471416
rect 580625 471411 580691 471414
rect 111885 471338 111951 471341
rect 109940 471336 111951 471338
rect 109940 471280 111890 471336
rect 111946 471280 111951 471336
rect 583520 471324 584960 471414
rect 109940 471278 111951 471280
rect 111885 471275 111951 471278
rect 111793 470658 111859 470661
rect 109940 470656 111859 470658
rect 109940 470600 111798 470656
rect 111854 470600 111859 470656
rect 109940 470598 111859 470600
rect 111793 470595 111859 470598
rect 251265 470522 251331 470525
rect 251265 470520 253644 470522
rect 251265 470464 251270 470520
rect 251326 470464 253644 470520
rect 251265 470462 253644 470464
rect 251265 470459 251331 470462
rect 111793 469978 111859 469981
rect 109940 469976 111859 469978
rect 109940 469920 111798 469976
rect 111854 469920 111859 469976
rect 109940 469918 111859 469920
rect 111793 469915 111859 469918
rect 111793 469298 111859 469301
rect 109940 469296 111859 469298
rect 109940 469240 111798 469296
rect 111854 469240 111859 469296
rect 109940 469238 111859 469240
rect 111793 469235 111859 469238
rect 251173 469298 251239 469301
rect 251173 469296 253644 469298
rect 251173 469240 251178 469296
rect 251234 469240 253644 469296
rect 251173 469238 253644 469240
rect 251173 469235 251239 469238
rect 111885 468618 111951 468621
rect 109940 468616 111951 468618
rect 109940 468560 111890 468616
rect 111946 468560 111951 468616
rect 109940 468558 111951 468560
rect 111885 468555 111951 468558
rect 252185 468074 252251 468077
rect 252185 468072 253644 468074
rect 252185 468016 252190 468072
rect 252246 468016 253644 468072
rect 252185 468014 253644 468016
rect 252185 468011 252251 468014
rect 111793 467938 111859 467941
rect 109940 467936 111859 467938
rect 109940 467880 111798 467936
rect 111854 467880 111859 467936
rect 109940 467878 111859 467880
rect 111793 467875 111859 467878
rect 111885 467258 111951 467261
rect 109940 467256 111951 467258
rect 109940 467200 111890 467256
rect 111946 467200 111951 467256
rect 109940 467198 111951 467200
rect 111885 467195 111951 467198
rect 251173 466850 251239 466853
rect 251173 466848 253644 466850
rect 251173 466792 251178 466848
rect 251234 466792 253644 466848
rect 251173 466790 253644 466792
rect 251173 466787 251239 466790
rect 111793 466578 111859 466581
rect 109940 466576 111859 466578
rect 109940 466520 111798 466576
rect 111854 466520 111859 466576
rect 109940 466518 111859 466520
rect 111793 466515 111859 466518
rect 111885 465898 111951 465901
rect 109940 465896 111951 465898
rect 109940 465840 111890 465896
rect 111946 465840 111951 465896
rect 109940 465838 111951 465840
rect 111885 465835 111951 465838
rect 251633 465626 251699 465629
rect 251633 465624 253644 465626
rect 251633 465568 251638 465624
rect 251694 465568 253644 465624
rect 251633 465566 253644 465568
rect 251633 465563 251699 465566
rect 111793 465218 111859 465221
rect 109940 465216 111859 465218
rect 109940 465160 111798 465216
rect 111854 465160 111859 465216
rect 109940 465158 111859 465160
rect 111793 465155 111859 465158
rect 111885 464538 111951 464541
rect 109940 464536 111951 464538
rect 109940 464480 111890 464536
rect 111946 464480 111951 464536
rect 109940 464478 111951 464480
rect 111885 464475 111951 464478
rect 251173 464402 251239 464405
rect 251173 464400 253644 464402
rect 251173 464344 251178 464400
rect 251234 464344 253644 464400
rect 251173 464342 253644 464344
rect 251173 464339 251239 464342
rect 111793 463858 111859 463861
rect 109940 463856 111859 463858
rect 109940 463800 111798 463856
rect 111854 463800 111859 463856
rect 109940 463798 111859 463800
rect 111793 463795 111859 463798
rect 111885 463178 111951 463181
rect 109940 463176 111951 463178
rect 109940 463120 111890 463176
rect 111946 463120 111951 463176
rect 109940 463118 111951 463120
rect 111885 463115 111951 463118
rect 251173 463178 251239 463181
rect 251173 463176 253644 463178
rect 251173 463120 251178 463176
rect 251234 463120 253644 463176
rect 251173 463118 253644 463120
rect 251173 463115 251239 463118
rect -960 462634 480 462724
rect 3693 462634 3759 462637
rect -960 462632 3759 462634
rect -960 462576 3698 462632
rect 3754 462576 3759 462632
rect -960 462574 3759 462576
rect -960 462484 480 462574
rect 3693 462571 3759 462574
rect 111793 462498 111859 462501
rect 109940 462496 111859 462498
rect 109940 462440 111798 462496
rect 111854 462440 111859 462496
rect 109940 462438 111859 462440
rect 111793 462435 111859 462438
rect 252461 461954 252527 461957
rect 252461 461952 253644 461954
rect 252461 461896 252466 461952
rect 252522 461896 253644 461952
rect 252461 461894 253644 461896
rect 252461 461891 252527 461894
rect 111885 461818 111951 461821
rect 109940 461816 111951 461818
rect 109940 461760 111890 461816
rect 111946 461760 111951 461816
rect 109940 461758 111951 461760
rect 111885 461755 111951 461758
rect 111793 461138 111859 461141
rect 109940 461136 111859 461138
rect 109940 461080 111798 461136
rect 111854 461080 111859 461136
rect 109940 461078 111859 461080
rect 111793 461075 111859 461078
rect 251173 460730 251239 460733
rect 251173 460728 253644 460730
rect 251173 460672 251178 460728
rect 251234 460672 253644 460728
rect 251173 460670 253644 460672
rect 251173 460667 251239 460670
rect 111793 460458 111859 460461
rect 109940 460456 111859 460458
rect 109940 460400 111798 460456
rect 111854 460400 111859 460456
rect 109940 460398 111859 460400
rect 111793 460395 111859 460398
rect 112345 459778 112411 459781
rect 109940 459776 112411 459778
rect 109940 459720 112350 459776
rect 112406 459720 112411 459776
rect 109940 459718 112411 459720
rect 112345 459715 112411 459718
rect 251173 459506 251239 459509
rect 251173 459504 253644 459506
rect 251173 459448 251178 459504
rect 251234 459448 253644 459504
rect 251173 459446 253644 459448
rect 251173 459443 251239 459446
rect 111885 459098 111951 459101
rect 109940 459096 111951 459098
rect 109940 459040 111890 459096
rect 111946 459040 111951 459096
rect 109940 459038 111951 459040
rect 111885 459035 111951 459038
rect 111793 458418 111859 458421
rect 109940 458416 111859 458418
rect 109940 458360 111798 458416
rect 111854 458360 111859 458416
rect 109940 458358 111859 458360
rect 111793 458355 111859 458358
rect 252093 458282 252159 458285
rect 252093 458280 253644 458282
rect 252093 458224 252098 458280
rect 252154 458224 253644 458280
rect 252093 458222 253644 458224
rect 252093 458219 252159 458222
rect 580165 458146 580231 458149
rect 583520 458146 584960 458236
rect 580165 458144 584960 458146
rect 580165 458088 580170 458144
rect 580226 458088 584960 458144
rect 580165 458086 584960 458088
rect 580165 458083 580231 458086
rect 583520 457996 584960 458086
rect 112253 457738 112319 457741
rect 109940 457736 112319 457738
rect 109940 457680 112258 457736
rect 112314 457680 112319 457736
rect 109940 457678 112319 457680
rect 112253 457675 112319 457678
rect 111793 457058 111859 457061
rect 109940 457056 111859 457058
rect 109940 457000 111798 457056
rect 111854 457000 111859 457056
rect 109940 456998 111859 457000
rect 111793 456995 111859 456998
rect 251173 457058 251239 457061
rect 251173 457056 253644 457058
rect 251173 457000 251178 457056
rect 251234 457000 253644 457056
rect 251173 456998 253644 457000
rect 251173 456995 251239 456998
rect 111885 456378 111951 456381
rect 109940 456376 111951 456378
rect 109940 456320 111890 456376
rect 111946 456320 111951 456376
rect 109940 456318 111951 456320
rect 111885 456315 111951 456318
rect 251173 455834 251239 455837
rect 251173 455832 253644 455834
rect 251173 455776 251178 455832
rect 251234 455776 253644 455832
rect 251173 455774 253644 455776
rect 251173 455771 251239 455774
rect 111793 455698 111859 455701
rect 109940 455696 111859 455698
rect 109940 455640 111798 455696
rect 111854 455640 111859 455696
rect 109940 455638 111859 455640
rect 111793 455635 111859 455638
rect 111793 455018 111859 455021
rect 109940 455016 111859 455018
rect 109940 454960 111798 455016
rect 111854 454960 111859 455016
rect 109940 454958 111859 454960
rect 111793 454955 111859 454958
rect 251173 454610 251239 454613
rect 251173 454608 253644 454610
rect 251173 454552 251178 454608
rect 251234 454552 253644 454608
rect 251173 454550 253644 454552
rect 251173 454547 251239 454550
rect 111793 454338 111859 454341
rect 109940 454336 111859 454338
rect 109940 454280 111798 454336
rect 111854 454280 111859 454336
rect 109940 454278 111859 454280
rect 111793 454275 111859 454278
rect 111885 453658 111951 453661
rect 109940 453656 111951 453658
rect 109940 453600 111890 453656
rect 111946 453600 111951 453656
rect 109940 453598 111951 453600
rect 111885 453595 111951 453598
rect 251725 453386 251791 453389
rect 251725 453384 253644 453386
rect 251725 453328 251730 453384
rect 251786 453328 253644 453384
rect 251725 453326 253644 453328
rect 251725 453323 251791 453326
rect 111793 452978 111859 452981
rect 109940 452976 111859 452978
rect 109940 452920 111798 452976
rect 111854 452920 111859 452976
rect 109940 452918 111859 452920
rect 111793 452915 111859 452918
rect 111885 452298 111951 452301
rect 109940 452296 111951 452298
rect 109940 452240 111890 452296
rect 111946 452240 111951 452296
rect 109940 452238 111951 452240
rect 111885 452235 111951 452238
rect 251173 452162 251239 452165
rect 251173 452160 253644 452162
rect 251173 452104 251178 452160
rect 251234 452104 253644 452160
rect 251173 452102 253644 452104
rect 251173 452099 251239 452102
rect 111793 451618 111859 451621
rect 109940 451616 111859 451618
rect 109940 451560 111798 451616
rect 111854 451560 111859 451616
rect 109940 451558 111859 451560
rect 111793 451555 111859 451558
rect 111885 450938 111951 450941
rect 109940 450936 111951 450938
rect 109940 450880 111890 450936
rect 111946 450880 111951 450936
rect 109940 450878 111951 450880
rect 111885 450875 111951 450878
rect 251173 450938 251239 450941
rect 251173 450936 253644 450938
rect 251173 450880 251178 450936
rect 251234 450880 253644 450936
rect 251173 450878 253644 450880
rect 251173 450875 251239 450878
rect 111793 450258 111859 450261
rect 109940 450256 111859 450258
rect 109940 450200 111798 450256
rect 111854 450200 111859 450256
rect 109940 450198 111859 450200
rect 111793 450195 111859 450198
rect 251173 449714 251239 449717
rect 251173 449712 253644 449714
rect -960 449578 480 449668
rect 251173 449656 251178 449712
rect 251234 449656 253644 449712
rect 251173 449654 253644 449656
rect 251173 449651 251239 449654
rect 3785 449578 3851 449581
rect 111885 449578 111951 449581
rect -960 449576 3851 449578
rect -960 449520 3790 449576
rect 3846 449520 3851 449576
rect -960 449518 3851 449520
rect 109940 449576 111951 449578
rect 109940 449520 111890 449576
rect 111946 449520 111951 449576
rect 109940 449518 111951 449520
rect -960 449428 480 449518
rect 3785 449515 3851 449518
rect 111885 449515 111951 449518
rect 111793 448898 111859 448901
rect 109940 448896 111859 448898
rect 109940 448840 111798 448896
rect 111854 448840 111859 448896
rect 109940 448838 111859 448840
rect 111793 448835 111859 448838
rect 252369 448490 252435 448493
rect 252369 448488 253644 448490
rect 252369 448432 252374 448488
rect 252430 448432 253644 448488
rect 252369 448430 253644 448432
rect 252369 448427 252435 448430
rect 111793 448218 111859 448221
rect 109940 448216 111859 448218
rect 109940 448160 111798 448216
rect 111854 448160 111859 448216
rect 109940 448158 111859 448160
rect 111793 448155 111859 448158
rect 251173 447266 251239 447269
rect 251173 447264 253644 447266
rect 251173 447208 251178 447264
rect 251234 447208 253644 447264
rect 251173 447206 253644 447208
rect 251173 447203 251239 447206
rect 251173 446042 251239 446045
rect 251173 446040 253644 446042
rect 251173 445984 251178 446040
rect 251234 445984 253644 446040
rect 251173 445982 253644 445984
rect 251173 445979 251239 445982
rect 251173 444818 251239 444821
rect 251173 444816 253644 444818
rect 251173 444760 251178 444816
rect 251234 444760 253644 444816
rect 251173 444758 253644 444760
rect 251173 444755 251239 444758
rect 583520 444668 584960 444908
rect 250897 443594 250963 443597
rect 250897 443592 253644 443594
rect 250897 443536 250902 443592
rect 250958 443536 253644 443592
rect 250897 443534 253644 443536
rect 250897 443531 250963 443534
rect 251173 442370 251239 442373
rect 251173 442368 253644 442370
rect 251173 442312 251178 442368
rect 251234 442312 253644 442368
rect 251173 442310 253644 442312
rect 251173 442307 251239 442310
rect 251173 441146 251239 441149
rect 251173 441144 253644 441146
rect 251173 441088 251178 441144
rect 251234 441088 253644 441144
rect 251173 441086 253644 441088
rect 251173 441083 251239 441086
rect 251173 439922 251239 439925
rect 251173 439920 253644 439922
rect 251173 439864 251178 439920
rect 251234 439864 253644 439920
rect 251173 439862 253644 439864
rect 251173 439859 251239 439862
rect 251173 438698 251239 438701
rect 251173 438696 253644 438698
rect 251173 438640 251178 438696
rect 251234 438640 253644 438696
rect 251173 438638 253644 438640
rect 251173 438635 251239 438638
rect 251265 437474 251331 437477
rect 251265 437472 253644 437474
rect 251265 437416 251270 437472
rect 251326 437416 253644 437472
rect 251265 437414 253644 437416
rect 251265 437411 251331 437414
rect -960 436508 480 436748
rect 251173 436250 251239 436253
rect 251173 436248 253644 436250
rect 251173 436192 251178 436248
rect 251234 436192 253644 436248
rect 251173 436190 253644 436192
rect 251173 436187 251239 436190
rect 251173 435026 251239 435029
rect 251173 435024 253644 435026
rect 251173 434968 251178 435024
rect 251234 434968 253644 435024
rect 251173 434966 253644 434968
rect 251173 434963 251239 434966
rect 251173 433802 251239 433805
rect 251173 433800 253644 433802
rect 251173 433744 251178 433800
rect 251234 433744 253644 433800
rect 251173 433742 253644 433744
rect 251173 433739 251239 433742
rect 251173 432578 251239 432581
rect 251173 432576 253644 432578
rect 251173 432520 251178 432576
rect 251234 432520 253644 432576
rect 251173 432518 253644 432520
rect 251173 432515 251239 432518
rect 580717 431626 580783 431629
rect 583520 431626 584960 431716
rect 580717 431624 584960 431626
rect 580717 431568 580722 431624
rect 580778 431568 584960 431624
rect 580717 431566 584960 431568
rect 580717 431563 580783 431566
rect 583520 431476 584960 431566
rect 251173 431354 251239 431357
rect 251173 431352 253644 431354
rect 251173 431296 251178 431352
rect 251234 431296 253644 431352
rect 251173 431294 253644 431296
rect 251173 431291 251239 431294
rect 251173 430130 251239 430133
rect 251173 430128 253644 430130
rect 251173 430072 251178 430128
rect 251234 430072 253644 430128
rect 251173 430070 253644 430072
rect 251173 430067 251239 430070
rect 251173 428906 251239 428909
rect 251173 428904 253644 428906
rect 251173 428848 251178 428904
rect 251234 428848 253644 428904
rect 251173 428846 253644 428848
rect 251173 428843 251239 428846
rect 251265 427682 251331 427685
rect 251265 427680 253644 427682
rect 251265 427624 251270 427680
rect 251326 427624 253644 427680
rect 251265 427622 253644 427624
rect 251265 427619 251331 427622
rect 251173 426458 251239 426461
rect 251173 426456 253644 426458
rect 251173 426400 251178 426456
rect 251234 426400 253644 426456
rect 251173 426398 253644 426400
rect 251173 426395 251239 426398
rect 251173 425234 251239 425237
rect 251173 425232 253644 425234
rect 251173 425176 251178 425232
rect 251234 425176 253644 425232
rect 251173 425174 253644 425176
rect 251173 425171 251239 425174
rect 251173 424010 251239 424013
rect 251173 424008 253644 424010
rect 251173 423952 251178 424008
rect 251234 423952 253644 424008
rect 251173 423950 253644 423952
rect 251173 423947 251239 423950
rect -960 423602 480 423692
rect 3325 423602 3391 423605
rect -960 423600 3391 423602
rect -960 423544 3330 423600
rect 3386 423544 3391 423600
rect -960 423542 3391 423544
rect -960 423452 480 423542
rect 3325 423539 3391 423542
rect 250989 422786 251055 422789
rect 250989 422784 253644 422786
rect 250989 422728 250994 422784
rect 251050 422728 253644 422784
rect 250989 422726 253644 422728
rect 250989 422723 251055 422726
rect 251173 421562 251239 421565
rect 251173 421560 253644 421562
rect 251173 421504 251178 421560
rect 251234 421504 253644 421560
rect 251173 421502 253644 421504
rect 251173 421499 251239 421502
rect 251173 420338 251239 420341
rect 251173 420336 253644 420338
rect 251173 420280 251178 420336
rect 251234 420280 253644 420336
rect 251173 420278 253644 420280
rect 251173 420275 251239 420278
rect 251173 419114 251239 419117
rect 251173 419112 253644 419114
rect 251173 419056 251178 419112
rect 251234 419056 253644 419112
rect 251173 419054 253644 419056
rect 251173 419051 251239 419054
rect 580809 418298 580875 418301
rect 583520 418298 584960 418388
rect 580809 418296 584960 418298
rect 580809 418240 580814 418296
rect 580870 418240 584960 418296
rect 580809 418238 584960 418240
rect 580809 418235 580875 418238
rect 583520 418148 584960 418238
rect 251173 417890 251239 417893
rect 251173 417888 253644 417890
rect 251173 417832 251178 417888
rect 251234 417832 253644 417888
rect 251173 417830 253644 417832
rect 251173 417827 251239 417830
rect 251265 416666 251331 416669
rect 251265 416664 253644 416666
rect 251265 416608 251270 416664
rect 251326 416608 253644 416664
rect 251265 416606 253644 416608
rect 251265 416603 251331 416606
rect 251173 415442 251239 415445
rect 251173 415440 253644 415442
rect 251173 415384 251178 415440
rect 251234 415384 253644 415440
rect 251173 415382 253644 415384
rect 251173 415379 251239 415382
rect 251173 414218 251239 414221
rect 251173 414216 253644 414218
rect 251173 414160 251178 414216
rect 251234 414160 253644 414216
rect 251173 414158 253644 414160
rect 251173 414155 251239 414158
rect 220721 413946 220787 413949
rect 217948 413944 220787 413946
rect 217948 413888 220726 413944
rect 220782 413888 220787 413944
rect 217948 413886 220787 413888
rect 220721 413883 220787 413886
rect 219985 413538 220051 413541
rect 217948 413536 220051 413538
rect 217948 413480 219990 413536
rect 220046 413480 220051 413536
rect 217948 413478 220051 413480
rect 219985 413475 220051 413478
rect 219709 413130 219775 413133
rect 217948 413128 219775 413130
rect 217948 413072 219714 413128
rect 219770 413072 219775 413128
rect 217948 413070 219775 413072
rect 219709 413067 219775 413070
rect 251173 412994 251239 412997
rect 251173 412992 253644 412994
rect 251173 412936 251178 412992
rect 251234 412936 253644 412992
rect 251173 412934 253644 412936
rect 251173 412931 251239 412934
rect 219801 412722 219867 412725
rect 217948 412720 219867 412722
rect 217948 412664 219806 412720
rect 219862 412664 219867 412720
rect 217948 412662 219867 412664
rect 219801 412659 219867 412662
rect 220721 412314 220787 412317
rect 217948 412312 220787 412314
rect 217948 412256 220726 412312
rect 220782 412256 220787 412312
rect 217948 412254 220787 412256
rect 220721 412251 220787 412254
rect 220077 411906 220143 411909
rect 217948 411904 220143 411906
rect 217948 411848 220082 411904
rect 220138 411848 220143 411904
rect 217948 411846 220143 411848
rect 220077 411843 220143 411846
rect 251173 411770 251239 411773
rect 251173 411768 253644 411770
rect 251173 411712 251178 411768
rect 251234 411712 253644 411768
rect 251173 411710 253644 411712
rect 251173 411707 251239 411710
rect 219893 411498 219959 411501
rect 217948 411496 219959 411498
rect 217948 411440 219898 411496
rect 219954 411440 219959 411496
rect 217948 411438 219959 411440
rect 219893 411435 219959 411438
rect 220721 411090 220787 411093
rect 217948 411088 220787 411090
rect 217948 411032 220726 411088
rect 220782 411032 220787 411088
rect 217948 411030 220787 411032
rect 220721 411027 220787 411030
rect 219801 410682 219867 410685
rect 217948 410680 219867 410682
rect -960 410546 480 410636
rect 217948 410624 219806 410680
rect 219862 410624 219867 410680
rect 217948 410622 219867 410624
rect 219801 410619 219867 410622
rect 3325 410546 3391 410549
rect -960 410544 3391 410546
rect -960 410488 3330 410544
rect 3386 410488 3391 410544
rect -960 410486 3391 410488
rect -960 410396 480 410486
rect 3325 410483 3391 410486
rect 251173 410546 251239 410549
rect 251173 410544 253644 410546
rect 251173 410488 251178 410544
rect 251234 410488 253644 410544
rect 251173 410486 253644 410488
rect 251173 410483 251239 410486
rect 220077 410274 220143 410277
rect 217948 410272 220143 410274
rect 217948 410216 220082 410272
rect 220138 410216 220143 410272
rect 217948 410214 220143 410216
rect 220077 410211 220143 410214
rect 220721 409866 220787 409869
rect 217948 409864 220787 409866
rect 217948 409808 220726 409864
rect 220782 409808 220787 409864
rect 217948 409806 220787 409808
rect 220721 409803 220787 409806
rect 219985 409458 220051 409461
rect 217948 409456 220051 409458
rect 217948 409400 219990 409456
rect 220046 409400 220051 409456
rect 217948 409398 220051 409400
rect 219985 409395 220051 409398
rect 251173 409322 251239 409325
rect 251173 409320 253644 409322
rect 251173 409264 251178 409320
rect 251234 409264 253644 409320
rect 251173 409262 253644 409264
rect 251173 409259 251239 409262
rect 220077 409050 220143 409053
rect 217948 409048 220143 409050
rect 217948 408992 220082 409048
rect 220138 408992 220143 409048
rect 217948 408990 220143 408992
rect 220077 408987 220143 408990
rect 219893 408642 219959 408645
rect 217948 408640 219959 408642
rect 217948 408584 219898 408640
rect 219954 408584 219959 408640
rect 217948 408582 219959 408584
rect 219893 408579 219959 408582
rect 220721 408234 220787 408237
rect 217948 408232 220787 408234
rect 217948 408176 220726 408232
rect 220782 408176 220787 408232
rect 217948 408174 220787 408176
rect 220721 408171 220787 408174
rect 251173 408098 251239 408101
rect 251173 408096 253644 408098
rect 251173 408040 251178 408096
rect 251234 408040 253644 408096
rect 251173 408038 253644 408040
rect 251173 408035 251239 408038
rect 219893 407826 219959 407829
rect 217948 407824 219959 407826
rect 217948 407768 219898 407824
rect 219954 407768 219959 407824
rect 217948 407766 219959 407768
rect 219893 407763 219959 407766
rect 154941 407418 155007 407421
rect 220077 407418 220143 407421
rect 154941 407416 158148 407418
rect 154941 407360 154946 407416
rect 155002 407360 158148 407416
rect 154941 407358 158148 407360
rect 217948 407416 220143 407418
rect 217948 407360 220082 407416
rect 220138 407360 220143 407416
rect 217948 407358 220143 407360
rect 154941 407355 155007 407358
rect 220077 407355 220143 407358
rect 155677 407146 155743 407149
rect 155677 407144 158148 407146
rect 155677 407088 155682 407144
rect 155738 407088 158148 407144
rect 155677 407086 158148 407088
rect 155677 407083 155743 407086
rect 220721 407010 220787 407013
rect 217948 407008 220787 407010
rect 217948 406952 220726 407008
rect 220782 406952 220787 407008
rect 217948 406950 220787 406952
rect 220721 406947 220787 406950
rect 154573 406874 154639 406877
rect 251633 406874 251699 406877
rect 154573 406872 158148 406874
rect 154573 406816 154578 406872
rect 154634 406816 158148 406872
rect 154573 406814 158148 406816
rect 251633 406872 253644 406874
rect 251633 406816 251638 406872
rect 251694 406816 253644 406872
rect 251633 406814 253644 406816
rect 154573 406811 154639 406814
rect 251633 406811 251699 406814
rect 154941 406602 155007 406605
rect 220721 406602 220787 406605
rect 154941 406600 158148 406602
rect 154941 406544 154946 406600
rect 155002 406544 158148 406600
rect 154941 406542 158148 406544
rect 217948 406600 220787 406602
rect 217948 406544 220726 406600
rect 220782 406544 220787 406600
rect 217948 406542 220787 406544
rect 154941 406539 155007 406542
rect 220721 406539 220787 406542
rect 154849 406330 154915 406333
rect 154849 406328 158148 406330
rect 154849 406272 154854 406328
rect 154910 406272 158148 406328
rect 154849 406270 158148 406272
rect 154849 406267 154915 406270
rect 219893 406194 219959 406197
rect 217948 406192 219959 406194
rect 217948 406136 219898 406192
rect 219954 406136 219959 406192
rect 217948 406134 219959 406136
rect 219893 406131 219959 406134
rect 154757 406058 154823 406061
rect 154757 406056 158148 406058
rect 154757 406000 154762 406056
rect 154818 406000 158148 406056
rect 154757 405998 158148 406000
rect 154757 405995 154823 405998
rect 154665 405786 154731 405789
rect 220077 405786 220143 405789
rect 154665 405784 158148 405786
rect 154665 405728 154670 405784
rect 154726 405728 158148 405784
rect 154665 405726 158148 405728
rect 217948 405784 220143 405786
rect 217948 405728 220082 405784
rect 220138 405728 220143 405784
rect 217948 405726 220143 405728
rect 154665 405723 154731 405726
rect 220077 405723 220143 405726
rect 251173 405650 251239 405653
rect 251173 405648 253644 405650
rect 251173 405592 251178 405648
rect 251234 405592 253644 405648
rect 251173 405590 253644 405592
rect 251173 405587 251239 405590
rect 154573 405514 154639 405517
rect 154573 405512 158148 405514
rect 154573 405456 154578 405512
rect 154634 405456 158148 405512
rect 154573 405454 158148 405456
rect 154573 405451 154639 405454
rect 220721 405378 220787 405381
rect 217948 405376 220787 405378
rect 217948 405320 220726 405376
rect 220782 405320 220787 405376
rect 217948 405318 220787 405320
rect 220721 405315 220787 405318
rect 154757 405242 154823 405245
rect 154757 405240 158148 405242
rect 154757 405184 154762 405240
rect 154818 405184 158148 405240
rect 154757 405182 158148 405184
rect 154757 405179 154823 405182
rect 154941 404970 155007 404973
rect 219893 404970 219959 404973
rect 154941 404968 158148 404970
rect 154941 404912 154946 404968
rect 155002 404912 158148 404968
rect 154941 404910 158148 404912
rect 217948 404968 219959 404970
rect 217948 404912 219898 404968
rect 219954 404912 219959 404968
rect 217948 404910 219959 404912
rect 154941 404907 155007 404910
rect 219893 404907 219959 404910
rect 580901 404970 580967 404973
rect 583520 404970 584960 405060
rect 580901 404968 584960 404970
rect 580901 404912 580906 404968
rect 580962 404912 584960 404968
rect 580901 404910 584960 404912
rect 580901 404907 580967 404910
rect 583520 404820 584960 404910
rect 154849 404698 154915 404701
rect 154849 404696 158148 404698
rect 154849 404640 154854 404696
rect 154910 404640 158148 404696
rect 154849 404638 158148 404640
rect 154849 404635 154915 404638
rect 220077 404562 220143 404565
rect 217948 404560 220143 404562
rect 217948 404504 220082 404560
rect 220138 404504 220143 404560
rect 217948 404502 220143 404504
rect 220077 404499 220143 404502
rect 155769 404426 155835 404429
rect 251725 404426 251791 404429
rect 155769 404424 158148 404426
rect 155769 404368 155774 404424
rect 155830 404368 158148 404424
rect 155769 404366 158148 404368
rect 251725 404424 253644 404426
rect 251725 404368 251730 404424
rect 251786 404368 253644 404424
rect 251725 404366 253644 404368
rect 155769 404363 155835 404366
rect 251725 404363 251791 404366
rect 154665 404154 154731 404157
rect 220721 404154 220787 404157
rect 154665 404152 158148 404154
rect 154665 404096 154670 404152
rect 154726 404096 158148 404152
rect 154665 404094 158148 404096
rect 217948 404152 220787 404154
rect 217948 404096 220726 404152
rect 220782 404096 220787 404152
rect 217948 404094 220787 404096
rect 154665 404091 154731 404094
rect 220721 404091 220787 404094
rect 154757 403882 154823 403885
rect 154757 403880 158148 403882
rect 154757 403824 154762 403880
rect 154818 403824 158148 403880
rect 154757 403822 158148 403824
rect 154757 403819 154823 403822
rect 220077 403746 220143 403749
rect 217948 403744 220143 403746
rect 217948 403688 220082 403744
rect 220138 403688 220143 403744
rect 217948 403686 220143 403688
rect 220077 403683 220143 403686
rect 154941 403610 155007 403613
rect 154941 403608 158148 403610
rect 154941 403552 154946 403608
rect 155002 403552 158148 403608
rect 154941 403550 158148 403552
rect 154941 403547 155007 403550
rect 154849 403338 154915 403341
rect 219985 403338 220051 403341
rect 154849 403336 158148 403338
rect 154849 403280 154854 403336
rect 154910 403280 158148 403336
rect 154849 403278 158148 403280
rect 217948 403336 220051 403338
rect 217948 403280 219990 403336
rect 220046 403280 220051 403336
rect 217948 403278 220051 403280
rect 154849 403275 154915 403278
rect 219985 403275 220051 403278
rect 251081 403202 251147 403205
rect 251081 403200 253644 403202
rect 251081 403144 251086 403200
rect 251142 403144 253644 403200
rect 251081 403142 253644 403144
rect 251081 403139 251147 403142
rect 155217 403066 155283 403069
rect 155217 403064 158148 403066
rect 155217 403008 155222 403064
rect 155278 403008 158148 403064
rect 155217 403006 158148 403008
rect 155217 403003 155283 403006
rect 219801 402930 219867 402933
rect 217948 402928 219867 402930
rect 217948 402872 219806 402928
rect 219862 402872 219867 402928
rect 217948 402870 219867 402872
rect 219801 402867 219867 402870
rect 154665 402794 154731 402797
rect 154665 402792 158148 402794
rect 154665 402736 154670 402792
rect 154726 402736 158148 402792
rect 154665 402734 158148 402736
rect 154665 402731 154731 402734
rect 154849 402522 154915 402525
rect 219709 402522 219775 402525
rect 154849 402520 158148 402522
rect 154849 402464 154854 402520
rect 154910 402464 158148 402520
rect 154849 402462 158148 402464
rect 217948 402520 219775 402522
rect 217948 402464 219714 402520
rect 219770 402464 219775 402520
rect 217948 402462 219775 402464
rect 154849 402459 154915 402462
rect 219709 402459 219775 402462
rect 154757 402250 154823 402253
rect 154757 402248 158148 402250
rect 154757 402192 154762 402248
rect 154818 402192 158148 402248
rect 154757 402190 158148 402192
rect 154757 402187 154823 402190
rect 220721 402114 220787 402117
rect 217948 402112 220787 402114
rect 217948 402056 220726 402112
rect 220782 402056 220787 402112
rect 217948 402054 220787 402056
rect 220721 402051 220787 402054
rect 155217 401978 155283 401981
rect 251173 401978 251239 401981
rect 155217 401976 158148 401978
rect 155217 401920 155222 401976
rect 155278 401920 158148 401976
rect 155217 401918 158148 401920
rect 251173 401976 253644 401978
rect 251173 401920 251178 401976
rect 251234 401920 253644 401976
rect 251173 401918 253644 401920
rect 155217 401915 155283 401918
rect 251173 401915 251239 401918
rect 154941 401706 155007 401709
rect 220169 401706 220235 401709
rect 154941 401704 158148 401706
rect 154941 401648 154946 401704
rect 155002 401648 158148 401704
rect 154941 401646 158148 401648
rect 217948 401704 220235 401706
rect 217948 401648 220174 401704
rect 220230 401648 220235 401704
rect 217948 401646 220235 401648
rect 154941 401643 155007 401646
rect 220169 401643 220235 401646
rect 155125 401434 155191 401437
rect 155125 401432 158148 401434
rect 155125 401376 155130 401432
rect 155186 401376 158148 401432
rect 155125 401374 158148 401376
rect 155125 401371 155191 401374
rect 220077 401298 220143 401301
rect 217948 401296 220143 401298
rect 217948 401240 220082 401296
rect 220138 401240 220143 401296
rect 217948 401238 220143 401240
rect 220077 401235 220143 401238
rect 154849 401162 154915 401165
rect 154849 401160 158148 401162
rect 154849 401104 154854 401160
rect 154910 401104 158148 401160
rect 154849 401102 158148 401104
rect 154849 401099 154915 401102
rect 154941 400890 155007 400893
rect 220721 400890 220787 400893
rect 154941 400888 158148 400890
rect 154941 400832 154946 400888
rect 155002 400832 158148 400888
rect 154941 400830 158148 400832
rect 217948 400888 220787 400890
rect 217948 400832 220726 400888
rect 220782 400832 220787 400888
rect 217948 400830 220787 400832
rect 154941 400827 155007 400830
rect 220721 400827 220787 400830
rect 251909 400754 251975 400757
rect 251909 400752 253644 400754
rect 251909 400696 251914 400752
rect 251970 400696 253644 400752
rect 251909 400694 253644 400696
rect 251909 400691 251975 400694
rect 155217 400618 155283 400621
rect 155217 400616 158148 400618
rect 155217 400560 155222 400616
rect 155278 400560 158148 400616
rect 155217 400558 158148 400560
rect 155217 400555 155283 400558
rect 220169 400482 220235 400485
rect 217948 400480 220235 400482
rect 217948 400424 220174 400480
rect 220230 400424 220235 400480
rect 217948 400422 220235 400424
rect 220169 400419 220235 400422
rect 155033 400346 155099 400349
rect 155033 400344 158148 400346
rect 155033 400288 155038 400344
rect 155094 400288 158148 400344
rect 155033 400286 158148 400288
rect 155033 400283 155099 400286
rect 154941 400074 155007 400077
rect 219985 400074 220051 400077
rect 154941 400072 158148 400074
rect 154941 400016 154946 400072
rect 155002 400016 158148 400072
rect 154941 400014 158148 400016
rect 217948 400072 220051 400074
rect 217948 400016 219990 400072
rect 220046 400016 220051 400072
rect 217948 400014 220051 400016
rect 154941 400011 155007 400014
rect 219985 400011 220051 400014
rect 154849 399802 154915 399805
rect 154849 399800 158148 399802
rect 154849 399744 154854 399800
rect 154910 399744 158148 399800
rect 154849 399742 158148 399744
rect 154849 399739 154915 399742
rect 220721 399666 220787 399669
rect 217948 399664 220787 399666
rect 217948 399608 220726 399664
rect 220782 399608 220787 399664
rect 217948 399606 220787 399608
rect 220721 399603 220787 399606
rect 155033 399530 155099 399533
rect 251173 399530 251239 399533
rect 155033 399528 158148 399530
rect 155033 399472 155038 399528
rect 155094 399472 158148 399528
rect 155033 399470 158148 399472
rect 251173 399528 253644 399530
rect 251173 399472 251178 399528
rect 251234 399472 253644 399528
rect 251173 399470 253644 399472
rect 155033 399467 155099 399470
rect 251173 399467 251239 399470
rect 154757 399258 154823 399261
rect 220077 399258 220143 399261
rect 154757 399256 158148 399258
rect 154757 399200 154762 399256
rect 154818 399200 158148 399256
rect 154757 399198 158148 399200
rect 217948 399256 220143 399258
rect 217948 399200 220082 399256
rect 220138 399200 220143 399256
rect 217948 399198 220143 399200
rect 154757 399195 154823 399198
rect 220077 399195 220143 399198
rect 155125 398986 155191 398989
rect 155125 398984 158148 398986
rect 155125 398928 155130 398984
rect 155186 398928 158148 398984
rect 155125 398926 158148 398928
rect 155125 398923 155191 398926
rect 220169 398850 220235 398853
rect 217948 398848 220235 398850
rect 217948 398792 220174 398848
rect 220230 398792 220235 398848
rect 217948 398790 220235 398792
rect 220169 398787 220235 398790
rect 154941 398714 155007 398717
rect 154941 398712 158148 398714
rect 154941 398656 154946 398712
rect 155002 398656 158148 398712
rect 154941 398654 158148 398656
rect 154941 398651 155007 398654
rect 154573 398442 154639 398445
rect 220721 398442 220787 398445
rect 154573 398440 158148 398442
rect 154573 398384 154578 398440
rect 154634 398384 158148 398440
rect 154573 398382 158148 398384
rect 217948 398440 220787 398442
rect 217948 398384 220726 398440
rect 220782 398384 220787 398440
rect 217948 398382 220787 398384
rect 154573 398379 154639 398382
rect 220721 398379 220787 398382
rect 251173 398306 251239 398309
rect 251173 398304 253644 398306
rect 251173 398248 251178 398304
rect 251234 398248 253644 398304
rect 251173 398246 253644 398248
rect 251173 398243 251239 398246
rect 154849 398170 154915 398173
rect 154849 398168 158148 398170
rect 154849 398112 154854 398168
rect 154910 398112 158148 398168
rect 154849 398110 158148 398112
rect 154849 398107 154915 398110
rect 220077 398034 220143 398037
rect 217948 398032 220143 398034
rect 217948 397976 220082 398032
rect 220138 397976 220143 398032
rect 217948 397974 220143 397976
rect 220077 397971 220143 397974
rect 155033 397898 155099 397901
rect 155033 397896 158148 397898
rect 155033 397840 155038 397896
rect 155094 397840 158148 397896
rect 155033 397838 158148 397840
rect 155033 397835 155099 397838
rect 154665 397626 154731 397629
rect 220169 397626 220235 397629
rect 154665 397624 158148 397626
rect -960 397490 480 397580
rect 154665 397568 154670 397624
rect 154726 397568 158148 397624
rect 154665 397566 158148 397568
rect 217948 397624 220235 397626
rect 217948 397568 220174 397624
rect 220230 397568 220235 397624
rect 217948 397566 220235 397568
rect 154665 397563 154731 397566
rect 220169 397563 220235 397566
rect 3325 397490 3391 397493
rect -960 397488 3391 397490
rect -960 397432 3330 397488
rect 3386 397432 3391 397488
rect -960 397430 3391 397432
rect -960 397340 480 397430
rect 3325 397427 3391 397430
rect 154941 397354 155007 397357
rect 154941 397352 158148 397354
rect 154941 397296 154946 397352
rect 155002 397296 158148 397352
rect 154941 397294 158148 397296
rect 154941 397291 155007 397294
rect 220721 397218 220787 397221
rect 217948 397216 220787 397218
rect 217948 397160 220726 397216
rect 220782 397160 220787 397216
rect 217948 397158 220787 397160
rect 220721 397155 220787 397158
rect 155033 397082 155099 397085
rect 251173 397082 251239 397085
rect 155033 397080 158148 397082
rect 155033 397024 155038 397080
rect 155094 397024 158148 397080
rect 155033 397022 158148 397024
rect 251173 397080 253644 397082
rect 251173 397024 251178 397080
rect 251234 397024 253644 397080
rect 251173 397022 253644 397024
rect 155033 397019 155099 397022
rect 251173 397019 251239 397022
rect 154849 396810 154915 396813
rect 220721 396810 220787 396813
rect 154849 396808 158148 396810
rect 154849 396752 154854 396808
rect 154910 396752 158148 396808
rect 154849 396750 158148 396752
rect 217948 396808 220787 396810
rect 217948 396752 220726 396808
rect 220782 396752 220787 396808
rect 217948 396750 220787 396752
rect 154849 396747 154915 396750
rect 220721 396747 220787 396750
rect 154757 396538 154823 396541
rect 154757 396536 158148 396538
rect 154757 396480 154762 396536
rect 154818 396480 158148 396536
rect 154757 396478 158148 396480
rect 154757 396475 154823 396478
rect 220169 396402 220235 396405
rect 217948 396400 220235 396402
rect 217948 396344 220174 396400
rect 220230 396344 220235 396400
rect 217948 396342 220235 396344
rect 220169 396339 220235 396342
rect 155125 396266 155191 396269
rect 155125 396264 158148 396266
rect 155125 396208 155130 396264
rect 155186 396208 158148 396264
rect 155125 396206 158148 396208
rect 155125 396203 155191 396206
rect 154941 395994 155007 395997
rect 219893 395994 219959 395997
rect 154941 395992 158148 395994
rect 154941 395936 154946 395992
rect 155002 395936 158148 395992
rect 154941 395934 158148 395936
rect 217948 395992 219959 395994
rect 217948 395936 219898 395992
rect 219954 395936 219959 395992
rect 217948 395934 219959 395936
rect 154941 395931 155007 395934
rect 219893 395931 219959 395934
rect 251173 395858 251239 395861
rect 251173 395856 253644 395858
rect 251173 395800 251178 395856
rect 251234 395800 253644 395856
rect 251173 395798 253644 395800
rect 251173 395795 251239 395798
rect 154665 395722 154731 395725
rect 154665 395720 158148 395722
rect 154665 395664 154670 395720
rect 154726 395664 158148 395720
rect 154665 395662 158148 395664
rect 154665 395659 154731 395662
rect 220077 395586 220143 395589
rect 217948 395584 220143 395586
rect 217948 395528 220082 395584
rect 220138 395528 220143 395584
rect 217948 395526 220143 395528
rect 220077 395523 220143 395526
rect 154849 395450 154915 395453
rect 154849 395448 158148 395450
rect 154849 395392 154854 395448
rect 154910 395392 158148 395448
rect 154849 395390 158148 395392
rect 154849 395387 154915 395390
rect 154757 395178 154823 395181
rect 220169 395178 220235 395181
rect 154757 395176 158148 395178
rect 154757 395120 154762 395176
rect 154818 395120 158148 395176
rect 154757 395118 158148 395120
rect 217948 395176 220235 395178
rect 217948 395120 220174 395176
rect 220230 395120 220235 395176
rect 217948 395118 220235 395120
rect 154757 395115 154823 395118
rect 220169 395115 220235 395118
rect 155033 394906 155099 394909
rect 155033 394904 158148 394906
rect 155033 394848 155038 394904
rect 155094 394848 158148 394904
rect 155033 394846 158148 394848
rect 155033 394843 155099 394846
rect 220721 394770 220787 394773
rect 217948 394768 220787 394770
rect 217948 394712 220726 394768
rect 220782 394712 220787 394768
rect 217948 394710 220787 394712
rect 220721 394707 220787 394710
rect 154665 394634 154731 394637
rect 251633 394634 251699 394637
rect 154665 394632 158148 394634
rect 154665 394576 154670 394632
rect 154726 394576 158148 394632
rect 154665 394574 158148 394576
rect 251633 394632 253644 394634
rect 251633 394576 251638 394632
rect 251694 394576 253644 394632
rect 251633 394574 253644 394576
rect 154665 394571 154731 394574
rect 251633 394571 251699 394574
rect 154573 394362 154639 394365
rect 220721 394362 220787 394365
rect 154573 394360 158148 394362
rect 154573 394304 154578 394360
rect 154634 394304 158148 394360
rect 154573 394302 158148 394304
rect 217948 394360 220787 394362
rect 217948 394304 220726 394360
rect 220782 394304 220787 394360
rect 217948 394302 220787 394304
rect 154573 394299 154639 394302
rect 220721 394299 220787 394302
rect 154757 394090 154823 394093
rect 154757 394088 158148 394090
rect 154757 394032 154762 394088
rect 154818 394032 158148 394088
rect 154757 394030 158148 394032
rect 154757 394027 154823 394030
rect 219985 393954 220051 393957
rect 217948 393952 220051 393954
rect 217948 393896 219990 393952
rect 220046 393896 220051 393952
rect 217948 393894 220051 393896
rect 219985 393891 220051 393894
rect 154941 393818 155007 393821
rect 154941 393816 158148 393818
rect 154941 393760 154946 393816
rect 155002 393760 158148 393816
rect 154941 393758 158148 393760
rect 154941 393755 155007 393758
rect 154849 393546 154915 393549
rect 220169 393546 220235 393549
rect 154849 393544 158148 393546
rect 154849 393488 154854 393544
rect 154910 393488 158148 393544
rect 154849 393486 158148 393488
rect 217948 393544 220235 393546
rect 217948 393488 220174 393544
rect 220230 393488 220235 393544
rect 217948 393486 220235 393488
rect 154849 393483 154915 393486
rect 220169 393483 220235 393486
rect 251173 393410 251239 393413
rect 251173 393408 253644 393410
rect 251173 393352 251178 393408
rect 251234 393352 253644 393408
rect 251173 393350 253644 393352
rect 251173 393347 251239 393350
rect 154941 393274 155007 393277
rect 154941 393272 158148 393274
rect 154941 393216 154946 393272
rect 155002 393216 158148 393272
rect 154941 393214 158148 393216
rect 154941 393211 155007 393214
rect 220721 393138 220787 393141
rect 217948 393136 220787 393138
rect 217948 393080 220726 393136
rect 220782 393080 220787 393136
rect 217948 393078 220787 393080
rect 220721 393075 220787 393078
rect 155033 393002 155099 393005
rect 155033 393000 158148 393002
rect 155033 392944 155038 393000
rect 155094 392944 158148 393000
rect 155033 392942 158148 392944
rect 155033 392939 155099 392942
rect 154941 392730 155007 392733
rect 220261 392730 220327 392733
rect 154941 392728 158148 392730
rect 154941 392672 154946 392728
rect 155002 392672 158148 392728
rect 154941 392670 158148 392672
rect 217948 392728 220327 392730
rect 217948 392672 220266 392728
rect 220322 392672 220327 392728
rect 217948 392670 220327 392672
rect 154941 392667 155007 392670
rect 220261 392667 220327 392670
rect 154849 392458 154915 392461
rect 154849 392456 158148 392458
rect 154849 392400 154854 392456
rect 154910 392400 158148 392456
rect 154849 392398 158148 392400
rect 154849 392395 154915 392398
rect 220169 392322 220235 392325
rect 217948 392320 220235 392322
rect 217948 392264 220174 392320
rect 220230 392264 220235 392320
rect 217948 392262 220235 392264
rect 220169 392259 220235 392262
rect 154757 392186 154823 392189
rect 251173 392186 251239 392189
rect 154757 392184 158148 392186
rect 154757 392128 154762 392184
rect 154818 392128 158148 392184
rect 154757 392126 158148 392128
rect 251173 392184 253644 392186
rect 251173 392128 251178 392184
rect 251234 392128 253644 392184
rect 251173 392126 253644 392128
rect 154757 392123 154823 392126
rect 251173 392123 251239 392126
rect 154941 391914 155007 391917
rect 220721 391914 220787 391917
rect 154941 391912 158148 391914
rect 154941 391856 154946 391912
rect 155002 391856 158148 391912
rect 154941 391854 158148 391856
rect 217948 391912 220787 391914
rect 217948 391856 220726 391912
rect 220782 391856 220787 391912
rect 217948 391854 220787 391856
rect 154941 391851 155007 391854
rect 220721 391851 220787 391854
rect 154665 391642 154731 391645
rect 154665 391640 158148 391642
rect 154665 391584 154670 391640
rect 154726 391584 158148 391640
rect 583520 391628 584960 391868
rect 154665 391582 158148 391584
rect 154665 391579 154731 391582
rect 220721 391506 220787 391509
rect 217948 391504 220787 391506
rect 217948 391448 220726 391504
rect 220782 391448 220787 391504
rect 217948 391446 220787 391448
rect 220721 391443 220787 391446
rect 154757 391370 154823 391373
rect 154757 391368 158148 391370
rect 154757 391312 154762 391368
rect 154818 391312 158148 391368
rect 154757 391310 158148 391312
rect 154757 391307 154823 391310
rect 154941 391098 155007 391101
rect 220261 391098 220327 391101
rect 154941 391096 158148 391098
rect 154941 391040 154946 391096
rect 155002 391040 158148 391096
rect 154941 391038 158148 391040
rect 217948 391096 220327 391098
rect 217948 391040 220266 391096
rect 220322 391040 220327 391096
rect 217948 391038 220327 391040
rect 154941 391035 155007 391038
rect 220261 391035 220327 391038
rect 251173 390962 251239 390965
rect 251173 390960 253644 390962
rect 251173 390904 251178 390960
rect 251234 390904 253644 390960
rect 251173 390902 253644 390904
rect 251173 390899 251239 390902
rect 153837 390826 153903 390829
rect 153837 390824 158148 390826
rect 153837 390768 153842 390824
rect 153898 390768 158148 390824
rect 153837 390766 158148 390768
rect 153837 390763 153903 390766
rect 220445 390690 220511 390693
rect 217948 390688 220511 390690
rect 217948 390632 220450 390688
rect 220506 390632 220511 390688
rect 217948 390630 220511 390632
rect 220445 390627 220511 390630
rect 154941 390554 155007 390557
rect 154941 390552 158148 390554
rect 154941 390496 154946 390552
rect 155002 390496 158148 390552
rect 154941 390494 158148 390496
rect 154941 390491 155007 390494
rect 155217 390282 155283 390285
rect 220721 390282 220787 390285
rect 155217 390280 158148 390282
rect 155217 390224 155222 390280
rect 155278 390224 158148 390280
rect 155217 390222 158148 390224
rect 217948 390280 220787 390282
rect 217948 390224 220726 390280
rect 220782 390224 220787 390280
rect 217948 390222 220787 390224
rect 155217 390219 155283 390222
rect 220721 390219 220787 390222
rect 154941 390010 155007 390013
rect 154941 390008 158148 390010
rect 154941 389952 154946 390008
rect 155002 389952 158148 390008
rect 154941 389950 158148 389952
rect 154941 389947 155007 389950
rect 219893 389874 219959 389877
rect 217948 389872 219959 389874
rect 217948 389816 219898 389872
rect 219954 389816 219959 389872
rect 217948 389814 219959 389816
rect 219893 389811 219959 389814
rect 154849 389738 154915 389741
rect 251173 389738 251239 389741
rect 154849 389736 158148 389738
rect 154849 389680 154854 389736
rect 154910 389680 158148 389736
rect 154849 389678 158148 389680
rect 251173 389736 253644 389738
rect 251173 389680 251178 389736
rect 251234 389680 253644 389736
rect 251173 389678 253644 389680
rect 154849 389675 154915 389678
rect 251173 389675 251239 389678
rect 154573 389466 154639 389469
rect 220353 389466 220419 389469
rect 154573 389464 158148 389466
rect 154573 389408 154578 389464
rect 154634 389408 158148 389464
rect 154573 389406 158148 389408
rect 217948 389464 220419 389466
rect 217948 389408 220358 389464
rect 220414 389408 220419 389464
rect 217948 389406 220419 389408
rect 154573 389403 154639 389406
rect 220353 389403 220419 389406
rect 155033 389194 155099 389197
rect 155033 389192 158148 389194
rect 155033 389136 155038 389192
rect 155094 389136 158148 389192
rect 155033 389134 158148 389136
rect 155033 389131 155099 389134
rect 220721 389058 220787 389061
rect 217948 389056 220787 389058
rect 217948 389000 220726 389056
rect 220782 389000 220787 389056
rect 217948 388998 220787 389000
rect 220721 388995 220787 388998
rect 154665 388922 154731 388925
rect 154665 388920 158148 388922
rect 154665 388864 154670 388920
rect 154726 388864 158148 388920
rect 154665 388862 158148 388864
rect 154665 388859 154731 388862
rect 154757 388650 154823 388653
rect 220445 388650 220511 388653
rect 154757 388648 158148 388650
rect 154757 388592 154762 388648
rect 154818 388592 158148 388648
rect 154757 388590 158148 388592
rect 217948 388648 220511 388650
rect 217948 388592 220450 388648
rect 220506 388592 220511 388648
rect 217948 388590 220511 388592
rect 154757 388587 154823 388590
rect 220445 388587 220511 388590
rect 251449 388514 251515 388517
rect 251449 388512 253644 388514
rect 251449 388456 251454 388512
rect 251510 388456 253644 388512
rect 251449 388454 253644 388456
rect 251449 388451 251515 388454
rect 154941 388378 155007 388381
rect 154941 388376 158148 388378
rect 154941 388320 154946 388376
rect 155002 388320 158148 388376
rect 154941 388318 158148 388320
rect 154941 388315 155007 388318
rect 220077 388242 220143 388245
rect 217948 388240 220143 388242
rect 217948 388184 220082 388240
rect 220138 388184 220143 388240
rect 217948 388182 220143 388184
rect 220077 388179 220143 388182
rect 154849 388106 154915 388109
rect 154849 388104 158148 388106
rect 154849 388048 154854 388104
rect 154910 388048 158148 388104
rect 154849 388046 158148 388048
rect 154849 388043 154915 388046
rect 155217 387834 155283 387837
rect 220169 387834 220235 387837
rect 155217 387832 158148 387834
rect 155217 387776 155222 387832
rect 155278 387776 158148 387832
rect 155217 387774 158148 387776
rect 217948 387832 220235 387834
rect 217948 387776 220174 387832
rect 220230 387776 220235 387832
rect 217948 387774 220235 387776
rect 155217 387771 155283 387774
rect 220169 387771 220235 387774
rect 154941 387562 155007 387565
rect 154941 387560 158148 387562
rect 154941 387504 154946 387560
rect 155002 387504 158148 387560
rect 154941 387502 158148 387504
rect 154941 387499 155007 387502
rect 220721 387426 220787 387429
rect 217948 387424 220787 387426
rect 217948 387368 220726 387424
rect 220782 387368 220787 387424
rect 217948 387366 220787 387368
rect 220721 387363 220787 387366
rect 154849 387290 154915 387293
rect 251725 387290 251791 387293
rect 154849 387288 158148 387290
rect 154849 387232 154854 387288
rect 154910 387232 158148 387288
rect 154849 387230 158148 387232
rect 251725 387288 253644 387290
rect 251725 387232 251730 387288
rect 251786 387232 253644 387288
rect 251725 387230 253644 387232
rect 154849 387227 154915 387230
rect 251725 387227 251791 387230
rect 155033 387018 155099 387021
rect 220261 387018 220327 387021
rect 155033 387016 158148 387018
rect 155033 386960 155038 387016
rect 155094 386960 158148 387016
rect 155033 386958 158148 386960
rect 217948 387016 220327 387018
rect 217948 386960 220266 387016
rect 220322 386960 220327 387016
rect 217948 386958 220327 386960
rect 155033 386955 155099 386958
rect 220261 386955 220327 386958
rect 154757 386746 154823 386749
rect 154757 386744 158148 386746
rect 154757 386688 154762 386744
rect 154818 386688 158148 386744
rect 154757 386686 158148 386688
rect 154757 386683 154823 386686
rect 220445 386610 220511 386613
rect 217948 386608 220511 386610
rect 217948 386552 220450 386608
rect 220506 386552 220511 386608
rect 217948 386550 220511 386552
rect 220445 386547 220511 386550
rect 155125 386474 155191 386477
rect 155125 386472 158148 386474
rect 155125 386416 155130 386472
rect 155186 386416 158148 386472
rect 155125 386414 158148 386416
rect 155125 386411 155191 386414
rect 154941 386202 155007 386205
rect 220721 386202 220787 386205
rect 154941 386200 158148 386202
rect 154941 386144 154946 386200
rect 155002 386144 158148 386200
rect 154941 386142 158148 386144
rect 217948 386200 220787 386202
rect 217948 386144 220726 386200
rect 220782 386144 220787 386200
rect 217948 386142 220787 386144
rect 154941 386139 155007 386142
rect 220721 386139 220787 386142
rect 251449 386066 251515 386069
rect 251449 386064 253644 386066
rect 251449 386008 251454 386064
rect 251510 386008 253644 386064
rect 251449 386006 253644 386008
rect 251449 386003 251515 386006
rect 154665 385930 154731 385933
rect 154665 385928 158148 385930
rect 154665 385872 154670 385928
rect 154726 385872 158148 385928
rect 154665 385870 158148 385872
rect 154665 385867 154731 385870
rect 220169 385794 220235 385797
rect 217948 385792 220235 385794
rect 217948 385736 220174 385792
rect 220230 385736 220235 385792
rect 217948 385734 220235 385736
rect 220169 385731 220235 385734
rect 155309 385658 155375 385661
rect 155309 385656 158148 385658
rect 155309 385600 155314 385656
rect 155370 385600 158148 385656
rect 155309 385598 158148 385600
rect 155309 385595 155375 385598
rect 154849 385386 154915 385389
rect 220445 385386 220511 385389
rect 154849 385384 158148 385386
rect 154849 385328 154854 385384
rect 154910 385328 158148 385384
rect 154849 385326 158148 385328
rect 217948 385384 220511 385386
rect 217948 385328 220450 385384
rect 220506 385328 220511 385384
rect 217948 385326 220511 385328
rect 154849 385323 154915 385326
rect 220445 385323 220511 385326
rect 155033 385114 155099 385117
rect 155033 385112 158148 385114
rect 155033 385056 155038 385112
rect 155094 385056 158148 385112
rect 155033 385054 158148 385056
rect 155033 385051 155099 385054
rect 220353 384978 220419 384981
rect 217948 384976 220419 384978
rect 217948 384920 220358 384976
rect 220414 384920 220419 384976
rect 217948 384918 220419 384920
rect 220353 384915 220419 384918
rect 154941 384842 155007 384845
rect 251173 384842 251239 384845
rect 154941 384840 158148 384842
rect 154941 384784 154946 384840
rect 155002 384784 158148 384840
rect 154941 384782 158148 384784
rect 251173 384840 253644 384842
rect 251173 384784 251178 384840
rect 251234 384784 253644 384840
rect 251173 384782 253644 384784
rect 154941 384779 155007 384782
rect 251173 384779 251239 384782
rect 155033 384570 155099 384573
rect 220721 384570 220787 384573
rect 155033 384568 158148 384570
rect -960 384284 480 384524
rect 155033 384512 155038 384568
rect 155094 384512 158148 384568
rect 155033 384510 158148 384512
rect 217948 384568 220787 384570
rect 217948 384512 220726 384568
rect 220782 384512 220787 384568
rect 217948 384510 220787 384512
rect 155033 384507 155099 384510
rect 220721 384507 220787 384510
rect 155125 384298 155191 384301
rect 155125 384296 158148 384298
rect 155125 384240 155130 384296
rect 155186 384240 158148 384296
rect 155125 384238 158148 384240
rect 155125 384235 155191 384238
rect 220261 384162 220327 384165
rect 217948 384160 220327 384162
rect 217948 384104 220266 384160
rect 220322 384104 220327 384160
rect 217948 384102 220327 384104
rect 220261 384099 220327 384102
rect 154849 384026 154915 384029
rect 154849 384024 158148 384026
rect 154849 383968 154854 384024
rect 154910 383968 158148 384024
rect 154849 383966 158148 383968
rect 154849 383963 154915 383966
rect 154665 383754 154731 383757
rect 220445 383754 220511 383757
rect 154665 383752 158148 383754
rect 154665 383696 154670 383752
rect 154726 383696 158148 383752
rect 154665 383694 158148 383696
rect 217948 383752 220511 383754
rect 217948 383696 220450 383752
rect 220506 383696 220511 383752
rect 217948 383694 220511 383696
rect 154665 383691 154731 383694
rect 220445 383691 220511 383694
rect 251173 383618 251239 383621
rect 251173 383616 253644 383618
rect 251173 383560 251178 383616
rect 251234 383560 253644 383616
rect 251173 383558 253644 383560
rect 251173 383555 251239 383558
rect 154941 383482 155007 383485
rect 154941 383480 158148 383482
rect 154941 383424 154946 383480
rect 155002 383424 158148 383480
rect 154941 383422 158148 383424
rect 154941 383419 155007 383422
rect 220077 383346 220143 383349
rect 217948 383344 220143 383346
rect 217948 383288 220082 383344
rect 220138 383288 220143 383344
rect 217948 383286 220143 383288
rect 220077 383283 220143 383286
rect 154849 383210 154915 383213
rect 154849 383208 158148 383210
rect 154849 383152 154854 383208
rect 154910 383152 158148 383208
rect 154849 383150 158148 383152
rect 154849 383147 154915 383150
rect 153929 382938 153995 382941
rect 220445 382938 220511 382941
rect 153929 382936 158148 382938
rect 153929 382880 153934 382936
rect 153990 382880 158148 382936
rect 153929 382878 158148 382880
rect 217948 382936 220511 382938
rect 217948 382880 220450 382936
rect 220506 382880 220511 382936
rect 217948 382878 220511 382880
rect 153929 382875 153995 382878
rect 220445 382875 220511 382878
rect 154941 382666 155007 382669
rect 154941 382664 158148 382666
rect 154941 382608 154946 382664
rect 155002 382608 158148 382664
rect 154941 382606 158148 382608
rect 154941 382603 155007 382606
rect 220537 382530 220603 382533
rect 217948 382528 220603 382530
rect 217948 382472 220542 382528
rect 220598 382472 220603 382528
rect 217948 382470 220603 382472
rect 220537 382467 220603 382470
rect 154665 382394 154731 382397
rect 154665 382392 158148 382394
rect 154665 382336 154670 382392
rect 154726 382336 158148 382392
rect 154665 382334 158148 382336
rect 154665 382331 154731 382334
rect 154941 382122 155007 382125
rect 220721 382122 220787 382125
rect 154941 382120 158148 382122
rect 154941 382064 154946 382120
rect 155002 382064 158148 382120
rect 154941 382062 158148 382064
rect 217948 382120 220787 382122
rect 217948 382064 220726 382120
rect 220782 382064 220787 382120
rect 217948 382062 220787 382064
rect 154941 382059 155007 382062
rect 220721 382059 220787 382062
rect 154573 381850 154639 381853
rect 154573 381848 158148 381850
rect 154573 381792 154578 381848
rect 154634 381792 158148 381848
rect 154573 381790 158148 381792
rect 154573 381787 154639 381790
rect 220629 381714 220695 381717
rect 217948 381712 220695 381714
rect 217948 381656 220634 381712
rect 220690 381656 220695 381712
rect 217948 381654 220695 381656
rect 220629 381651 220695 381654
rect 154849 381578 154915 381581
rect 154849 381576 158148 381578
rect 154849 381520 154854 381576
rect 154910 381520 158148 381576
rect 154849 381518 158148 381520
rect 154849 381515 154915 381518
rect 154941 381306 155007 381309
rect 220537 381306 220603 381309
rect 154941 381304 158148 381306
rect 154941 381248 154946 381304
rect 155002 381248 158148 381304
rect 154941 381246 158148 381248
rect 217948 381304 220603 381306
rect 217948 381248 220542 381304
rect 220598 381248 220603 381304
rect 217948 381246 220603 381248
rect 154941 381243 155007 381246
rect 220537 381243 220603 381246
rect 155493 381034 155559 381037
rect 155493 381032 158148 381034
rect 155493 380976 155498 381032
rect 155554 380976 158148 381032
rect 155493 380974 158148 380976
rect 155493 380971 155559 380974
rect 220721 380898 220787 380901
rect 217948 380896 220787 380898
rect 217948 380840 220726 380896
rect 220782 380840 220787 380896
rect 217948 380838 220787 380840
rect 220721 380835 220787 380838
rect 154941 380762 155007 380765
rect 154941 380760 158148 380762
rect 154941 380704 154946 380760
rect 155002 380704 158148 380760
rect 154941 380702 158148 380704
rect 154941 380699 155007 380702
rect 154941 380490 155007 380493
rect 220721 380490 220787 380493
rect 154941 380488 158148 380490
rect 154941 380432 154946 380488
rect 155002 380432 158148 380488
rect 154941 380430 158148 380432
rect 217948 380488 220787 380490
rect 217948 380432 220726 380488
rect 220782 380432 220787 380488
rect 217948 380430 220787 380432
rect 154941 380427 155007 380430
rect 220721 380427 220787 380430
rect 154849 380218 154915 380221
rect 154849 380216 158148 380218
rect 154849 380160 154854 380216
rect 154910 380160 158148 380216
rect 154849 380158 158148 380160
rect 154849 380155 154915 380158
rect 219709 380082 219775 380085
rect 217948 380080 219775 380082
rect 217948 380024 219714 380080
rect 219770 380024 219775 380080
rect 217948 380022 219775 380024
rect 219709 380019 219775 380022
rect 154757 379946 154823 379949
rect 154757 379944 158148 379946
rect 154757 379888 154762 379944
rect 154818 379888 158148 379944
rect 154757 379886 158148 379888
rect 154757 379883 154823 379886
rect 155033 379674 155099 379677
rect 220629 379674 220695 379677
rect 155033 379672 158148 379674
rect 155033 379616 155038 379672
rect 155094 379616 158148 379672
rect 155033 379614 158148 379616
rect 217948 379672 220695 379674
rect 217948 379616 220634 379672
rect 220690 379616 220695 379672
rect 217948 379614 220695 379616
rect 155033 379611 155099 379614
rect 220629 379611 220695 379614
rect 154941 379402 155007 379405
rect 154941 379400 158148 379402
rect 154941 379344 154946 379400
rect 155002 379344 158148 379400
rect 154941 379342 158148 379344
rect 154941 379339 155007 379342
rect 220721 379266 220787 379269
rect 217948 379264 220787 379266
rect 217948 379208 220726 379264
rect 220782 379208 220787 379264
rect 217948 379206 220787 379208
rect 220721 379203 220787 379206
rect 154849 379130 154915 379133
rect 154849 379128 158148 379130
rect 154849 379072 154854 379128
rect 154910 379072 158148 379128
rect 154849 379070 158148 379072
rect 154849 379067 154915 379070
rect 154941 378858 155007 378861
rect 220537 378858 220603 378861
rect 154941 378856 158148 378858
rect 154941 378800 154946 378856
rect 155002 378800 158148 378856
rect 154941 378798 158148 378800
rect 217948 378856 220603 378858
rect 217948 378800 220542 378856
rect 220598 378800 220603 378856
rect 217948 378798 220603 378800
rect 154941 378795 155007 378798
rect 220537 378795 220603 378798
rect 154021 378586 154087 378589
rect 154021 378584 158148 378586
rect 154021 378528 154026 378584
rect 154082 378528 158148 378584
rect 154021 378526 158148 378528
rect 154021 378523 154087 378526
rect 220629 378450 220695 378453
rect 217948 378448 220695 378450
rect 217948 378392 220634 378448
rect 220690 378392 220695 378448
rect 217948 378390 220695 378392
rect 220629 378387 220695 378390
rect 579797 378450 579863 378453
rect 583520 378450 584960 378540
rect 579797 378448 584960 378450
rect 579797 378392 579802 378448
rect 579858 378392 584960 378448
rect 579797 378390 584960 378392
rect 579797 378387 579863 378390
rect 155033 378314 155099 378317
rect 155033 378312 158148 378314
rect 155033 378256 155038 378312
rect 155094 378256 158148 378312
rect 583520 378300 584960 378390
rect 155033 378254 158148 378256
rect 155033 378251 155099 378254
rect 154941 378042 155007 378045
rect 220721 378042 220787 378045
rect 154941 378040 158148 378042
rect 154941 377984 154946 378040
rect 155002 377984 158148 378040
rect 154941 377982 158148 377984
rect 217948 378040 220787 378042
rect 217948 377984 220726 378040
rect 220782 377984 220787 378040
rect 217948 377982 220787 377984
rect 154941 377979 155007 377982
rect 220721 377979 220787 377982
rect 154941 377770 155007 377773
rect 154941 377768 158148 377770
rect 154941 377712 154946 377768
rect 155002 377712 158148 377768
rect 154941 377710 158148 377712
rect 154941 377707 155007 377710
rect 220629 377634 220695 377637
rect 217948 377632 220695 377634
rect 217948 377576 220634 377632
rect 220690 377576 220695 377632
rect 217948 377574 220695 377576
rect 220629 377571 220695 377574
rect 155033 377498 155099 377501
rect 155033 377496 158148 377498
rect 155033 377440 155038 377496
rect 155094 377440 158148 377496
rect 155033 377438 158148 377440
rect 155033 377435 155099 377438
rect 154757 377226 154823 377229
rect 220537 377226 220603 377229
rect 154757 377224 158148 377226
rect 154757 377168 154762 377224
rect 154818 377168 158148 377224
rect 154757 377166 158148 377168
rect 217948 377224 220603 377226
rect 217948 377168 220542 377224
rect 220598 377168 220603 377224
rect 217948 377166 220603 377168
rect 154757 377163 154823 377166
rect 220537 377163 220603 377166
rect 154849 376954 154915 376957
rect 154849 376952 158148 376954
rect 154849 376896 154854 376952
rect 154910 376896 158148 376952
rect 154849 376894 158148 376896
rect 154849 376891 154915 376894
rect 220445 376818 220511 376821
rect 217948 376816 220511 376818
rect 217948 376760 220450 376816
rect 220506 376760 220511 376816
rect 217948 376758 220511 376760
rect 220445 376755 220511 376758
rect 154941 376682 155007 376685
rect 154941 376680 158148 376682
rect 154941 376624 154946 376680
rect 155002 376624 158148 376680
rect 154941 376622 158148 376624
rect 154941 376619 155007 376622
rect 154941 376410 155007 376413
rect 220721 376410 220787 376413
rect 154941 376408 158148 376410
rect 154941 376352 154946 376408
rect 155002 376352 158148 376408
rect 154941 376350 158148 376352
rect 217948 376408 220787 376410
rect 217948 376352 220726 376408
rect 220782 376352 220787 376408
rect 217948 376350 220787 376352
rect 154941 376347 155007 376350
rect 220721 376347 220787 376350
rect 154849 376138 154915 376141
rect 154849 376136 158148 376138
rect 154849 376080 154854 376136
rect 154910 376080 158148 376136
rect 154849 376078 158148 376080
rect 154849 376075 154915 376078
rect 219985 376002 220051 376005
rect 217948 376000 220051 376002
rect 217948 375944 219990 376000
rect 220046 375944 220051 376000
rect 217948 375942 220051 375944
rect 219985 375939 220051 375942
rect 155033 375866 155099 375869
rect 155033 375864 158148 375866
rect 155033 375808 155038 375864
rect 155094 375808 158148 375864
rect 155033 375806 158148 375808
rect 155033 375803 155099 375806
rect 154665 375594 154731 375597
rect 219985 375594 220051 375597
rect 154665 375592 158148 375594
rect 154665 375536 154670 375592
rect 154726 375536 158148 375592
rect 154665 375534 158148 375536
rect 217948 375592 220051 375594
rect 217948 375536 219990 375592
rect 220046 375536 220051 375592
rect 217948 375534 220051 375536
rect 154665 375531 154731 375534
rect 219985 375531 220051 375534
rect 154941 375322 155007 375325
rect 154941 375320 158148 375322
rect 154941 375264 154946 375320
rect 155002 375264 158148 375320
rect 154941 375262 158148 375264
rect 154941 375259 155007 375262
rect 220721 375186 220787 375189
rect 217948 375184 220787 375186
rect 217948 375128 220726 375184
rect 220782 375128 220787 375184
rect 217948 375126 220787 375128
rect 220721 375123 220787 375126
rect 154849 375050 154915 375053
rect 154849 375048 158148 375050
rect 154849 374992 154854 375048
rect 154910 374992 158148 375048
rect 154849 374990 158148 374992
rect 154849 374987 154915 374990
rect 154573 374778 154639 374781
rect 219433 374778 219499 374781
rect 154573 374776 158148 374778
rect 154573 374720 154578 374776
rect 154634 374720 158148 374776
rect 154573 374718 158148 374720
rect 217948 374776 219499 374778
rect 217948 374720 219438 374776
rect 219494 374720 219499 374776
rect 217948 374718 219499 374720
rect 154573 374715 154639 374718
rect 219433 374715 219499 374718
rect 155125 374506 155191 374509
rect 155125 374504 158148 374506
rect 155125 374448 155130 374504
rect 155186 374448 158148 374504
rect 155125 374446 158148 374448
rect 155125 374443 155191 374446
rect 220629 374370 220695 374373
rect 217948 374368 220695 374370
rect 217948 374312 220634 374368
rect 220690 374312 220695 374368
rect 217948 374310 220695 374312
rect 220629 374307 220695 374310
rect 155401 374234 155467 374237
rect 155401 374232 158148 374234
rect 155401 374176 155406 374232
rect 155462 374176 158148 374232
rect 155401 374174 158148 374176
rect 155401 374171 155467 374174
rect 154573 373962 154639 373965
rect 220537 373962 220603 373965
rect 154573 373960 158148 373962
rect 154573 373904 154578 373960
rect 154634 373904 158148 373960
rect 154573 373902 158148 373904
rect 217948 373960 220603 373962
rect 217948 373904 220542 373960
rect 220598 373904 220603 373960
rect 217948 373902 220603 373904
rect 154573 373899 154639 373902
rect 220537 373899 220603 373902
rect 154941 373690 155007 373693
rect 154941 373688 158148 373690
rect 154941 373632 154946 373688
rect 155002 373632 158148 373688
rect 154941 373630 158148 373632
rect 154941 373627 155007 373630
rect 219893 373554 219959 373557
rect 217948 373552 219959 373554
rect 217948 373496 219898 373552
rect 219954 373496 219959 373552
rect 217948 373494 219959 373496
rect 219893 373491 219959 373494
rect 154849 373418 154915 373421
rect 154849 373416 158148 373418
rect 154849 373360 154854 373416
rect 154910 373360 158148 373416
rect 154849 373358 158148 373360
rect 154849 373355 154915 373358
rect 154757 373146 154823 373149
rect 220629 373146 220695 373149
rect 154757 373144 158148 373146
rect 154757 373088 154762 373144
rect 154818 373088 158148 373144
rect 154757 373086 158148 373088
rect 217948 373144 220695 373146
rect 217948 373088 220634 373144
rect 220690 373088 220695 373144
rect 217948 373086 220695 373088
rect 154757 373083 154823 373086
rect 220629 373083 220695 373086
rect 154665 372874 154731 372877
rect 154665 372872 158148 372874
rect 154665 372816 154670 372872
rect 154726 372816 158148 372872
rect 154665 372814 158148 372816
rect 154665 372811 154731 372814
rect 220721 372738 220787 372741
rect 217948 372736 220787 372738
rect 217948 372680 220726 372736
rect 220782 372680 220787 372736
rect 217948 372678 220787 372680
rect 220721 372675 220787 372678
rect 154941 372602 155007 372605
rect 154941 372600 158148 372602
rect 154941 372544 154946 372600
rect 155002 372544 158148 372600
rect 154941 372542 158148 372544
rect 154941 372539 155007 372542
rect 154757 372330 154823 372333
rect 220353 372330 220419 372333
rect 154757 372328 158148 372330
rect 154757 372272 154762 372328
rect 154818 372272 158148 372328
rect 154757 372270 158148 372272
rect 217948 372328 220419 372330
rect 217948 372272 220358 372328
rect 220414 372272 220419 372328
rect 217948 372270 220419 372272
rect 154757 372267 154823 372270
rect 220353 372267 220419 372270
rect 154941 372058 155007 372061
rect 154941 372056 158148 372058
rect 154941 372000 154946 372056
rect 155002 372000 158148 372056
rect 154941 371998 158148 372000
rect 154941 371995 155007 371998
rect 220445 371922 220511 371925
rect 217948 371920 220511 371922
rect 217948 371864 220450 371920
rect 220506 371864 220511 371920
rect 217948 371862 220511 371864
rect 220445 371859 220511 371862
rect 155125 371786 155191 371789
rect 155125 371784 158148 371786
rect 155125 371728 155130 371784
rect 155186 371728 158148 371784
rect 155125 371726 158148 371728
rect 155125 371723 155191 371726
rect 154849 371514 154915 371517
rect 219985 371514 220051 371517
rect 154849 371512 158148 371514
rect -960 371378 480 371468
rect 154849 371456 154854 371512
rect 154910 371456 158148 371512
rect 154849 371454 158148 371456
rect 217948 371512 220051 371514
rect 217948 371456 219990 371512
rect 220046 371456 220051 371512
rect 217948 371454 220051 371456
rect 154849 371451 154915 371454
rect 219985 371451 220051 371454
rect 3325 371378 3391 371381
rect -960 371376 3391 371378
rect -960 371320 3330 371376
rect 3386 371320 3391 371376
rect -960 371318 3391 371320
rect -960 371228 480 371318
rect 3325 371315 3391 371318
rect 155125 371242 155191 371245
rect 155125 371240 158148 371242
rect 155125 371184 155130 371240
rect 155186 371184 158148 371240
rect 155125 371182 158148 371184
rect 155125 371179 155191 371182
rect 220629 371106 220695 371109
rect 217948 371104 220695 371106
rect 217948 371048 220634 371104
rect 220690 371048 220695 371104
rect 217948 371046 220695 371048
rect 220629 371043 220695 371046
rect 154941 370970 155007 370973
rect 154941 370968 158148 370970
rect 154941 370912 154946 370968
rect 155002 370912 158148 370968
rect 154941 370910 158148 370912
rect 154941 370907 155007 370910
rect 154849 370698 154915 370701
rect 220721 370698 220787 370701
rect 154849 370696 158148 370698
rect 154849 370640 154854 370696
rect 154910 370640 158148 370696
rect 154849 370638 158148 370640
rect 217948 370696 220787 370698
rect 217948 370640 220726 370696
rect 220782 370640 220787 370696
rect 217948 370638 220787 370640
rect 154849 370635 154915 370638
rect 220721 370635 220787 370638
rect 154757 370426 154823 370429
rect 154757 370424 158148 370426
rect 154757 370368 154762 370424
rect 154818 370368 158148 370424
rect 154757 370366 158148 370368
rect 154757 370363 154823 370366
rect 220537 370290 220603 370293
rect 217948 370288 220603 370290
rect 217948 370232 220542 370288
rect 220598 370232 220603 370288
rect 217948 370230 220603 370232
rect 220537 370227 220603 370230
rect 154665 370154 154731 370157
rect 154665 370152 158148 370154
rect 154665 370096 154670 370152
rect 154726 370096 158148 370152
rect 154665 370094 158148 370096
rect 154665 370091 154731 370094
rect 155309 369882 155375 369885
rect 220537 369882 220603 369885
rect 155309 369880 158148 369882
rect 155309 369824 155314 369880
rect 155370 369824 158148 369880
rect 155309 369822 158148 369824
rect 217948 369880 220603 369882
rect 217948 369824 220542 369880
rect 220598 369824 220603 369880
rect 217948 369822 220603 369824
rect 155309 369819 155375 369822
rect 220537 369819 220603 369822
rect 154941 369610 155007 369613
rect 154941 369608 158148 369610
rect 154941 369552 154946 369608
rect 155002 369552 158148 369608
rect 154941 369550 158148 369552
rect 154941 369547 155007 369550
rect 220629 369474 220695 369477
rect 217948 369472 220695 369474
rect 217948 369416 220634 369472
rect 220690 369416 220695 369472
rect 217948 369414 220695 369416
rect 220629 369411 220695 369414
rect 154849 369338 154915 369341
rect 154849 369336 158148 369338
rect 154849 369280 154854 369336
rect 154910 369280 158148 369336
rect 154849 369278 158148 369280
rect 154849 369275 154915 369278
rect 155125 369066 155191 369069
rect 220629 369066 220695 369069
rect 155125 369064 158148 369066
rect 155125 369008 155130 369064
rect 155186 369008 158148 369064
rect 155125 369006 158148 369008
rect 217948 369064 220695 369066
rect 217948 369008 220634 369064
rect 220690 369008 220695 369064
rect 217948 369006 220695 369008
rect 155125 369003 155191 369006
rect 220629 369003 220695 369006
rect 154665 368794 154731 368797
rect 154665 368792 158148 368794
rect 154665 368736 154670 368792
rect 154726 368736 158148 368792
rect 154665 368734 158148 368736
rect 154665 368731 154731 368734
rect 219709 368658 219775 368661
rect 217948 368656 219775 368658
rect 217948 368600 219714 368656
rect 219770 368600 219775 368656
rect 217948 368598 219775 368600
rect 219709 368595 219775 368598
rect 154757 368522 154823 368525
rect 154757 368520 158148 368522
rect 154757 368464 154762 368520
rect 154818 368464 158148 368520
rect 154757 368462 158148 368464
rect 154757 368459 154823 368462
rect 154573 368250 154639 368253
rect 220721 368250 220787 368253
rect 154573 368248 158148 368250
rect 154573 368192 154578 368248
rect 154634 368192 158148 368248
rect 154573 368190 158148 368192
rect 217948 368248 220787 368250
rect 217948 368192 220726 368248
rect 220782 368192 220787 368248
rect 217948 368190 220787 368192
rect 154573 368187 154639 368190
rect 220721 368187 220787 368190
rect 154941 367978 155007 367981
rect 154941 367976 158148 367978
rect 154941 367920 154946 367976
rect 155002 367920 158148 367976
rect 154941 367918 158148 367920
rect 154941 367915 155007 367918
rect 220537 367842 220603 367845
rect 217948 367840 220603 367842
rect 217948 367784 220542 367840
rect 220598 367784 220603 367840
rect 217948 367782 220603 367784
rect 220537 367779 220603 367782
rect 155493 367706 155559 367709
rect 155493 367704 158148 367706
rect 155493 367648 155498 367704
rect 155554 367648 158148 367704
rect 155493 367646 158148 367648
rect 155493 367643 155559 367646
rect 154757 367434 154823 367437
rect 219893 367434 219959 367437
rect 154757 367432 158148 367434
rect 154757 367376 154762 367432
rect 154818 367376 158148 367432
rect 154757 367374 158148 367376
rect 217948 367432 219959 367434
rect 217948 367376 219898 367432
rect 219954 367376 219959 367432
rect 217948 367374 219959 367376
rect 154757 367371 154823 367374
rect 219893 367371 219959 367374
rect 154849 367162 154915 367165
rect 154849 367160 158148 367162
rect 154849 367104 154854 367160
rect 154910 367104 158148 367160
rect 154849 367102 158148 367104
rect 154849 367099 154915 367102
rect 220721 367026 220787 367029
rect 217948 367024 220787 367026
rect 217948 366968 220726 367024
rect 220782 366968 220787 367024
rect 217948 366966 220787 366968
rect 220721 366963 220787 366966
rect 154941 366890 155007 366893
rect 154941 366888 158148 366890
rect 154941 366832 154946 366888
rect 155002 366832 158148 366888
rect 154941 366830 158148 366832
rect 154941 366827 155007 366830
rect 155125 366618 155191 366621
rect 220537 366618 220603 366621
rect 155125 366616 158148 366618
rect 155125 366560 155130 366616
rect 155186 366560 158148 366616
rect 155125 366558 158148 366560
rect 217948 366616 220603 366618
rect 217948 366560 220542 366616
rect 220598 366560 220603 366616
rect 217948 366558 220603 366560
rect 155125 366555 155191 366558
rect 220537 366555 220603 366558
rect 154665 366346 154731 366349
rect 154665 366344 158148 366346
rect 154665 366288 154670 366344
rect 154726 366288 158148 366344
rect 154665 366286 158148 366288
rect 154665 366283 154731 366286
rect 220629 366210 220695 366213
rect 217948 366208 220695 366210
rect 217948 366152 220634 366208
rect 220690 366152 220695 366208
rect 217948 366150 220695 366152
rect 220629 366147 220695 366150
rect 154849 366074 154915 366077
rect 154849 366072 158148 366074
rect 154849 366016 154854 366072
rect 154910 366016 158148 366072
rect 154849 366014 158148 366016
rect 154849 366011 154915 366014
rect 155585 365802 155651 365805
rect 219617 365802 219683 365805
rect 155585 365800 158148 365802
rect 155585 365744 155590 365800
rect 155646 365744 158148 365800
rect 155585 365742 158148 365744
rect 217948 365800 219683 365802
rect 217948 365744 219622 365800
rect 219678 365744 219683 365800
rect 217948 365742 219683 365744
rect 155585 365739 155651 365742
rect 219617 365739 219683 365742
rect 154665 365530 154731 365533
rect 154665 365528 158148 365530
rect 154665 365472 154670 365528
rect 154726 365472 158148 365528
rect 154665 365470 158148 365472
rect 154665 365467 154731 365470
rect 219985 365394 220051 365397
rect 217948 365392 220051 365394
rect 217948 365336 219990 365392
rect 220046 365336 220051 365392
rect 217948 365334 220051 365336
rect 219985 365331 220051 365334
rect 154941 365258 155007 365261
rect 154941 365256 158148 365258
rect 154941 365200 154946 365256
rect 155002 365200 158148 365256
rect 154941 365198 158148 365200
rect 154941 365195 155007 365198
rect 579981 365122 580047 365125
rect 583520 365122 584960 365212
rect 579981 365120 584960 365122
rect 579981 365064 579986 365120
rect 580042 365064 584960 365120
rect 579981 365062 584960 365064
rect 579981 365059 580047 365062
rect 154757 364986 154823 364989
rect 220629 364986 220695 364989
rect 154757 364984 158148 364986
rect 154757 364928 154762 364984
rect 154818 364928 158148 364984
rect 154757 364926 158148 364928
rect 217948 364984 220695 364986
rect 217948 364928 220634 364984
rect 220690 364928 220695 364984
rect 583520 364972 584960 365062
rect 217948 364926 220695 364928
rect 154757 364923 154823 364926
rect 220629 364923 220695 364926
rect 154849 364714 154915 364717
rect 154849 364712 158148 364714
rect 154849 364656 154854 364712
rect 154910 364656 158148 364712
rect 154849 364654 158148 364656
rect 154849 364651 154915 364654
rect 219709 364578 219775 364581
rect 217948 364576 219775 364578
rect 217948 364520 219714 364576
rect 219770 364520 219775 364576
rect 217948 364518 219775 364520
rect 219709 364515 219775 364518
rect 155125 364442 155191 364445
rect 155125 364440 158148 364442
rect 155125 364384 155130 364440
rect 155186 364384 158148 364440
rect 155125 364382 158148 364384
rect 155125 364379 155191 364382
rect 154941 364170 155007 364173
rect 220537 364170 220603 364173
rect 154941 364168 158148 364170
rect 154941 364112 154946 364168
rect 155002 364112 158148 364168
rect 154941 364110 158148 364112
rect 217948 364168 220603 364170
rect 217948 364112 220542 364168
rect 220598 364112 220603 364168
rect 217948 364110 220603 364112
rect 154941 364107 155007 364110
rect 220537 364107 220603 364110
rect 154757 363898 154823 363901
rect 154757 363896 158148 363898
rect 154757 363840 154762 363896
rect 154818 363840 158148 363896
rect 154757 363838 158148 363840
rect 154757 363835 154823 363838
rect 220721 363762 220787 363765
rect 217948 363760 220787 363762
rect 217948 363704 220726 363760
rect 220782 363704 220787 363760
rect 217948 363702 220787 363704
rect 220721 363699 220787 363702
rect 154849 363626 154915 363629
rect 154849 363624 158148 363626
rect 154849 363568 154854 363624
rect 154910 363568 158148 363624
rect 154849 363566 158148 363568
rect 154849 363563 154915 363566
rect 155033 363354 155099 363357
rect 220629 363354 220695 363357
rect 155033 363352 158148 363354
rect 155033 363296 155038 363352
rect 155094 363296 158148 363352
rect 155033 363294 158148 363296
rect 217948 363352 220695 363354
rect 217948 363296 220634 363352
rect 220690 363296 220695 363352
rect 217948 363294 220695 363296
rect 155033 363291 155099 363294
rect 220629 363291 220695 363294
rect 155217 363082 155283 363085
rect 155217 363080 158148 363082
rect 155217 363024 155222 363080
rect 155278 363024 158148 363080
rect 155217 363022 158148 363024
rect 155217 363019 155283 363022
rect 220721 362946 220787 362949
rect 217948 362944 220787 362946
rect 217948 362888 220726 362944
rect 220782 362888 220787 362944
rect 217948 362886 220787 362888
rect 220721 362883 220787 362886
rect 154941 362810 155007 362813
rect 154941 362808 158148 362810
rect 154941 362752 154946 362808
rect 155002 362752 158148 362808
rect 154941 362750 158148 362752
rect 154941 362747 155007 362750
rect 155401 362538 155467 362541
rect 220629 362538 220695 362541
rect 155401 362536 158148 362538
rect 155401 362480 155406 362536
rect 155462 362480 158148 362536
rect 155401 362478 158148 362480
rect 217948 362536 220695 362538
rect 217948 362480 220634 362536
rect 220690 362480 220695 362536
rect 217948 362478 220695 362480
rect 155401 362475 155467 362478
rect 220629 362475 220695 362478
rect 154849 362266 154915 362269
rect 154849 362264 158148 362266
rect 154849 362208 154854 362264
rect 154910 362208 158148 362264
rect 154849 362206 158148 362208
rect 154849 362203 154915 362206
rect 220445 362130 220511 362133
rect 217948 362128 220511 362130
rect 217948 362072 220450 362128
rect 220506 362072 220511 362128
rect 217948 362070 220511 362072
rect 220445 362067 220511 362070
rect 155033 361994 155099 361997
rect 155033 361992 158148 361994
rect 155033 361936 155038 361992
rect 155094 361936 158148 361992
rect 155033 361934 158148 361936
rect 155033 361931 155099 361934
rect 154573 361722 154639 361725
rect 220537 361722 220603 361725
rect 154573 361720 158148 361722
rect 154573 361664 154578 361720
rect 154634 361664 158148 361720
rect 154573 361662 158148 361664
rect 217948 361720 220603 361722
rect 217948 361664 220542 361720
rect 220598 361664 220603 361720
rect 217948 361662 220603 361664
rect 154573 361659 154639 361662
rect 220537 361659 220603 361662
rect 154941 361450 155007 361453
rect 154941 361448 158148 361450
rect 154941 361392 154946 361448
rect 155002 361392 158148 361448
rect 154941 361390 158148 361392
rect 154941 361387 155007 361390
rect 220721 361314 220787 361317
rect 217948 361312 220787 361314
rect 217948 361256 220726 361312
rect 220782 361256 220787 361312
rect 217948 361254 220787 361256
rect 220721 361251 220787 361254
rect 154573 361178 154639 361181
rect 154573 361176 158148 361178
rect 154573 361120 154578 361176
rect 154634 361120 158148 361176
rect 154573 361118 158148 361120
rect 154573 361115 154639 361118
rect 154849 360906 154915 360909
rect 220445 360906 220511 360909
rect 154849 360904 158148 360906
rect 154849 360848 154854 360904
rect 154910 360848 158148 360904
rect 154849 360846 158148 360848
rect 217948 360904 220511 360906
rect 217948 360848 220450 360904
rect 220506 360848 220511 360904
rect 217948 360846 220511 360848
rect 154849 360843 154915 360846
rect 220445 360843 220511 360846
rect 154757 360634 154823 360637
rect 154757 360632 158148 360634
rect 154757 360576 154762 360632
rect 154818 360576 158148 360632
rect 154757 360574 158148 360576
rect 154757 360571 154823 360574
rect 219893 360498 219959 360501
rect 217948 360496 219959 360498
rect 217948 360440 219898 360496
rect 219954 360440 219959 360496
rect 217948 360438 219959 360440
rect 219893 360435 219959 360438
rect 155033 360362 155099 360365
rect 155033 360360 158148 360362
rect 155033 360304 155038 360360
rect 155094 360304 158148 360360
rect 155033 360302 158148 360304
rect 155033 360299 155099 360302
rect 154941 360090 155007 360093
rect 220629 360090 220695 360093
rect 154941 360088 158148 360090
rect 154941 360032 154946 360088
rect 155002 360032 158148 360088
rect 154941 360030 158148 360032
rect 217948 360088 220695 360090
rect 217948 360032 220634 360088
rect 220690 360032 220695 360088
rect 217948 360030 220695 360032
rect 154941 360027 155007 360030
rect 220629 360027 220695 360030
rect 155033 359818 155099 359821
rect 155033 359816 158148 359818
rect 155033 359760 155038 359816
rect 155094 359760 158148 359816
rect 155033 359758 158148 359760
rect 155033 359755 155099 359758
rect 220721 359682 220787 359685
rect 217948 359680 220787 359682
rect 217948 359624 220726 359680
rect 220782 359624 220787 359680
rect 217948 359622 220787 359624
rect 220721 359619 220787 359622
rect 154573 359546 154639 359549
rect 154573 359544 158148 359546
rect 154573 359488 154578 359544
rect 154634 359488 158148 359544
rect 154573 359486 158148 359488
rect 154573 359483 154639 359486
rect 154849 359274 154915 359277
rect 220721 359274 220787 359277
rect 154849 359272 158148 359274
rect 154849 359216 154854 359272
rect 154910 359216 158148 359272
rect 154849 359214 158148 359216
rect 217948 359272 220787 359274
rect 217948 359216 220726 359272
rect 220782 359216 220787 359272
rect 217948 359214 220787 359216
rect 154849 359211 154915 359214
rect 220721 359211 220787 359214
rect 154941 359002 155007 359005
rect 154941 359000 158148 359002
rect 154941 358944 154946 359000
rect 155002 358944 158148 359000
rect 154941 358942 158148 358944
rect 154941 358939 155007 358942
rect 219709 358866 219775 358869
rect 217948 358864 219775 358866
rect 217948 358808 219714 358864
rect 219770 358808 219775 358864
rect 217948 358806 219775 358808
rect 219709 358803 219775 358806
rect 154573 358730 154639 358733
rect 154573 358728 158148 358730
rect 154573 358672 154578 358728
rect 154634 358672 158148 358728
rect 154573 358670 158148 358672
rect 154573 358667 154639 358670
rect -960 358458 480 358548
rect 2957 358458 3023 358461
rect -960 358456 3023 358458
rect -960 358400 2962 358456
rect 3018 358400 3023 358456
rect -960 358398 3023 358400
rect -960 358308 480 358398
rect 2957 358395 3023 358398
rect 155125 358458 155191 358461
rect 219433 358458 219499 358461
rect 155125 358456 158148 358458
rect 155125 358400 155130 358456
rect 155186 358400 158148 358456
rect 155125 358398 158148 358400
rect 217948 358456 219499 358458
rect 217948 358400 219438 358456
rect 219494 358400 219499 358456
rect 217948 358398 219499 358400
rect 155125 358395 155191 358398
rect 219433 358395 219499 358398
rect 155585 358186 155651 358189
rect 155585 358184 158148 358186
rect 155585 358128 155590 358184
rect 155646 358128 158148 358184
rect 155585 358126 158148 358128
rect 155585 358123 155651 358126
rect 220629 358050 220695 358053
rect 217948 358048 220695 358050
rect 217948 357992 220634 358048
rect 220690 357992 220695 358048
rect 217948 357990 220695 357992
rect 220629 357987 220695 357990
rect 154941 357914 155007 357917
rect 154941 357912 158148 357914
rect 154941 357856 154946 357912
rect 155002 357856 158148 357912
rect 154941 357854 158148 357856
rect 154941 357851 155007 357854
rect 154757 357642 154823 357645
rect 219985 357642 220051 357645
rect 154757 357640 158148 357642
rect 154757 357584 154762 357640
rect 154818 357584 158148 357640
rect 154757 357582 158148 357584
rect 217948 357640 220051 357642
rect 217948 357584 219990 357640
rect 220046 357584 220051 357640
rect 217948 357582 220051 357584
rect 154757 357579 154823 357582
rect 219985 357579 220051 357582
rect 154941 357370 155007 357373
rect 154941 357368 158148 357370
rect 154941 357312 154946 357368
rect 155002 357312 158148 357368
rect 154941 357310 158148 357312
rect 154941 357307 155007 357310
rect 220629 357234 220695 357237
rect 217948 357232 220695 357234
rect 217948 357176 220634 357232
rect 220690 357176 220695 357232
rect 217948 357174 220695 357176
rect 220629 357171 220695 357174
rect 155033 357098 155099 357101
rect 155033 357096 158148 357098
rect 155033 357040 155038 357096
rect 155094 357040 158148 357096
rect 155033 357038 158148 357040
rect 155033 357035 155099 357038
rect 154941 356826 155007 356829
rect 219893 356826 219959 356829
rect 154941 356824 158148 356826
rect 154941 356768 154946 356824
rect 155002 356768 158148 356824
rect 154941 356766 158148 356768
rect 217948 356824 219959 356826
rect 217948 356768 219898 356824
rect 219954 356768 219959 356824
rect 217948 356766 219959 356768
rect 154941 356763 155007 356766
rect 219893 356763 219959 356766
rect 154849 356554 154915 356557
rect 154849 356552 158148 356554
rect 154849 356496 154854 356552
rect 154910 356496 158148 356552
rect 154849 356494 158148 356496
rect 154849 356491 154915 356494
rect 220721 356418 220787 356421
rect 217948 356416 220787 356418
rect 217948 356360 220726 356416
rect 220782 356360 220787 356416
rect 217948 356358 220787 356360
rect 220721 356355 220787 356358
rect 154757 356282 154823 356285
rect 154757 356280 158148 356282
rect 154757 356224 154762 356280
rect 154818 356224 158148 356280
rect 154757 356222 158148 356224
rect 154757 356219 154823 356222
rect 154573 356010 154639 356013
rect 220721 356010 220787 356013
rect 154573 356008 158148 356010
rect 154573 355952 154578 356008
rect 154634 355952 158148 356008
rect 154573 355950 158148 355952
rect 217948 356008 220787 356010
rect 217948 355952 220726 356008
rect 220782 355952 220787 356008
rect 217948 355950 220787 355952
rect 154573 355947 154639 355950
rect 220721 355947 220787 355950
rect 154941 355738 155007 355741
rect 154941 355736 158148 355738
rect 154941 355680 154946 355736
rect 155002 355680 158148 355736
rect 154941 355678 158148 355680
rect 154941 355675 155007 355678
rect 220721 355602 220787 355605
rect 217948 355600 220787 355602
rect 217948 355544 220726 355600
rect 220782 355544 220787 355600
rect 217948 355542 220787 355544
rect 220721 355539 220787 355542
rect 154849 355466 154915 355469
rect 154849 355464 158148 355466
rect 154849 355408 154854 355464
rect 154910 355408 158148 355464
rect 154849 355406 158148 355408
rect 154849 355403 154915 355406
rect 155033 355194 155099 355197
rect 220537 355194 220603 355197
rect 155033 355192 158148 355194
rect 155033 355136 155038 355192
rect 155094 355136 158148 355192
rect 155033 355134 158148 355136
rect 217948 355192 220603 355194
rect 217948 355136 220542 355192
rect 220598 355136 220603 355192
rect 217948 355134 220603 355136
rect 155033 355131 155099 355134
rect 220537 355131 220603 355134
rect 155309 354922 155375 354925
rect 155309 354920 158148 354922
rect 155309 354864 155314 354920
rect 155370 354864 158148 354920
rect 155309 354862 158148 354864
rect 155309 354859 155375 354862
rect 219801 354786 219867 354789
rect 217948 354784 219867 354786
rect 217948 354728 219806 354784
rect 219862 354728 219867 354784
rect 217948 354726 219867 354728
rect 219801 354723 219867 354726
rect 154573 354650 154639 354653
rect 154573 354648 158148 354650
rect 154573 354592 154578 354648
rect 154634 354592 158148 354648
rect 154573 354590 158148 354592
rect 154573 354587 154639 354590
rect 154941 354378 155007 354381
rect 220629 354378 220695 354381
rect 154941 354376 158148 354378
rect 154941 354320 154946 354376
rect 155002 354320 158148 354376
rect 154941 354318 158148 354320
rect 217948 354376 220695 354378
rect 217948 354320 220634 354376
rect 220690 354320 220695 354376
rect 217948 354318 220695 354320
rect 154941 354315 155007 354318
rect 220629 354315 220695 354318
rect 154757 354106 154823 354109
rect 154757 354104 158148 354106
rect 154757 354048 154762 354104
rect 154818 354048 158148 354104
rect 154757 354046 158148 354048
rect 154757 354043 154823 354046
rect 220721 353970 220787 353973
rect 217948 353968 220787 353970
rect 217948 353912 220726 353968
rect 220782 353912 220787 353968
rect 217948 353910 220787 353912
rect 220721 353907 220787 353910
rect 155585 353834 155651 353837
rect 155585 353832 158148 353834
rect 155585 353776 155590 353832
rect 155646 353776 158148 353832
rect 155585 353774 158148 353776
rect 155585 353771 155651 353774
rect 154849 353562 154915 353565
rect 220537 353562 220603 353565
rect 154849 353560 158148 353562
rect 154849 353504 154854 353560
rect 154910 353504 158148 353560
rect 154849 353502 158148 353504
rect 217948 353560 220603 353562
rect 217948 353504 220542 353560
rect 220598 353504 220603 353560
rect 217948 353502 220603 353504
rect 154849 353499 154915 353502
rect 220537 353499 220603 353502
rect 154849 353290 154915 353293
rect 154849 353288 158148 353290
rect 154849 353232 154854 353288
rect 154910 353232 158148 353288
rect 154849 353230 158148 353232
rect 154849 353227 154915 353230
rect 220721 353154 220787 353157
rect 217948 353152 220787 353154
rect 217948 353096 220726 353152
rect 220782 353096 220787 353152
rect 217948 353094 220787 353096
rect 220721 353091 220787 353094
rect 154941 353018 155007 353021
rect 154941 353016 158148 353018
rect 154941 352960 154946 353016
rect 155002 352960 158148 353016
rect 154941 352958 158148 352960
rect 154941 352955 155007 352958
rect 155033 352746 155099 352749
rect 220445 352746 220511 352749
rect 155033 352744 158148 352746
rect 155033 352688 155038 352744
rect 155094 352688 158148 352744
rect 155033 352686 158148 352688
rect 217948 352744 220511 352746
rect 217948 352688 220450 352744
rect 220506 352688 220511 352744
rect 217948 352686 220511 352688
rect 155033 352683 155099 352686
rect 220445 352683 220511 352686
rect 154757 352474 154823 352477
rect 154757 352472 158148 352474
rect 154757 352416 154762 352472
rect 154818 352416 158148 352472
rect 154757 352414 158148 352416
rect 154757 352411 154823 352414
rect 220445 352338 220511 352341
rect 217948 352336 220511 352338
rect 217948 352280 220450 352336
rect 220506 352280 220511 352336
rect 217948 352278 220511 352280
rect 220445 352275 220511 352278
rect 154849 352202 154915 352205
rect 154849 352200 158148 352202
rect 154849 352144 154854 352200
rect 154910 352144 158148 352200
rect 154849 352142 158148 352144
rect 154849 352139 154915 352142
rect 155401 351930 155467 351933
rect 219893 351930 219959 351933
rect 155401 351928 158148 351930
rect 155401 351872 155406 351928
rect 155462 351872 158148 351928
rect 155401 351870 158148 351872
rect 217948 351928 219959 351930
rect 217948 351872 219898 351928
rect 219954 351872 219959 351928
rect 217948 351870 219959 351872
rect 155401 351867 155467 351870
rect 219893 351867 219959 351870
rect 580165 351930 580231 351933
rect 583520 351930 584960 352020
rect 580165 351928 584960 351930
rect 580165 351872 580170 351928
rect 580226 351872 584960 351928
rect 580165 351870 584960 351872
rect 580165 351867 580231 351870
rect 583520 351780 584960 351870
rect 154941 351658 155007 351661
rect 154941 351656 158148 351658
rect 154941 351600 154946 351656
rect 155002 351600 158148 351656
rect 154941 351598 158148 351600
rect 154941 351595 155007 351598
rect 220721 351522 220787 351525
rect 217948 351520 220787 351522
rect 217948 351464 220726 351520
rect 220782 351464 220787 351520
rect 217948 351462 220787 351464
rect 220721 351459 220787 351462
rect 154757 351386 154823 351389
rect 154757 351384 158148 351386
rect 154757 351328 154762 351384
rect 154818 351328 158148 351384
rect 154757 351326 158148 351328
rect 154757 351323 154823 351326
rect 154849 351114 154915 351117
rect 219985 351114 220051 351117
rect 154849 351112 158148 351114
rect 154849 351056 154854 351112
rect 154910 351056 158148 351112
rect 154849 351054 158148 351056
rect 217948 351112 220051 351114
rect 217948 351056 219990 351112
rect 220046 351056 220051 351112
rect 217948 351054 220051 351056
rect 154849 351051 154915 351054
rect 219985 351051 220051 351054
rect 155125 350842 155191 350845
rect 155125 350840 158148 350842
rect 155125 350784 155130 350840
rect 155186 350784 158148 350840
rect 155125 350782 158148 350784
rect 155125 350779 155191 350782
rect 219893 350706 219959 350709
rect 217948 350704 219959 350706
rect 217948 350648 219898 350704
rect 219954 350648 219959 350704
rect 217948 350646 219959 350648
rect 219893 350643 219959 350646
rect 155033 350570 155099 350573
rect 155033 350568 158148 350570
rect 155033 350512 155038 350568
rect 155094 350512 158148 350568
rect 155033 350510 158148 350512
rect 155033 350507 155099 350510
rect 154573 350298 154639 350301
rect 220353 350298 220419 350301
rect 154573 350296 158148 350298
rect 154573 350240 154578 350296
rect 154634 350240 158148 350296
rect 154573 350238 158148 350240
rect 217948 350296 220419 350298
rect 217948 350240 220358 350296
rect 220414 350240 220419 350296
rect 217948 350238 220419 350240
rect 154573 350235 154639 350238
rect 220353 350235 220419 350238
rect 154941 350026 155007 350029
rect 154941 350024 158148 350026
rect 154941 349968 154946 350024
rect 155002 349968 158148 350024
rect 154941 349966 158148 349968
rect 154941 349963 155007 349966
rect 220537 349890 220603 349893
rect 217948 349888 220603 349890
rect 217948 349832 220542 349888
rect 220598 349832 220603 349888
rect 217948 349830 220603 349832
rect 220537 349827 220603 349830
rect 154941 349754 155007 349757
rect 154941 349752 158148 349754
rect 154941 349696 154946 349752
rect 155002 349696 158148 349752
rect 154941 349694 158148 349696
rect 154941 349691 155007 349694
rect 154849 349482 154915 349485
rect 219893 349482 219959 349485
rect 154849 349480 158148 349482
rect 154849 349424 154854 349480
rect 154910 349424 158148 349480
rect 154849 349422 158148 349424
rect 217948 349480 219959 349482
rect 217948 349424 219898 349480
rect 219954 349424 219959 349480
rect 217948 349422 219959 349424
rect 154849 349419 154915 349422
rect 219893 349419 219959 349422
rect 155493 349210 155559 349213
rect 155493 349208 158148 349210
rect 155493 349152 155498 349208
rect 155554 349152 158148 349208
rect 155493 349150 158148 349152
rect 155493 349147 155559 349150
rect 220537 349074 220603 349077
rect 217948 349072 220603 349074
rect 217948 349016 220542 349072
rect 220598 349016 220603 349072
rect 217948 349014 220603 349016
rect 220537 349011 220603 349014
rect 155033 348938 155099 348941
rect 155033 348936 158148 348938
rect 155033 348880 155038 348936
rect 155094 348880 158148 348936
rect 155033 348878 158148 348880
rect 155033 348875 155099 348878
rect 154849 348666 154915 348669
rect 220721 348666 220787 348669
rect 154849 348664 158148 348666
rect 154849 348608 154854 348664
rect 154910 348608 158148 348664
rect 154849 348606 158148 348608
rect 217948 348664 220787 348666
rect 217948 348608 220726 348664
rect 220782 348608 220787 348664
rect 217948 348606 220787 348608
rect 154849 348603 154915 348606
rect 220721 348603 220787 348606
rect 154757 348394 154823 348397
rect 154757 348392 158148 348394
rect 154757 348336 154762 348392
rect 154818 348336 158148 348392
rect 154757 348334 158148 348336
rect 154757 348331 154823 348334
rect 220629 348258 220695 348261
rect 217948 348256 220695 348258
rect 217948 348200 220634 348256
rect 220690 348200 220695 348256
rect 217948 348198 220695 348200
rect 220629 348195 220695 348198
rect 154941 348122 155007 348125
rect 154941 348120 158148 348122
rect 154941 348064 154946 348120
rect 155002 348064 158148 348120
rect 154941 348062 158148 348064
rect 154941 348059 155007 348062
rect 154941 347850 155007 347853
rect 220445 347850 220511 347853
rect 154941 347848 158148 347850
rect 154941 347792 154946 347848
rect 155002 347792 158148 347848
rect 154941 347790 158148 347792
rect 217948 347848 220511 347850
rect 217948 347792 220450 347848
rect 220506 347792 220511 347848
rect 217948 347790 220511 347792
rect 154941 347787 155007 347790
rect 220445 347787 220511 347790
rect 155033 347578 155099 347581
rect 155033 347576 158148 347578
rect 155033 347520 155038 347576
rect 155094 347520 158148 347576
rect 155033 347518 158148 347520
rect 155033 347515 155099 347518
rect 220721 347442 220787 347445
rect 217948 347440 220787 347442
rect 217948 347384 220726 347440
rect 220782 347384 220787 347440
rect 217948 347382 220787 347384
rect 220721 347379 220787 347382
rect 154849 347306 154915 347309
rect 154849 347304 158148 347306
rect 154849 347248 154854 347304
rect 154910 347248 158148 347304
rect 154849 347246 158148 347248
rect 154849 347243 154915 347246
rect 154573 347034 154639 347037
rect 220445 347034 220511 347037
rect 154573 347032 158148 347034
rect 154573 346976 154578 347032
rect 154634 346976 158148 347032
rect 154573 346974 158148 346976
rect 217948 347032 220511 347034
rect 217948 346976 220450 347032
rect 220506 346976 220511 347032
rect 217948 346974 220511 346976
rect 154573 346971 154639 346974
rect 220445 346971 220511 346974
rect 154941 346762 155007 346765
rect 154941 346760 158148 346762
rect 154941 346704 154946 346760
rect 155002 346704 158148 346760
rect 154941 346702 158148 346704
rect 154941 346699 155007 346702
rect 220629 346626 220695 346629
rect 217948 346624 220695 346626
rect 217948 346568 220634 346624
rect 220690 346568 220695 346624
rect 217948 346566 220695 346568
rect 220629 346563 220695 346566
rect 154849 346490 154915 346493
rect 154849 346488 158148 346490
rect 154849 346432 154854 346488
rect 154910 346432 158148 346488
rect 154849 346430 158148 346432
rect 154849 346427 154915 346430
rect 155033 346218 155099 346221
rect 220721 346218 220787 346221
rect 155033 346216 158148 346218
rect 155033 346160 155038 346216
rect 155094 346160 158148 346216
rect 155033 346158 158148 346160
rect 217948 346216 220787 346218
rect 217948 346160 220726 346216
rect 220782 346160 220787 346216
rect 217948 346158 220787 346160
rect 155033 346155 155099 346158
rect 220721 346155 220787 346158
rect 154941 345946 155007 345949
rect 154941 345944 158148 345946
rect 154941 345888 154946 345944
rect 155002 345888 158148 345944
rect 154941 345886 158148 345888
rect 154941 345883 155007 345886
rect 220721 345810 220787 345813
rect 217948 345808 220787 345810
rect 217948 345752 220726 345808
rect 220782 345752 220787 345808
rect 217948 345750 220787 345752
rect 220721 345747 220787 345750
rect 154990 345614 158148 345674
rect 154849 345538 154915 345541
rect 154990 345538 155050 345614
rect 154849 345536 155050 345538
rect -960 345402 480 345492
rect 154849 345480 154854 345536
rect 154910 345480 155050 345536
rect 154849 345478 155050 345480
rect 154849 345475 154915 345478
rect 3049 345402 3115 345405
rect -960 345400 3115 345402
rect -960 345344 3054 345400
rect 3110 345344 3115 345400
rect -960 345342 3115 345344
rect -960 345252 480 345342
rect 3049 345339 3115 345342
rect 155585 345402 155651 345405
rect 220629 345402 220695 345405
rect 155585 345400 158148 345402
rect 155585 345344 155590 345400
rect 155646 345344 158148 345400
rect 155585 345342 158148 345344
rect 217948 345400 220695 345402
rect 217948 345344 220634 345400
rect 220690 345344 220695 345400
rect 217948 345342 220695 345344
rect 155585 345339 155651 345342
rect 220629 345339 220695 345342
rect 154941 345130 155007 345133
rect 154941 345128 158148 345130
rect 154941 345072 154946 345128
rect 155002 345072 158148 345128
rect 154941 345070 158148 345072
rect 154941 345067 155007 345070
rect 220353 344994 220419 344997
rect 217948 344992 220419 344994
rect 217948 344936 220358 344992
rect 220414 344936 220419 344992
rect 217948 344934 220419 344936
rect 220353 344931 220419 344934
rect 155033 344858 155099 344861
rect 155033 344856 158148 344858
rect 155033 344800 155038 344856
rect 155094 344800 158148 344856
rect 155033 344798 158148 344800
rect 155033 344795 155099 344798
rect 154941 344586 155007 344589
rect 220721 344586 220787 344589
rect 154941 344584 158148 344586
rect 154941 344528 154946 344584
rect 155002 344528 158148 344584
rect 154941 344526 158148 344528
rect 217948 344584 220787 344586
rect 217948 344528 220726 344584
rect 220782 344528 220787 344584
rect 217948 344526 220787 344528
rect 154941 344523 155007 344526
rect 220721 344523 220787 344526
rect 154849 344314 154915 344317
rect 154849 344312 158148 344314
rect 154849 344256 154854 344312
rect 154910 344256 158148 344312
rect 154849 344254 158148 344256
rect 154849 344251 154915 344254
rect 220629 344178 220695 344181
rect 217948 344176 220695 344178
rect 217948 344120 220634 344176
rect 220690 344120 220695 344176
rect 217948 344118 220695 344120
rect 220629 344115 220695 344118
rect 154573 344042 154639 344045
rect 154573 344040 158148 344042
rect 154573 343984 154578 344040
rect 154634 343984 158148 344040
rect 154573 343982 158148 343984
rect 154573 343979 154639 343982
rect 154573 343770 154639 343773
rect 219893 343770 219959 343773
rect 154573 343768 158148 343770
rect 154573 343712 154578 343768
rect 154634 343712 158148 343768
rect 154573 343710 158148 343712
rect 217948 343768 219959 343770
rect 217948 343712 219898 343768
rect 219954 343712 219959 343768
rect 217948 343710 219959 343712
rect 154573 343707 154639 343710
rect 219893 343707 219959 343710
rect 155033 343498 155099 343501
rect 155033 343496 158148 343498
rect 155033 343440 155038 343496
rect 155094 343440 158148 343496
rect 155033 343438 158148 343440
rect 155033 343435 155099 343438
rect 220629 343362 220695 343365
rect 217948 343360 220695 343362
rect 217948 343304 220634 343360
rect 220690 343304 220695 343360
rect 217948 343302 220695 343304
rect 220629 343299 220695 343302
rect 155493 343226 155559 343229
rect 155493 343224 158148 343226
rect 155493 343168 155498 343224
rect 155554 343168 158148 343224
rect 155493 343166 158148 343168
rect 155493 343163 155559 343166
rect 154849 342954 154915 342957
rect 220721 342954 220787 342957
rect 154849 342952 158148 342954
rect 154849 342896 154854 342952
rect 154910 342896 158148 342952
rect 154849 342894 158148 342896
rect 217948 342952 220787 342954
rect 217948 342896 220726 342952
rect 220782 342896 220787 342952
rect 217948 342894 220787 342896
rect 154849 342891 154915 342894
rect 220721 342891 220787 342894
rect 155677 342682 155743 342685
rect 155677 342680 158148 342682
rect 155677 342624 155682 342680
rect 155738 342624 158148 342680
rect 155677 342622 158148 342624
rect 155677 342619 155743 342622
rect 220445 342546 220511 342549
rect 217948 342544 220511 342546
rect 217948 342488 220450 342544
rect 220506 342488 220511 342544
rect 217948 342486 220511 342488
rect 220445 342483 220511 342486
rect 154941 342410 155007 342413
rect 154941 342408 158148 342410
rect 154941 342352 154946 342408
rect 155002 342352 158148 342408
rect 154941 342350 158148 342352
rect 154941 342347 155007 342350
rect 154757 342138 154823 342141
rect 220721 342138 220787 342141
rect 154757 342136 158148 342138
rect 154757 342080 154762 342136
rect 154818 342080 158148 342136
rect 154757 342078 158148 342080
rect 217948 342136 220787 342138
rect 217948 342080 220726 342136
rect 220782 342080 220787 342136
rect 217948 342078 220787 342080
rect 154757 342075 154823 342078
rect 220721 342075 220787 342078
rect 154941 341866 155007 341869
rect 154941 341864 158148 341866
rect 154941 341808 154946 341864
rect 155002 341808 158148 341864
rect 154941 341806 158148 341808
rect 154941 341803 155007 341806
rect 219801 341730 219867 341733
rect 217948 341728 219867 341730
rect 217948 341672 219806 341728
rect 219862 341672 219867 341728
rect 217948 341670 219867 341672
rect 219801 341667 219867 341670
rect 155033 341594 155099 341597
rect 155033 341592 158148 341594
rect 155033 341536 155038 341592
rect 155094 341536 158148 341592
rect 155033 341534 158148 341536
rect 155033 341531 155099 341534
rect 154849 341322 154915 341325
rect 220537 341322 220603 341325
rect 154849 341320 158148 341322
rect 154849 341264 154854 341320
rect 154910 341264 158148 341320
rect 154849 341262 158148 341264
rect 217948 341320 220603 341322
rect 217948 341264 220542 341320
rect 220598 341264 220603 341320
rect 217948 341262 220603 341264
rect 154849 341259 154915 341262
rect 220537 341259 220603 341262
rect 155125 341050 155191 341053
rect 155125 341048 158148 341050
rect 155125 340992 155130 341048
rect 155186 340992 158148 341048
rect 155125 340990 158148 340992
rect 155125 340987 155191 340990
rect 220261 340914 220327 340917
rect 217948 340912 220327 340914
rect 217948 340856 220266 340912
rect 220322 340856 220327 340912
rect 217948 340854 220327 340856
rect 220261 340851 220327 340854
rect 155033 340778 155099 340781
rect 155033 340776 158148 340778
rect 155033 340720 155038 340776
rect 155094 340720 158148 340776
rect 155033 340718 158148 340720
rect 155033 340715 155099 340718
rect 154757 340506 154823 340509
rect 219893 340506 219959 340509
rect 154757 340504 158148 340506
rect 154757 340448 154762 340504
rect 154818 340448 158148 340504
rect 154757 340446 158148 340448
rect 217948 340504 219959 340506
rect 217948 340448 219898 340504
rect 219954 340448 219959 340504
rect 217948 340446 219959 340448
rect 154757 340443 154823 340446
rect 219893 340443 219959 340446
rect 154941 340234 155007 340237
rect 154941 340232 158148 340234
rect 154941 340176 154946 340232
rect 155002 340176 158148 340232
rect 154941 340174 158148 340176
rect 154941 340171 155007 340174
rect 220169 340098 220235 340101
rect 217948 340096 220235 340098
rect 217948 340040 220174 340096
rect 220230 340040 220235 340096
rect 217948 340038 220235 340040
rect 220169 340035 220235 340038
rect 154849 339962 154915 339965
rect 154849 339960 158148 339962
rect 154849 339904 154854 339960
rect 154910 339904 158148 339960
rect 154849 339902 158148 339904
rect 154849 339899 154915 339902
rect 154941 339690 155007 339693
rect 219525 339690 219591 339693
rect 154941 339688 158148 339690
rect 154941 339632 154946 339688
rect 155002 339632 158148 339688
rect 154941 339630 158148 339632
rect 217948 339688 219591 339690
rect 217948 339632 219530 339688
rect 219586 339632 219591 339688
rect 217948 339630 219591 339632
rect 154941 339627 155007 339630
rect 219525 339627 219591 339630
rect 154665 339418 154731 339421
rect 154665 339416 158148 339418
rect 154665 339360 154670 339416
rect 154726 339360 158148 339416
rect 154665 339358 158148 339360
rect 154665 339355 154731 339358
rect 220721 339282 220787 339285
rect 217948 339280 220787 339282
rect 217948 339224 220726 339280
rect 220782 339224 220787 339280
rect 217948 339222 220787 339224
rect 220721 339219 220787 339222
rect 154849 339146 154915 339149
rect 154849 339144 158148 339146
rect 154849 339088 154854 339144
rect 154910 339088 158148 339144
rect 154849 339086 158148 339088
rect 154849 339083 154915 339086
rect 155033 338874 155099 338877
rect 220629 338874 220695 338877
rect 155033 338872 158148 338874
rect 155033 338816 155038 338872
rect 155094 338816 158148 338872
rect 155033 338814 158148 338816
rect 217948 338872 220695 338874
rect 217948 338816 220634 338872
rect 220690 338816 220695 338872
rect 217948 338814 220695 338816
rect 155033 338811 155099 338814
rect 220629 338811 220695 338814
rect 154941 338602 155007 338605
rect 154941 338600 158148 338602
rect 154941 338544 154946 338600
rect 155002 338544 158148 338600
rect 154941 338542 158148 338544
rect 154941 338539 155007 338542
rect 220445 338466 220511 338469
rect 217948 338464 220511 338466
rect 217948 338408 220450 338464
rect 220506 338408 220511 338464
rect 583520 338452 584960 338692
rect 217948 338406 220511 338408
rect 220445 338403 220511 338406
rect 155217 338330 155283 338333
rect 155217 338328 158148 338330
rect 155217 338272 155222 338328
rect 155278 338272 158148 338328
rect 155217 338270 158148 338272
rect 155217 338267 155283 338270
rect 154757 338058 154823 338061
rect 219893 338058 219959 338061
rect 154757 338056 158148 338058
rect 154757 338000 154762 338056
rect 154818 338000 158148 338056
rect 154757 337998 158148 338000
rect 217948 338056 219959 338058
rect 217948 338000 219898 338056
rect 219954 338000 219959 338056
rect 217948 337998 219959 338000
rect 154757 337995 154823 337998
rect 219893 337995 219959 337998
rect 154849 337786 154915 337789
rect 154849 337784 158148 337786
rect 154849 337728 154854 337784
rect 154910 337728 158148 337784
rect 154849 337726 158148 337728
rect 154849 337723 154915 337726
rect 220629 337650 220695 337653
rect 217948 337648 220695 337650
rect 217948 337592 220634 337648
rect 220690 337592 220695 337648
rect 217948 337590 220695 337592
rect 220629 337587 220695 337590
rect 155033 337514 155099 337517
rect 155033 337512 158148 337514
rect 155033 337456 155038 337512
rect 155094 337456 158148 337512
rect 155033 337454 158148 337456
rect 155033 337451 155099 337454
rect 154573 337242 154639 337245
rect 220721 337242 220787 337245
rect 154573 337240 158148 337242
rect 154573 337184 154578 337240
rect 154634 337184 158148 337240
rect 154573 337182 158148 337184
rect 217948 337240 220787 337242
rect 217948 337184 220726 337240
rect 220782 337184 220787 337240
rect 217948 337182 220787 337184
rect 154573 337179 154639 337182
rect 220721 337179 220787 337182
rect 154941 336970 155007 336973
rect 154941 336968 158148 336970
rect 154941 336912 154946 336968
rect 155002 336912 158148 336968
rect 154941 336910 158148 336912
rect 154941 336907 155007 336910
rect 220537 336834 220603 336837
rect 217948 336832 220603 336834
rect 217948 336776 220542 336832
rect 220598 336776 220603 336832
rect 217948 336774 220603 336776
rect 220537 336771 220603 336774
rect 154757 336698 154823 336701
rect 154757 336696 158148 336698
rect 154757 336640 154762 336696
rect 154818 336640 158148 336696
rect 154757 336638 158148 336640
rect 154757 336635 154823 336638
rect 154665 336426 154731 336429
rect 220629 336426 220695 336429
rect 154665 336424 158148 336426
rect 154665 336368 154670 336424
rect 154726 336368 158148 336424
rect 154665 336366 158148 336368
rect 217948 336424 220695 336426
rect 217948 336368 220634 336424
rect 220690 336368 220695 336424
rect 217948 336366 220695 336368
rect 154665 336363 154731 336366
rect 220629 336363 220695 336366
rect 155033 336154 155099 336157
rect 155033 336152 158148 336154
rect 155033 336096 155038 336152
rect 155094 336096 158148 336152
rect 155033 336094 158148 336096
rect 155033 336091 155099 336094
rect 220537 336018 220603 336021
rect 217948 336016 220603 336018
rect 217948 335960 220542 336016
rect 220598 335960 220603 336016
rect 217948 335958 220603 335960
rect 220537 335955 220603 335958
rect 154849 335882 154915 335885
rect 154849 335880 158148 335882
rect 154849 335824 154854 335880
rect 154910 335824 158148 335880
rect 154849 335822 158148 335824
rect 154849 335819 154915 335822
rect 154941 335610 155007 335613
rect 220721 335610 220787 335613
rect 154941 335608 158148 335610
rect 154941 335552 154946 335608
rect 155002 335552 158148 335608
rect 154941 335550 158148 335552
rect 217948 335608 220787 335610
rect 217948 335552 220726 335608
rect 220782 335552 220787 335608
rect 217948 335550 220787 335552
rect 154941 335547 155007 335550
rect 220721 335547 220787 335550
rect 155585 335338 155651 335341
rect 155585 335336 158148 335338
rect 155585 335280 155590 335336
rect 155646 335280 158148 335336
rect 155585 335278 158148 335280
rect 155585 335275 155651 335278
rect 220169 335202 220235 335205
rect 217948 335200 220235 335202
rect 217948 335144 220174 335200
rect 220230 335144 220235 335200
rect 217948 335142 220235 335144
rect 220169 335139 220235 335142
rect 155861 335066 155927 335069
rect 155861 335064 158148 335066
rect 155861 335008 155866 335064
rect 155922 335008 158148 335064
rect 155861 335006 158148 335008
rect 155861 335003 155927 335006
rect 154757 334794 154823 334797
rect 219985 334794 220051 334797
rect 154757 334792 158148 334794
rect 154757 334736 154762 334792
rect 154818 334736 158148 334792
rect 154757 334734 158148 334736
rect 217948 334792 220051 334794
rect 217948 334736 219990 334792
rect 220046 334736 220051 334792
rect 217948 334734 220051 334736
rect 154757 334731 154823 334734
rect 219985 334731 220051 334734
rect 155125 334522 155191 334525
rect 155125 334520 158148 334522
rect 155125 334464 155130 334520
rect 155186 334464 158148 334520
rect 155125 334462 158148 334464
rect 155125 334459 155191 334462
rect 220353 334386 220419 334389
rect 217948 334384 220419 334386
rect 217948 334328 220358 334384
rect 220414 334328 220419 334384
rect 217948 334326 220419 334328
rect 220353 334323 220419 334326
rect 154941 334250 155007 334253
rect 154941 334248 158148 334250
rect 154941 334192 154946 334248
rect 155002 334192 158148 334248
rect 154941 334190 158148 334192
rect 154941 334187 155007 334190
rect 154849 333978 154915 333981
rect 220445 333978 220511 333981
rect 154849 333976 158148 333978
rect 154849 333920 154854 333976
rect 154910 333920 158148 333976
rect 154849 333918 158148 333920
rect 217948 333976 220511 333978
rect 217948 333920 220450 333976
rect 220506 333920 220511 333976
rect 217948 333918 220511 333920
rect 154849 333915 154915 333918
rect 220445 333915 220511 333918
rect 154941 333706 155007 333709
rect 154941 333704 158148 333706
rect 154941 333648 154946 333704
rect 155002 333648 158148 333704
rect 154941 333646 158148 333648
rect 154941 333643 155007 333646
rect 220629 333570 220695 333573
rect 217948 333568 220695 333570
rect 217948 333512 220634 333568
rect 220690 333512 220695 333568
rect 217948 333510 220695 333512
rect 220629 333507 220695 333510
rect 154757 333434 154823 333437
rect 154757 333432 158148 333434
rect 154757 333376 154762 333432
rect 154818 333376 158148 333432
rect 154757 333374 158148 333376
rect 154757 333371 154823 333374
rect 154021 333162 154087 333165
rect 219801 333162 219867 333165
rect 154021 333160 158148 333162
rect 154021 333104 154026 333160
rect 154082 333104 158148 333160
rect 154021 333102 158148 333104
rect 217948 333160 219867 333162
rect 217948 333104 219806 333160
rect 219862 333104 219867 333160
rect 217948 333102 219867 333104
rect 154021 333099 154087 333102
rect 219801 333099 219867 333102
rect 154573 332890 154639 332893
rect 154573 332888 158148 332890
rect 154573 332832 154578 332888
rect 154634 332832 158148 332888
rect 154573 332830 158148 332832
rect 154573 332827 154639 332830
rect 220721 332754 220787 332757
rect 217948 332752 220787 332754
rect 217948 332696 220726 332752
rect 220782 332696 220787 332752
rect 217948 332694 220787 332696
rect 220721 332691 220787 332694
rect 154757 332618 154823 332621
rect 154757 332616 158148 332618
rect 154757 332560 154762 332616
rect 154818 332560 158148 332616
rect 154757 332558 158148 332560
rect 154757 332555 154823 332558
rect -960 332196 480 332436
rect 155769 332346 155835 332349
rect 219893 332346 219959 332349
rect 155769 332344 158148 332346
rect 155769 332288 155774 332344
rect 155830 332288 158148 332344
rect 155769 332286 158148 332288
rect 217948 332344 219959 332346
rect 217948 332288 219898 332344
rect 219954 332288 219959 332344
rect 217948 332286 219959 332288
rect 155769 332283 155835 332286
rect 219893 332283 219959 332286
rect 154941 332074 155007 332077
rect 154941 332072 158148 332074
rect 154941 332016 154946 332072
rect 155002 332016 158148 332072
rect 154941 332014 158148 332016
rect 154941 332011 155007 332014
rect 220537 331938 220603 331941
rect 217948 331936 220603 331938
rect 217948 331880 220542 331936
rect 220598 331880 220603 331936
rect 217948 331878 220603 331880
rect 220537 331875 220603 331878
rect 155033 331802 155099 331805
rect 155033 331800 158148 331802
rect 155033 331744 155038 331800
rect 155094 331744 158148 331800
rect 155033 331742 158148 331744
rect 155033 331739 155099 331742
rect 154849 331530 154915 331533
rect 219893 331530 219959 331533
rect 154849 331528 158148 331530
rect 154849 331472 154854 331528
rect 154910 331472 158148 331528
rect 154849 331470 158148 331472
rect 217948 331528 219959 331530
rect 217948 331472 219898 331528
rect 219954 331472 219959 331528
rect 217948 331470 219959 331472
rect 154849 331467 154915 331470
rect 219893 331467 219959 331470
rect 154941 331258 155007 331261
rect 154941 331256 158148 331258
rect 154941 331200 154946 331256
rect 155002 331200 158148 331256
rect 154941 331198 158148 331200
rect 154941 331195 155007 331198
rect 220537 331122 220603 331125
rect 217948 331120 220603 331122
rect 217948 331064 220542 331120
rect 220598 331064 220603 331120
rect 217948 331062 220603 331064
rect 220537 331059 220603 331062
rect 155033 330986 155099 330989
rect 155033 330984 158148 330986
rect 155033 330928 155038 330984
rect 155094 330928 158148 330984
rect 155033 330926 158148 330928
rect 155033 330923 155099 330926
rect 155125 330714 155191 330717
rect 219709 330714 219775 330717
rect 155125 330712 158148 330714
rect 155125 330656 155130 330712
rect 155186 330656 158148 330712
rect 155125 330654 158148 330656
rect 217948 330712 219775 330714
rect 217948 330656 219714 330712
rect 219770 330656 219775 330712
rect 217948 330654 219775 330656
rect 155125 330651 155191 330654
rect 219709 330651 219775 330654
rect 154849 330442 154915 330445
rect 154849 330440 158148 330442
rect 154849 330384 154854 330440
rect 154910 330384 158148 330440
rect 154849 330382 158148 330384
rect 154849 330379 154915 330382
rect 220721 330306 220787 330309
rect 217948 330304 220787 330306
rect 217948 330248 220726 330304
rect 220782 330248 220787 330304
rect 217948 330246 220787 330248
rect 220721 330243 220787 330246
rect 154941 330170 155007 330173
rect 154941 330168 158148 330170
rect 154941 330112 154946 330168
rect 155002 330112 158148 330168
rect 154941 330110 158148 330112
rect 154941 330107 155007 330110
rect 154573 329898 154639 329901
rect 220629 329898 220695 329901
rect 154573 329896 158148 329898
rect 154573 329840 154578 329896
rect 154634 329840 158148 329896
rect 154573 329838 158148 329840
rect 217948 329896 220695 329898
rect 217948 329840 220634 329896
rect 220690 329840 220695 329896
rect 217948 329838 220695 329840
rect 154573 329835 154639 329838
rect 220629 329835 220695 329838
rect 154849 329626 154915 329629
rect 154849 329624 158148 329626
rect 154849 329568 154854 329624
rect 154910 329568 158148 329624
rect 154849 329566 158148 329568
rect 154849 329563 154915 329566
rect 220537 329490 220603 329493
rect 217948 329488 220603 329490
rect 217948 329432 220542 329488
rect 220598 329432 220603 329488
rect 217948 329430 220603 329432
rect 220537 329427 220603 329430
rect 155125 329354 155191 329357
rect 155125 329352 158148 329354
rect 155125 329296 155130 329352
rect 155186 329296 158148 329352
rect 155125 329294 158148 329296
rect 155125 329291 155191 329294
rect 155033 329082 155099 329085
rect 219525 329082 219591 329085
rect 155033 329080 158148 329082
rect 155033 329024 155038 329080
rect 155094 329024 158148 329080
rect 155033 329022 158148 329024
rect 217948 329080 219591 329082
rect 217948 329024 219530 329080
rect 219586 329024 219591 329080
rect 217948 329022 219591 329024
rect 155033 329019 155099 329022
rect 219525 329019 219591 329022
rect 154941 328810 155007 328813
rect 154941 328808 158148 328810
rect 154941 328752 154946 328808
rect 155002 328752 158148 328808
rect 154941 328750 158148 328752
rect 154941 328747 155007 328750
rect 220721 328674 220787 328677
rect 217948 328672 220787 328674
rect 217948 328616 220726 328672
rect 220782 328616 220787 328672
rect 217948 328614 220787 328616
rect 220721 328611 220787 328614
rect 154573 328538 154639 328541
rect 154573 328536 158148 328538
rect 154573 328480 154578 328536
rect 154634 328480 158148 328536
rect 154573 328478 158148 328480
rect 154573 328475 154639 328478
rect 155033 328266 155099 328269
rect 220261 328266 220327 328269
rect 155033 328264 158148 328266
rect 155033 328208 155038 328264
rect 155094 328208 158148 328264
rect 155033 328206 158148 328208
rect 217948 328264 220327 328266
rect 217948 328208 220266 328264
rect 220322 328208 220327 328264
rect 217948 328206 220327 328208
rect 155033 328203 155099 328206
rect 220261 328203 220327 328206
rect 154665 327994 154731 327997
rect 154665 327992 158148 327994
rect 154665 327936 154670 327992
rect 154726 327936 158148 327992
rect 154665 327934 158148 327936
rect 154665 327931 154731 327934
rect 220261 327858 220327 327861
rect 217948 327856 220327 327858
rect 217948 327800 220266 327856
rect 220322 327800 220327 327856
rect 217948 327798 220327 327800
rect 220261 327795 220327 327798
rect 154849 327722 154915 327725
rect 154849 327720 158148 327722
rect 154849 327664 154854 327720
rect 154910 327664 158148 327720
rect 154849 327662 158148 327664
rect 154849 327659 154915 327662
rect 154941 327450 155007 327453
rect 220721 327450 220787 327453
rect 154941 327448 158148 327450
rect 154941 327392 154946 327448
rect 155002 327392 158148 327448
rect 154941 327390 158148 327392
rect 217948 327448 220787 327450
rect 217948 327392 220726 327448
rect 220782 327392 220787 327448
rect 217948 327390 220787 327392
rect 154941 327387 155007 327390
rect 220721 327387 220787 327390
rect 154757 327178 154823 327181
rect 154757 327176 158148 327178
rect 154757 327120 154762 327176
rect 154818 327120 158148 327176
rect 154757 327118 158148 327120
rect 154757 327115 154823 327118
rect 219525 327042 219591 327045
rect 217948 327040 219591 327042
rect 217948 326984 219530 327040
rect 219586 326984 219591 327040
rect 217948 326982 219591 326984
rect 219525 326979 219591 326982
rect 154849 326906 154915 326909
rect 154849 326904 158148 326906
rect 154849 326848 154854 326904
rect 154910 326848 158148 326904
rect 154849 326846 158148 326848
rect 154849 326843 154915 326846
rect 154941 326634 155007 326637
rect 220629 326634 220695 326637
rect 154941 326632 158148 326634
rect 154941 326576 154946 326632
rect 155002 326576 158148 326632
rect 154941 326574 158148 326576
rect 217948 326632 220695 326634
rect 217948 326576 220634 326632
rect 220690 326576 220695 326632
rect 217948 326574 220695 326576
rect 154941 326571 155007 326574
rect 220629 326571 220695 326574
rect 154757 326362 154823 326365
rect 154757 326360 158148 326362
rect 154757 326304 154762 326360
rect 154818 326304 158148 326360
rect 154757 326302 158148 326304
rect 154757 326299 154823 326302
rect 220353 326226 220419 326229
rect 217948 326224 220419 326226
rect 217948 326168 220358 326224
rect 220414 326168 220419 326224
rect 217948 326166 220419 326168
rect 220353 326163 220419 326166
rect 155033 326090 155099 326093
rect 155033 326088 158148 326090
rect 155033 326032 155038 326088
rect 155094 326032 158148 326088
rect 155033 326030 158148 326032
rect 155033 326027 155099 326030
rect 154573 325818 154639 325821
rect 220721 325818 220787 325821
rect 154573 325816 158148 325818
rect 154573 325760 154578 325816
rect 154634 325760 158148 325816
rect 154573 325758 158148 325760
rect 217948 325816 220787 325818
rect 217948 325760 220726 325816
rect 220782 325760 220787 325816
rect 217948 325758 220787 325760
rect 154573 325755 154639 325758
rect 220721 325755 220787 325758
rect 155033 325546 155099 325549
rect 155033 325544 158148 325546
rect 155033 325488 155038 325544
rect 155094 325488 158148 325544
rect 155033 325486 158148 325488
rect 155033 325483 155099 325486
rect 220261 325410 220327 325413
rect 217948 325408 220327 325410
rect 217948 325352 220266 325408
rect 220322 325352 220327 325408
rect 217948 325350 220327 325352
rect 220261 325347 220327 325350
rect 154757 325274 154823 325277
rect 580165 325274 580231 325277
rect 583520 325274 584960 325364
rect 154757 325272 158148 325274
rect 154757 325216 154762 325272
rect 154818 325216 158148 325272
rect 154757 325214 158148 325216
rect 580165 325272 584960 325274
rect 580165 325216 580170 325272
rect 580226 325216 584960 325272
rect 580165 325214 584960 325216
rect 154757 325211 154823 325214
rect 580165 325211 580231 325214
rect 583520 325124 584960 325214
rect 154849 325002 154915 325005
rect 219893 325002 219959 325005
rect 154849 325000 158148 325002
rect 154849 324944 154854 325000
rect 154910 324944 158148 325000
rect 154849 324942 158148 324944
rect 217948 325000 219959 325002
rect 217948 324944 219898 325000
rect 219954 324944 219959 325000
rect 217948 324942 219959 324944
rect 154849 324939 154915 324942
rect 219893 324939 219959 324942
rect 154941 324730 155007 324733
rect 154941 324728 158148 324730
rect 154941 324672 154946 324728
rect 155002 324672 158148 324728
rect 154941 324670 158148 324672
rect 154941 324667 155007 324670
rect 220721 324594 220787 324597
rect 217948 324592 220787 324594
rect 217948 324536 220726 324592
rect 220782 324536 220787 324592
rect 217948 324534 220787 324536
rect 220721 324531 220787 324534
rect 154941 324458 155007 324461
rect 154941 324456 158148 324458
rect 154941 324400 154946 324456
rect 155002 324400 158148 324456
rect 154941 324398 158148 324400
rect 154941 324395 155007 324398
rect 155033 324186 155099 324189
rect 220261 324186 220327 324189
rect 155033 324184 158148 324186
rect 155033 324128 155038 324184
rect 155094 324128 158148 324184
rect 155033 324126 158148 324128
rect 217948 324184 220327 324186
rect 217948 324128 220266 324184
rect 220322 324128 220327 324184
rect 217948 324126 220327 324128
rect 155033 324123 155099 324126
rect 220261 324123 220327 324126
rect 153929 323914 153995 323917
rect 153929 323912 158148 323914
rect 153929 323856 153934 323912
rect 153990 323856 158148 323912
rect 153929 323854 158148 323856
rect 153929 323851 153995 323854
rect 220629 323778 220695 323781
rect 217948 323776 220695 323778
rect 217948 323720 220634 323776
rect 220690 323720 220695 323776
rect 217948 323718 220695 323720
rect 220629 323715 220695 323718
rect 154941 323642 155007 323645
rect 154941 323640 158148 323642
rect 154941 323584 154946 323640
rect 155002 323584 158148 323640
rect 154941 323582 158148 323584
rect 154941 323579 155007 323582
rect 154849 323370 154915 323373
rect 219709 323370 219775 323373
rect 154849 323368 158148 323370
rect 154849 323312 154854 323368
rect 154910 323312 158148 323368
rect 154849 323310 158148 323312
rect 217948 323368 219775 323370
rect 217948 323312 219714 323368
rect 219770 323312 219775 323368
rect 217948 323310 219775 323312
rect 154849 323307 154915 323310
rect 219709 323307 219775 323310
rect 154941 323098 155007 323101
rect 154941 323096 158148 323098
rect 154941 323040 154946 323096
rect 155002 323040 158148 323096
rect 154941 323038 158148 323040
rect 154941 323035 155007 323038
rect 220721 322962 220787 322965
rect 217948 322960 220787 322962
rect 217948 322904 220726 322960
rect 220782 322904 220787 322960
rect 217948 322902 220787 322904
rect 220721 322899 220787 322902
rect 155033 322826 155099 322829
rect 155033 322824 158148 322826
rect 155033 322768 155038 322824
rect 155094 322768 158148 322824
rect 155033 322766 158148 322768
rect 155033 322763 155099 322766
rect 154757 322554 154823 322557
rect 220537 322554 220603 322557
rect 154757 322552 158148 322554
rect 154757 322496 154762 322552
rect 154818 322496 158148 322552
rect 154757 322494 158148 322496
rect 217948 322552 220603 322554
rect 217948 322496 220542 322552
rect 220598 322496 220603 322552
rect 217948 322494 220603 322496
rect 154757 322491 154823 322494
rect 220537 322491 220603 322494
rect 154849 322282 154915 322285
rect 154849 322280 158148 322282
rect 154849 322224 154854 322280
rect 154910 322224 158148 322280
rect 154849 322222 158148 322224
rect 154849 322219 154915 322222
rect 220629 322146 220695 322149
rect 217948 322144 220695 322146
rect 217948 322088 220634 322144
rect 220690 322088 220695 322144
rect 217948 322086 220695 322088
rect 220629 322083 220695 322086
rect 154941 322010 155007 322013
rect 154941 322008 158148 322010
rect 154941 321952 154946 322008
rect 155002 321952 158148 322008
rect 154941 321950 158148 321952
rect 154941 321947 155007 321950
rect 154573 321738 154639 321741
rect 220721 321738 220787 321741
rect 154573 321736 158148 321738
rect 154573 321680 154578 321736
rect 154634 321680 158148 321736
rect 154573 321678 158148 321680
rect 217948 321736 220787 321738
rect 217948 321680 220726 321736
rect 220782 321680 220787 321736
rect 217948 321678 220787 321680
rect 154573 321675 154639 321678
rect 220721 321675 220787 321678
rect 155033 321466 155099 321469
rect 155033 321464 158148 321466
rect 155033 321408 155038 321464
rect 155094 321408 158148 321464
rect 155033 321406 158148 321408
rect 155033 321403 155099 321406
rect 220261 321330 220327 321333
rect 217948 321328 220327 321330
rect 217948 321272 220266 321328
rect 220322 321272 220327 321328
rect 217948 321270 220327 321272
rect 220261 321267 220327 321270
rect 154757 321194 154823 321197
rect 154757 321192 158148 321194
rect 154757 321136 154762 321192
rect 154818 321136 158148 321192
rect 154757 321134 158148 321136
rect 154757 321131 154823 321134
rect 154941 320922 155007 320925
rect 220721 320922 220787 320925
rect 154941 320920 158148 320922
rect 154941 320864 154946 320920
rect 155002 320864 158148 320920
rect 154941 320862 158148 320864
rect 217948 320920 220787 320922
rect 217948 320864 220726 320920
rect 220782 320864 220787 320920
rect 217948 320862 220787 320864
rect 154941 320859 155007 320862
rect 220721 320859 220787 320862
rect 154849 320650 154915 320653
rect 154849 320648 158148 320650
rect 154849 320592 154854 320648
rect 154910 320592 158148 320648
rect 154849 320590 158148 320592
rect 154849 320587 154915 320590
rect 220261 320514 220327 320517
rect 217948 320512 220327 320514
rect 217948 320456 220266 320512
rect 220322 320456 220327 320512
rect 217948 320454 220327 320456
rect 220261 320451 220327 320454
rect 154941 320378 155007 320381
rect 154941 320376 158148 320378
rect 154941 320320 154946 320376
rect 155002 320320 158148 320376
rect 154941 320318 158148 320320
rect 154941 320315 155007 320318
rect 154849 320106 154915 320109
rect 220445 320106 220511 320109
rect 154849 320104 158148 320106
rect 154849 320048 154854 320104
rect 154910 320048 158148 320104
rect 154849 320046 158148 320048
rect 217948 320104 220511 320106
rect 217948 320048 220450 320104
rect 220506 320048 220511 320104
rect 217948 320046 220511 320048
rect 154849 320043 154915 320046
rect 220445 320043 220511 320046
rect 154757 319834 154823 319837
rect 154757 319832 158148 319834
rect 154757 319776 154762 319832
rect 154818 319776 158148 319832
rect 154757 319774 158148 319776
rect 154757 319771 154823 319774
rect 220445 319698 220511 319701
rect 217948 319696 220511 319698
rect 217948 319640 220450 319696
rect 220506 319640 220511 319696
rect 217948 319638 220511 319640
rect 220445 319635 220511 319638
rect 155033 319562 155099 319565
rect 155033 319560 158148 319562
rect 155033 319504 155038 319560
rect 155094 319504 158148 319560
rect 155033 319502 158148 319504
rect 155033 319499 155099 319502
rect -960 319290 480 319380
rect 3417 319290 3483 319293
rect -960 319288 3483 319290
rect -960 319232 3422 319288
rect 3478 319232 3483 319288
rect -960 319230 3483 319232
rect -960 319140 480 319230
rect 3417 319227 3483 319230
rect 154941 319290 155007 319293
rect 220353 319290 220419 319293
rect 154941 319288 158148 319290
rect 154941 319232 154946 319288
rect 155002 319232 158148 319288
rect 154941 319230 158148 319232
rect 217948 319288 220419 319290
rect 217948 319232 220358 319288
rect 220414 319232 220419 319288
rect 217948 319230 220419 319232
rect 154941 319227 155007 319230
rect 220353 319227 220419 319230
rect 155493 319018 155559 319021
rect 155493 319016 158148 319018
rect 155493 318960 155498 319016
rect 155554 318960 158148 319016
rect 155493 318958 158148 318960
rect 155493 318955 155559 318958
rect 220721 318882 220787 318885
rect 217948 318880 220787 318882
rect 217948 318824 220726 318880
rect 220782 318824 220787 318880
rect 217948 318822 220787 318824
rect 220721 318819 220787 318822
rect 154665 318746 154731 318749
rect 154665 318744 158148 318746
rect 154665 318688 154670 318744
rect 154726 318688 158148 318744
rect 154665 318686 158148 318688
rect 154665 318683 154731 318686
rect 154757 318474 154823 318477
rect 219985 318474 220051 318477
rect 154757 318472 158148 318474
rect 154757 318416 154762 318472
rect 154818 318416 158148 318472
rect 154757 318414 158148 318416
rect 217948 318472 220051 318474
rect 217948 318416 219990 318472
rect 220046 318416 220051 318472
rect 217948 318414 220051 318416
rect 154757 318411 154823 318414
rect 219985 318411 220051 318414
rect 155033 318202 155099 318205
rect 155033 318200 158148 318202
rect 155033 318144 155038 318200
rect 155094 318144 158148 318200
rect 155033 318142 158148 318144
rect 155033 318139 155099 318142
rect 220629 318066 220695 318069
rect 217948 318064 220695 318066
rect 217948 318008 220634 318064
rect 220690 318008 220695 318064
rect 217948 318006 220695 318008
rect 220629 318003 220695 318006
rect 154849 317930 154915 317933
rect 154849 317928 158148 317930
rect 154849 317872 154854 317928
rect 154910 317872 158148 317928
rect 154849 317870 158148 317872
rect 154849 317867 154915 317870
rect 154941 317658 155007 317661
rect 220721 317658 220787 317661
rect 154941 317656 158148 317658
rect 154941 317600 154946 317656
rect 155002 317600 158148 317656
rect 154941 317598 158148 317600
rect 217948 317656 220787 317658
rect 217948 317600 220726 317656
rect 220782 317600 220787 317656
rect 217948 317598 220787 317600
rect 154941 317595 155007 317598
rect 220721 317595 220787 317598
rect 154757 317386 154823 317389
rect 154757 317384 158148 317386
rect 154757 317328 154762 317384
rect 154818 317328 158148 317384
rect 154757 317326 158148 317328
rect 154757 317323 154823 317326
rect 220721 317250 220787 317253
rect 217948 317248 220787 317250
rect 217948 317192 220726 317248
rect 220782 317192 220787 317248
rect 217948 317190 220787 317192
rect 220721 317187 220787 317190
rect 154849 317114 154915 317117
rect 154849 317112 158148 317114
rect 154849 317056 154854 317112
rect 154910 317056 158148 317112
rect 154849 317054 158148 317056
rect 154849 317051 154915 317054
rect 154573 316842 154639 316845
rect 220629 316842 220695 316845
rect 154573 316840 158148 316842
rect 154573 316784 154578 316840
rect 154634 316784 158148 316840
rect 154573 316782 158148 316784
rect 217948 316840 220695 316842
rect 217948 316784 220634 316840
rect 220690 316784 220695 316840
rect 217948 316782 220695 316784
rect 154573 316779 154639 316782
rect 220629 316779 220695 316782
rect 155033 316570 155099 316573
rect 155033 316568 158148 316570
rect 155033 316512 155038 316568
rect 155094 316512 158148 316568
rect 155033 316510 158148 316512
rect 155033 316507 155099 316510
rect 220445 316434 220511 316437
rect 217948 316432 220511 316434
rect 217948 316376 220450 316432
rect 220506 316376 220511 316432
rect 217948 316374 220511 316376
rect 220445 316371 220511 316374
rect 154941 316298 155007 316301
rect 154941 316296 158148 316298
rect 154941 316240 154946 316296
rect 155002 316240 158148 316296
rect 154941 316238 158148 316240
rect 154941 316235 155007 316238
rect 155033 316026 155099 316029
rect 220629 316026 220695 316029
rect 155033 316024 158148 316026
rect 155033 315968 155038 316024
rect 155094 315968 158148 316024
rect 155033 315966 158148 315968
rect 217948 316024 220695 316026
rect 217948 315968 220634 316024
rect 220690 315968 220695 316024
rect 217948 315966 220695 315968
rect 155033 315963 155099 315966
rect 220629 315963 220695 315966
rect 154849 315754 154915 315757
rect 154849 315752 158148 315754
rect 154849 315696 154854 315752
rect 154910 315696 158148 315752
rect 154849 315694 158148 315696
rect 154849 315691 154915 315694
rect 219985 315618 220051 315621
rect 217948 315616 220051 315618
rect 217948 315560 219990 315616
rect 220046 315560 220051 315616
rect 217948 315558 220051 315560
rect 219985 315555 220051 315558
rect 154757 315482 154823 315485
rect 154757 315480 158148 315482
rect 154757 315424 154762 315480
rect 154818 315424 158148 315480
rect 154757 315422 158148 315424
rect 154757 315419 154823 315422
rect 154941 315210 155007 315213
rect 220721 315210 220787 315213
rect 154941 315208 158148 315210
rect 154941 315152 154946 315208
rect 155002 315152 158148 315208
rect 154941 315150 158148 315152
rect 217948 315208 220787 315210
rect 217948 315152 220726 315208
rect 220782 315152 220787 315208
rect 217948 315150 220787 315152
rect 154941 315147 155007 315150
rect 220721 315147 220787 315150
rect 155585 314938 155651 314941
rect 155585 314936 158148 314938
rect 155585 314880 155590 314936
rect 155646 314880 158148 314936
rect 155585 314878 158148 314880
rect 155585 314875 155651 314878
rect 220537 314802 220603 314805
rect 217948 314800 220603 314802
rect 217948 314744 220542 314800
rect 220598 314744 220603 314800
rect 217948 314742 220603 314744
rect 220537 314739 220603 314742
rect 154757 314666 154823 314669
rect 154757 314664 158148 314666
rect 154757 314608 154762 314664
rect 154818 314608 158148 314664
rect 154757 314606 158148 314608
rect 154757 314603 154823 314606
rect 154849 314394 154915 314397
rect 220629 314394 220695 314397
rect 154849 314392 158148 314394
rect 154849 314336 154854 314392
rect 154910 314336 158148 314392
rect 154849 314334 158148 314336
rect 217948 314392 220695 314394
rect 217948 314336 220634 314392
rect 220690 314336 220695 314392
rect 217948 314334 220695 314336
rect 154849 314331 154915 314334
rect 220629 314331 220695 314334
rect 111793 314258 111859 314261
rect 109910 314256 111859 314258
rect 109910 314200 111798 314256
rect 111854 314200 111859 314256
rect 109910 314198 111859 314200
rect 109910 313752 109970 314198
rect 111793 314195 111859 314198
rect 155677 314122 155743 314125
rect 155677 314120 158148 314122
rect 155677 314064 155682 314120
rect 155738 314064 158148 314120
rect 155677 314062 158148 314064
rect 155677 314059 155743 314062
rect 220445 313986 220511 313989
rect 217948 313984 220511 313986
rect 217948 313928 220450 313984
rect 220506 313928 220511 313984
rect 217948 313926 220511 313928
rect 220445 313923 220511 313926
rect 154573 313850 154639 313853
rect 154573 313848 158148 313850
rect 154573 313792 154578 313848
rect 154634 313792 158148 313848
rect 154573 313790 158148 313792
rect 154573 313787 154639 313790
rect 154941 313578 155007 313581
rect 220721 313578 220787 313581
rect 154941 313576 158148 313578
rect 154941 313520 154946 313576
rect 155002 313520 158148 313576
rect 154941 313518 158148 313520
rect 217948 313576 220787 313578
rect 217948 313520 220726 313576
rect 220782 313520 220787 313576
rect 217948 313518 220787 313520
rect 154941 313515 155007 313518
rect 220721 313515 220787 313518
rect 154941 313306 155007 313309
rect 154941 313304 158148 313306
rect 154941 313248 154946 313304
rect 155002 313248 158148 313304
rect 154941 313246 158148 313248
rect 154941 313243 155007 313246
rect 111793 313170 111859 313173
rect 219893 313170 219959 313173
rect 109910 313168 111859 313170
rect 109910 313112 111798 313168
rect 111854 313112 111859 313168
rect 109910 313110 111859 313112
rect 217948 313168 219959 313170
rect 217948 313112 219898 313168
rect 219954 313112 219959 313168
rect 217948 313110 219959 313112
rect 109910 313072 109970 313110
rect 111793 313107 111859 313110
rect 219893 313107 219959 313110
rect 154849 313034 154915 313037
rect 154849 313032 158148 313034
rect 154849 312976 154854 313032
rect 154910 312976 158148 313032
rect 154849 312974 158148 312976
rect 154849 312971 154915 312974
rect 111885 312762 111951 312765
rect 109910 312760 111951 312762
rect 109910 312704 111890 312760
rect 111946 312704 111951 312760
rect 109910 312702 111951 312704
rect 109910 312392 109970 312702
rect 111885 312699 111951 312702
rect 154757 312762 154823 312765
rect 220445 312762 220511 312765
rect 154757 312760 158148 312762
rect 154757 312704 154762 312760
rect 154818 312704 158148 312760
rect 154757 312702 158148 312704
rect 217948 312760 220511 312762
rect 217948 312704 220450 312760
rect 220506 312704 220511 312760
rect 217948 312702 220511 312704
rect 154757 312699 154823 312702
rect 220445 312699 220511 312702
rect 154573 312490 154639 312493
rect 154573 312488 158148 312490
rect 154573 312432 154578 312488
rect 154634 312432 158148 312488
rect 154573 312430 158148 312432
rect 154573 312427 154639 312430
rect 220445 312354 220511 312357
rect 217948 312352 220511 312354
rect 217948 312296 220450 312352
rect 220506 312296 220511 312352
rect 217948 312294 220511 312296
rect 220445 312291 220511 312294
rect 154941 312218 155007 312221
rect 154941 312216 158148 312218
rect 154941 312160 154946 312216
rect 155002 312160 158148 312216
rect 154941 312158 158148 312160
rect 154941 312155 155007 312158
rect 580441 312082 580507 312085
rect 583520 312082 584960 312172
rect 580441 312080 584960 312082
rect 580441 312024 580446 312080
rect 580502 312024 584960 312080
rect 580441 312022 584960 312024
rect 580441 312019 580507 312022
rect 154573 311946 154639 311949
rect 220721 311946 220787 311949
rect 154573 311944 158148 311946
rect 154573 311888 154578 311944
rect 154634 311888 158148 311944
rect 154573 311886 158148 311888
rect 217948 311944 220787 311946
rect 217948 311888 220726 311944
rect 220782 311888 220787 311944
rect 583520 311932 584960 312022
rect 217948 311886 220787 311888
rect 154573 311883 154639 311886
rect 220721 311883 220787 311886
rect 111793 311810 111859 311813
rect 109910 311808 111859 311810
rect 109910 311752 111798 311808
rect 111854 311752 111859 311808
rect 109910 311750 111859 311752
rect 109910 311712 109970 311750
rect 111793 311747 111859 311750
rect 154757 311674 154823 311677
rect 154757 311672 158148 311674
rect 154757 311616 154762 311672
rect 154818 311616 158148 311672
rect 154757 311614 158148 311616
rect 154757 311611 154823 311614
rect 220629 311538 220695 311541
rect 217948 311536 220695 311538
rect 217948 311480 220634 311536
rect 220690 311480 220695 311536
rect 217948 311478 220695 311480
rect 220629 311475 220695 311478
rect 111885 311402 111951 311405
rect 109910 311400 111951 311402
rect 109910 311344 111890 311400
rect 111946 311344 111951 311400
rect 109910 311342 111951 311344
rect 109910 311032 109970 311342
rect 111885 311339 111951 311342
rect 154849 311402 154915 311405
rect 154849 311400 158148 311402
rect 154849 311344 154854 311400
rect 154910 311344 158148 311400
rect 154849 311342 158148 311344
rect 154849 311339 154915 311342
rect 155033 311130 155099 311133
rect 220721 311130 220787 311133
rect 155033 311128 158148 311130
rect 155033 311072 155038 311128
rect 155094 311072 158148 311128
rect 155033 311070 158148 311072
rect 217948 311128 220787 311130
rect 217948 311072 220726 311128
rect 220782 311072 220787 311128
rect 217948 311070 220787 311072
rect 155033 311067 155099 311070
rect 220721 311067 220787 311070
rect 154941 310858 155007 310861
rect 154941 310856 158148 310858
rect 154941 310800 154946 310856
rect 155002 310800 158148 310856
rect 154941 310798 158148 310800
rect 154941 310795 155007 310798
rect 220537 310722 220603 310725
rect 217948 310720 220603 310722
rect 217948 310664 220542 310720
rect 220598 310664 220603 310720
rect 217948 310662 220603 310664
rect 220537 310659 220603 310662
rect 154849 310586 154915 310589
rect 256693 310586 256759 310589
rect 154849 310584 158148 310586
rect 154849 310528 154854 310584
rect 154910 310528 158148 310584
rect 154849 310526 158148 310528
rect 256693 310584 260084 310586
rect 256693 310528 256698 310584
rect 256754 310528 260084 310584
rect 256693 310526 260084 310528
rect 154849 310523 154915 310526
rect 256693 310523 256759 310526
rect 111793 310450 111859 310453
rect 109910 310448 111859 310450
rect 109910 310392 111798 310448
rect 111854 310392 111859 310448
rect 109910 310390 111859 310392
rect 109910 310352 109970 310390
rect 111793 310387 111859 310390
rect 154849 310314 154915 310317
rect 220721 310314 220787 310317
rect 154849 310312 158148 310314
rect 154849 310256 154854 310312
rect 154910 310256 158148 310312
rect 154849 310254 158148 310256
rect 217948 310312 220787 310314
rect 217948 310256 220726 310312
rect 220782 310256 220787 310312
rect 217948 310254 220787 310256
rect 154849 310251 154915 310254
rect 220721 310251 220787 310254
rect 111885 310042 111951 310045
rect 109910 310040 111951 310042
rect 109910 309984 111890 310040
rect 111946 309984 111951 310040
rect 109910 309982 111951 309984
rect 109910 309672 109970 309982
rect 111885 309979 111951 309982
rect 154757 310042 154823 310045
rect 154757 310040 158148 310042
rect 154757 309984 154762 310040
rect 154818 309984 158148 310040
rect 154757 309982 158148 309984
rect 154757 309979 154823 309982
rect 220537 309906 220603 309909
rect 217948 309904 220603 309906
rect 217948 309848 220542 309904
rect 220598 309848 220603 309904
rect 217948 309846 220603 309848
rect 220537 309843 220603 309846
rect 154573 309770 154639 309773
rect 154573 309768 158148 309770
rect 154573 309712 154578 309768
rect 154634 309712 158148 309768
rect 154573 309710 158148 309712
rect 154573 309707 154639 309710
rect 154941 309498 155007 309501
rect 220629 309498 220695 309501
rect 154941 309496 158148 309498
rect 154941 309440 154946 309496
rect 155002 309440 158148 309496
rect 154941 309438 158148 309440
rect 217948 309496 220695 309498
rect 217948 309440 220634 309496
rect 220690 309440 220695 309496
rect 217948 309438 220695 309440
rect 154941 309435 155007 309438
rect 220629 309435 220695 309438
rect 154941 309226 155007 309229
rect 154941 309224 158148 309226
rect 154941 309168 154946 309224
rect 155002 309168 158148 309224
rect 154941 309166 158148 309168
rect 154941 309163 155007 309166
rect 111793 309090 111859 309093
rect 219709 309090 219775 309093
rect 109910 309088 111859 309090
rect 109910 309032 111798 309088
rect 111854 309032 111859 309088
rect 109910 309030 111859 309032
rect 217948 309088 219775 309090
rect 217948 309032 219714 309088
rect 219770 309032 219775 309088
rect 217948 309030 219775 309032
rect 109910 308992 109970 309030
rect 111793 309027 111859 309030
rect 219709 309027 219775 309030
rect 155033 308954 155099 308957
rect 155033 308952 158148 308954
rect 155033 308896 155038 308952
rect 155094 308896 158148 308952
rect 155033 308894 158148 308896
rect 155033 308891 155099 308894
rect 111885 308682 111951 308685
rect 109910 308680 111951 308682
rect 109910 308624 111890 308680
rect 111946 308624 111951 308680
rect 109910 308622 111951 308624
rect 109910 308312 109970 308622
rect 111885 308619 111951 308622
rect 154757 308682 154823 308685
rect 219893 308682 219959 308685
rect 154757 308680 158148 308682
rect 154757 308624 154762 308680
rect 154818 308624 158148 308680
rect 154757 308622 158148 308624
rect 217948 308680 219959 308682
rect 217948 308624 219898 308680
rect 219954 308624 219959 308680
rect 217948 308622 219959 308624
rect 154757 308619 154823 308622
rect 219893 308619 219959 308622
rect 256693 308546 256759 308549
rect 256693 308544 260084 308546
rect 256693 308488 256698 308544
rect 256754 308488 260084 308544
rect 256693 308486 260084 308488
rect 256693 308483 256759 308486
rect 154849 308410 154915 308413
rect 154849 308408 158148 308410
rect 154849 308352 154854 308408
rect 154910 308352 158148 308408
rect 154849 308350 158148 308352
rect 154849 308347 154915 308350
rect 220629 308274 220695 308277
rect 217948 308272 220695 308274
rect 217948 308216 220634 308272
rect 220690 308216 220695 308272
rect 217948 308214 220695 308216
rect 220629 308211 220695 308214
rect 154573 308138 154639 308141
rect 154573 308136 158148 308138
rect 154573 308080 154578 308136
rect 154634 308080 158148 308136
rect 154573 308078 158148 308080
rect 154573 308075 154639 308078
rect 154941 307866 155007 307869
rect 220721 307866 220787 307869
rect 154941 307864 158148 307866
rect 154941 307808 154946 307864
rect 155002 307808 158148 307864
rect 154941 307806 158148 307808
rect 217948 307864 220787 307866
rect 217948 307808 220726 307864
rect 220782 307808 220787 307864
rect 217948 307806 220787 307808
rect 154941 307803 155007 307806
rect 220721 307803 220787 307806
rect 111793 307730 111859 307733
rect 109910 307728 111859 307730
rect 109910 307672 111798 307728
rect 111854 307672 111859 307728
rect 109910 307670 111859 307672
rect 109910 307632 109970 307670
rect 111793 307667 111859 307670
rect 155033 307594 155099 307597
rect 155033 307592 158148 307594
rect 155033 307536 155038 307592
rect 155094 307536 158148 307592
rect 155033 307534 158148 307536
rect 155033 307531 155099 307534
rect 220537 307458 220603 307461
rect 217948 307456 220603 307458
rect 217948 307400 220542 307456
rect 220598 307400 220603 307456
rect 217948 307398 220603 307400
rect 220537 307395 220603 307398
rect 111793 307322 111859 307325
rect 109910 307320 111859 307322
rect 109910 307264 111798 307320
rect 111854 307264 111859 307320
rect 109910 307262 111859 307264
rect 109910 306952 109970 307262
rect 111793 307259 111859 307262
rect 154757 307322 154823 307325
rect 154757 307320 158148 307322
rect 154757 307264 154762 307320
rect 154818 307264 158148 307320
rect 154757 307262 158148 307264
rect 154757 307259 154823 307262
rect 154941 307050 155007 307053
rect 220629 307050 220695 307053
rect 154941 307048 158148 307050
rect 154941 306992 154946 307048
rect 155002 306992 158148 307048
rect 154941 306990 158148 306992
rect 217948 307048 220695 307050
rect 217948 306992 220634 307048
rect 220690 306992 220695 307048
rect 217948 306990 220695 306992
rect 154941 306987 155007 306990
rect 220629 306987 220695 306990
rect 154849 306778 154915 306781
rect 154849 306776 158148 306778
rect 154849 306720 154854 306776
rect 154910 306720 158148 306776
rect 154849 306718 158148 306720
rect 154849 306715 154915 306718
rect 220721 306642 220787 306645
rect 217948 306640 220787 306642
rect 217948 306584 220726 306640
rect 220782 306584 220787 306640
rect 217948 306582 220787 306584
rect 220721 306579 220787 306582
rect 154941 306506 155007 306509
rect 256785 306506 256851 306509
rect 154941 306504 158148 306506
rect 154941 306448 154946 306504
rect 155002 306448 158148 306504
rect 154941 306446 158148 306448
rect 256785 306504 260084 306506
rect 256785 306448 256790 306504
rect 256846 306448 260084 306504
rect 256785 306446 260084 306448
rect 154941 306443 155007 306446
rect 256785 306443 256851 306446
rect 111793 306370 111859 306373
rect 109910 306368 111859 306370
rect -960 306234 480 306324
rect 109910 306312 111798 306368
rect 111854 306312 111859 306368
rect 109910 306310 111859 306312
rect 109910 306272 109970 306310
rect 111793 306307 111859 306310
rect 3233 306234 3299 306237
rect -960 306232 3299 306234
rect -960 306176 3238 306232
rect 3294 306176 3299 306232
rect -960 306174 3299 306176
rect -960 306084 480 306174
rect 3233 306171 3299 306174
rect 154849 306234 154915 306237
rect 220537 306234 220603 306237
rect 154849 306232 158148 306234
rect 154849 306176 154854 306232
rect 154910 306176 158148 306232
rect 154849 306174 158148 306176
rect 217948 306232 220603 306234
rect 217948 306176 220542 306232
rect 220598 306176 220603 306232
rect 217948 306174 220603 306176
rect 154849 306171 154915 306174
rect 220537 306171 220603 306174
rect 111885 305962 111951 305965
rect 109910 305960 111951 305962
rect 109910 305904 111890 305960
rect 111946 305904 111951 305960
rect 109910 305902 111951 305904
rect 109910 305592 109970 305902
rect 111885 305899 111951 305902
rect 154757 305962 154823 305965
rect 154757 305960 158148 305962
rect 154757 305904 154762 305960
rect 154818 305904 158148 305960
rect 154757 305902 158148 305904
rect 154757 305899 154823 305902
rect 220629 305826 220695 305829
rect 217948 305824 220695 305826
rect 217948 305768 220634 305824
rect 220690 305768 220695 305824
rect 217948 305766 220695 305768
rect 220629 305763 220695 305766
rect 155585 305690 155651 305693
rect 155585 305688 158148 305690
rect 155585 305632 155590 305688
rect 155646 305632 158148 305688
rect 155585 305630 158148 305632
rect 155585 305627 155651 305630
rect 154941 305418 155007 305421
rect 220721 305418 220787 305421
rect 154941 305416 158148 305418
rect 154941 305360 154946 305416
rect 155002 305360 158148 305416
rect 154941 305358 158148 305360
rect 217948 305416 220787 305418
rect 217948 305360 220726 305416
rect 220782 305360 220787 305416
rect 217948 305358 220787 305360
rect 154941 305355 155007 305358
rect 220721 305355 220787 305358
rect 155125 305146 155191 305149
rect 155125 305144 158148 305146
rect 155125 305088 155130 305144
rect 155186 305088 158148 305144
rect 155125 305086 158148 305088
rect 155125 305083 155191 305086
rect 220721 305010 220787 305013
rect 217948 305008 220787 305010
rect 217948 304952 220726 305008
rect 220782 304952 220787 305008
rect 217948 304950 220787 304952
rect 220721 304947 220787 304950
rect 109910 304874 109970 304912
rect 111793 304874 111859 304877
rect 109910 304872 111859 304874
rect 109910 304816 111798 304872
rect 111854 304816 111859 304872
rect 109910 304814 111859 304816
rect 111793 304811 111859 304814
rect 154849 304874 154915 304877
rect 154849 304872 158148 304874
rect 154849 304816 154854 304872
rect 154910 304816 158148 304872
rect 154849 304814 158148 304816
rect 154849 304811 154915 304814
rect 111885 304602 111951 304605
rect 109910 304600 111951 304602
rect 109910 304544 111890 304600
rect 111946 304544 111951 304600
rect 109910 304542 111951 304544
rect 109910 304232 109970 304542
rect 111885 304539 111951 304542
rect 154941 304602 155007 304605
rect 220445 304602 220511 304605
rect 154941 304600 158148 304602
rect 154941 304544 154946 304600
rect 155002 304544 158148 304600
rect 154941 304542 158148 304544
rect 217948 304600 220511 304602
rect 217948 304544 220450 304600
rect 220506 304544 220511 304600
rect 217948 304542 220511 304544
rect 154941 304539 155007 304542
rect 220445 304539 220511 304542
rect 257705 304466 257771 304469
rect 257705 304464 260084 304466
rect 257705 304408 257710 304464
rect 257766 304408 260084 304464
rect 257705 304406 260084 304408
rect 257705 304403 257771 304406
rect 155493 304330 155559 304333
rect 155493 304328 158148 304330
rect 155493 304272 155498 304328
rect 155554 304272 158148 304328
rect 155493 304270 158148 304272
rect 155493 304267 155559 304270
rect 220629 304194 220695 304197
rect 217948 304192 220695 304194
rect 217948 304136 220634 304192
rect 220690 304136 220695 304192
rect 217948 304134 220695 304136
rect 220629 304131 220695 304134
rect 154573 304058 154639 304061
rect 154573 304056 158148 304058
rect 154573 304000 154578 304056
rect 154634 304000 158148 304056
rect 154573 303998 158148 304000
rect 154573 303995 154639 303998
rect 154757 303786 154823 303789
rect 220721 303786 220787 303789
rect 154757 303784 158148 303786
rect 154757 303728 154762 303784
rect 154818 303728 158148 303784
rect 154757 303726 158148 303728
rect 217948 303784 220787 303786
rect 217948 303728 220726 303784
rect 220782 303728 220787 303784
rect 217948 303726 220787 303728
rect 154757 303723 154823 303726
rect 220721 303723 220787 303726
rect 109910 303514 109970 303552
rect 111793 303514 111859 303517
rect 109910 303512 111859 303514
rect 109910 303456 111798 303512
rect 111854 303456 111859 303512
rect 109910 303454 111859 303456
rect 111793 303451 111859 303454
rect 154941 303514 155007 303517
rect 154941 303512 158148 303514
rect 154941 303456 154946 303512
rect 155002 303456 158148 303512
rect 154941 303454 158148 303456
rect 154941 303451 155007 303454
rect 220537 303378 220603 303381
rect 217948 303376 220603 303378
rect 217948 303320 220542 303376
rect 220598 303320 220603 303376
rect 217948 303318 220603 303320
rect 220537 303315 220603 303318
rect 111885 303242 111951 303245
rect 109910 303240 111951 303242
rect 109910 303184 111890 303240
rect 111946 303184 111951 303240
rect 109910 303182 111951 303184
rect 109910 302872 109970 303182
rect 111885 303179 111951 303182
rect 155125 303242 155191 303245
rect 155125 303240 158148 303242
rect 155125 303184 155130 303240
rect 155186 303184 158148 303240
rect 155125 303182 158148 303184
rect 155125 303179 155191 303182
rect 154849 302970 154915 302973
rect 219893 302970 219959 302973
rect 154849 302968 158148 302970
rect 154849 302912 154854 302968
rect 154910 302912 158148 302968
rect 154849 302910 158148 302912
rect 217948 302968 219959 302970
rect 217948 302912 219898 302968
rect 219954 302912 219959 302968
rect 217948 302910 219959 302912
rect 154849 302907 154915 302910
rect 219893 302907 219959 302910
rect 153837 302698 153903 302701
rect 153837 302696 158148 302698
rect 153837 302640 153842 302696
rect 153898 302640 158148 302696
rect 153837 302638 158148 302640
rect 153837 302635 153903 302638
rect 220721 302562 220787 302565
rect 217948 302560 220787 302562
rect 217948 302504 220726 302560
rect 220782 302504 220787 302560
rect 217948 302502 220787 302504
rect 220721 302499 220787 302502
rect 154665 302426 154731 302429
rect 256693 302426 256759 302429
rect 154665 302424 158148 302426
rect 154665 302368 154670 302424
rect 154726 302368 158148 302424
rect 154665 302366 158148 302368
rect 256693 302424 260084 302426
rect 256693 302368 256698 302424
rect 256754 302368 260084 302424
rect 256693 302366 260084 302368
rect 154665 302363 154731 302366
rect 256693 302363 256759 302366
rect 109910 302154 109970 302192
rect 111793 302154 111859 302157
rect 109910 302152 111859 302154
rect 109910 302096 111798 302152
rect 111854 302096 111859 302152
rect 109910 302094 111859 302096
rect 111793 302091 111859 302094
rect 154849 302154 154915 302157
rect 220629 302154 220695 302157
rect 154849 302152 158148 302154
rect 154849 302096 154854 302152
rect 154910 302096 158148 302152
rect 154849 302094 158148 302096
rect 217948 302152 220695 302154
rect 217948 302096 220634 302152
rect 220690 302096 220695 302152
rect 217948 302094 220695 302096
rect 154849 302091 154915 302094
rect 220629 302091 220695 302094
rect 111885 301882 111951 301885
rect 109910 301880 111951 301882
rect 109910 301824 111890 301880
rect 111946 301824 111951 301880
rect 109910 301822 111951 301824
rect 109910 301512 109970 301822
rect 111885 301819 111951 301822
rect 154757 301882 154823 301885
rect 154757 301880 158148 301882
rect 154757 301824 154762 301880
rect 154818 301824 158148 301880
rect 154757 301822 158148 301824
rect 154757 301819 154823 301822
rect 220537 301746 220603 301749
rect 217948 301744 220603 301746
rect 217948 301688 220542 301744
rect 220598 301688 220603 301744
rect 217948 301686 220603 301688
rect 220537 301683 220603 301686
rect 154665 301610 154731 301613
rect 154665 301608 158148 301610
rect 154665 301552 154670 301608
rect 154726 301552 158148 301608
rect 154665 301550 158148 301552
rect 154665 301547 154731 301550
rect 154573 301338 154639 301341
rect 219985 301338 220051 301341
rect 154573 301336 158148 301338
rect 154573 301280 154578 301336
rect 154634 301280 158148 301336
rect 154573 301278 158148 301280
rect 217948 301336 220051 301338
rect 217948 301280 219990 301336
rect 220046 301280 220051 301336
rect 217948 301278 220051 301280
rect 154573 301275 154639 301278
rect 219985 301275 220051 301278
rect 155585 301066 155651 301069
rect 155585 301064 158148 301066
rect 155585 301008 155590 301064
rect 155646 301008 158148 301064
rect 155585 301006 158148 301008
rect 155585 301003 155651 301006
rect 220721 300930 220787 300933
rect 217948 300928 220787 300930
rect 217948 300872 220726 300928
rect 220782 300872 220787 300928
rect 217948 300870 220787 300872
rect 220721 300867 220787 300870
rect 109910 300794 109970 300832
rect 111885 300794 111951 300797
rect 109910 300792 111951 300794
rect 109910 300736 111890 300792
rect 111946 300736 111951 300792
rect 109910 300734 111951 300736
rect 111885 300731 111951 300734
rect 155309 300794 155375 300797
rect 155309 300792 158148 300794
rect 155309 300736 155314 300792
rect 155370 300736 158148 300792
rect 155309 300734 158148 300736
rect 155309 300731 155375 300734
rect 154849 300522 154915 300525
rect 154849 300520 158148 300522
rect 154849 300464 154854 300520
rect 154910 300464 158148 300520
rect 154849 300462 158148 300464
rect 154849 300459 154915 300462
rect 111793 300386 111859 300389
rect 109910 300384 111859 300386
rect 109910 300328 111798 300384
rect 111854 300328 111859 300384
rect 109910 300326 111859 300328
rect 217918 300386 217978 300492
rect 224166 300386 224172 300388
rect 217918 300326 224172 300386
rect 109910 300152 109970 300326
rect 111793 300323 111859 300326
rect 224166 300324 224172 300326
rect 224236 300324 224242 300388
rect 256693 300386 256759 300389
rect 256693 300384 260084 300386
rect 256693 300328 256698 300384
rect 256754 300328 260084 300384
rect 256693 300326 260084 300328
rect 256693 300323 256759 300326
rect 154757 300250 154823 300253
rect 154757 300248 158148 300250
rect 154757 300192 154762 300248
rect 154818 300192 158148 300248
rect 154757 300190 158148 300192
rect 154757 300187 154823 300190
rect 220629 300114 220695 300117
rect 217948 300112 220695 300114
rect 217948 300056 220634 300112
rect 220690 300056 220695 300112
rect 217948 300054 220695 300056
rect 220629 300051 220695 300054
rect 111977 299978 112043 299981
rect 109910 299976 112043 299978
rect 109910 299920 111982 299976
rect 112038 299920 112043 299976
rect 109910 299918 112043 299920
rect 109910 299472 109970 299918
rect 111977 299915 112043 299918
rect 154665 299978 154731 299981
rect 154665 299976 158148 299978
rect 154665 299920 154670 299976
rect 154726 299920 158148 299976
rect 154665 299918 158148 299920
rect 154665 299915 154731 299918
rect 154573 299706 154639 299709
rect 220721 299706 220787 299709
rect 154573 299704 158148 299706
rect 154573 299648 154578 299704
rect 154634 299648 158148 299704
rect 154573 299646 158148 299648
rect 217948 299704 220787 299706
rect 217948 299648 220726 299704
rect 220782 299648 220787 299704
rect 217948 299646 220787 299648
rect 154573 299643 154639 299646
rect 220721 299643 220787 299646
rect 154757 299434 154823 299437
rect 154757 299432 158148 299434
rect 154757 299376 154762 299432
rect 154818 299376 158148 299432
rect 154757 299374 158148 299376
rect 154757 299371 154823 299374
rect 220537 299298 220603 299301
rect 217948 299296 220603 299298
rect 217948 299240 220542 299296
rect 220598 299240 220603 299296
rect 217948 299238 220603 299240
rect 220537 299235 220603 299238
rect 154941 299162 155007 299165
rect 154941 299160 158148 299162
rect 154941 299104 154946 299160
rect 155002 299104 158148 299160
rect 154941 299102 158148 299104
rect 154941 299099 155007 299102
rect 111793 299026 111859 299029
rect 109910 299024 111859 299026
rect 109910 298968 111798 299024
rect 111854 298968 111859 299024
rect 109910 298966 111859 298968
rect 109910 298792 109970 298966
rect 111793 298963 111859 298966
rect 154573 298890 154639 298893
rect 219985 298890 220051 298893
rect 154573 298888 158148 298890
rect 154573 298832 154578 298888
rect 154634 298832 158148 298888
rect 154573 298830 158148 298832
rect 217948 298888 220051 298890
rect 217948 298832 219990 298888
rect 220046 298832 220051 298888
rect 217948 298830 220051 298832
rect 154573 298827 154639 298830
rect 219985 298827 220051 298830
rect 580257 298754 580323 298757
rect 583520 298754 584960 298844
rect 580257 298752 584960 298754
rect 580257 298696 580262 298752
rect 580318 298696 584960 298752
rect 580257 298694 584960 298696
rect 580257 298691 580323 298694
rect 154849 298618 154915 298621
rect 154849 298616 158148 298618
rect 154849 298560 154854 298616
rect 154910 298560 158148 298616
rect 583520 298604 584960 298694
rect 154849 298558 158148 298560
rect 154849 298555 154915 298558
rect 111793 298482 111859 298485
rect 220721 298482 220787 298485
rect 109910 298480 111859 298482
rect 109910 298424 111798 298480
rect 111854 298424 111859 298480
rect 109910 298422 111859 298424
rect 217948 298480 220787 298482
rect 217948 298424 220726 298480
rect 220782 298424 220787 298480
rect 217948 298422 220787 298424
rect 109910 298112 109970 298422
rect 111793 298419 111859 298422
rect 220721 298419 220787 298422
rect 154665 298346 154731 298349
rect 256693 298346 256759 298349
rect 154665 298344 158148 298346
rect 154665 298288 154670 298344
rect 154726 298288 158148 298344
rect 154665 298286 158148 298288
rect 256693 298344 260084 298346
rect 256693 298288 256698 298344
rect 256754 298288 260084 298344
rect 256693 298286 260084 298288
rect 154665 298283 154731 298286
rect 256693 298283 256759 298286
rect 154941 298074 155007 298077
rect 220629 298074 220695 298077
rect 154941 298072 158148 298074
rect 154941 298016 154946 298072
rect 155002 298016 158148 298072
rect 154941 298014 158148 298016
rect 217948 298072 220695 298074
rect 217948 298016 220634 298072
rect 220690 298016 220695 298072
rect 217948 298014 220695 298016
rect 154941 298011 155007 298014
rect 220629 298011 220695 298014
rect 154757 297802 154823 297805
rect 154757 297800 158148 297802
rect 154757 297744 154762 297800
rect 154818 297744 158148 297800
rect 154757 297742 158148 297744
rect 154757 297739 154823 297742
rect 111793 297666 111859 297669
rect 220721 297666 220787 297669
rect 109910 297664 111859 297666
rect 109910 297608 111798 297664
rect 111854 297608 111859 297664
rect 109910 297606 111859 297608
rect 217948 297664 220787 297666
rect 217948 297608 220726 297664
rect 220782 297608 220787 297664
rect 217948 297606 220787 297608
rect 109910 297432 109970 297606
rect 111793 297603 111859 297606
rect 220721 297603 220787 297606
rect 154573 297530 154639 297533
rect 154573 297528 158148 297530
rect 154573 297472 154578 297528
rect 154634 297472 158148 297528
rect 154573 297470 158148 297472
rect 154573 297467 154639 297470
rect 111885 297258 111951 297261
rect 109910 297256 111951 297258
rect 109910 297200 111890 297256
rect 111946 297200 111951 297256
rect 109910 297198 111951 297200
rect 109910 296752 109970 297198
rect 111885 297195 111951 297198
rect 155033 297258 155099 297261
rect 220721 297258 220787 297261
rect 155033 297256 158148 297258
rect 155033 297200 155038 297256
rect 155094 297200 158148 297256
rect 155033 297198 158148 297200
rect 217948 297256 220787 297258
rect 217948 297200 220726 297256
rect 220782 297200 220787 297256
rect 217948 297198 220787 297200
rect 155033 297195 155099 297198
rect 220721 297195 220787 297198
rect 155493 296986 155559 296989
rect 155493 296984 158148 296986
rect 155493 296928 155498 296984
rect 155554 296928 158148 296984
rect 155493 296926 158148 296928
rect 155493 296923 155559 296926
rect 220353 296850 220419 296853
rect 217948 296848 220419 296850
rect 217948 296792 220358 296848
rect 220414 296792 220419 296848
rect 217948 296790 220419 296792
rect 220353 296787 220419 296790
rect 154849 296714 154915 296717
rect 154849 296712 158148 296714
rect 154849 296656 154854 296712
rect 154910 296656 158148 296712
rect 154849 296654 158148 296656
rect 154849 296651 154915 296654
rect 111793 296442 111859 296445
rect 109910 296440 111859 296442
rect 109910 296384 111798 296440
rect 111854 296384 111859 296440
rect 109910 296382 111859 296384
rect 109910 296072 109970 296382
rect 111793 296379 111859 296382
rect 154941 296442 155007 296445
rect 220629 296442 220695 296445
rect 154941 296440 158148 296442
rect 154941 296384 154946 296440
rect 155002 296384 158148 296440
rect 154941 296382 158148 296384
rect 217948 296440 220695 296442
rect 217948 296384 220634 296440
rect 220690 296384 220695 296440
rect 217948 296382 220695 296384
rect 154941 296379 155007 296382
rect 220629 296379 220695 296382
rect 256693 296306 256759 296309
rect 256693 296304 260084 296306
rect 256693 296248 256698 296304
rect 256754 296248 260084 296304
rect 256693 296246 260084 296248
rect 256693 296243 256759 296246
rect 154757 296170 154823 296173
rect 154757 296168 158148 296170
rect 154757 296112 154762 296168
rect 154818 296112 158148 296168
rect 154757 296110 158148 296112
rect 154757 296107 154823 296110
rect 219893 296034 219959 296037
rect 217948 296032 219959 296034
rect 217948 295976 219898 296032
rect 219954 295976 219959 296032
rect 217948 295974 219959 295976
rect 219893 295971 219959 295974
rect 111885 295898 111951 295901
rect 109910 295896 111951 295898
rect 109910 295840 111890 295896
rect 111946 295840 111951 295896
rect 109910 295838 111951 295840
rect 109910 295392 109970 295838
rect 111885 295835 111951 295838
rect 154665 295898 154731 295901
rect 154665 295896 158148 295898
rect 154665 295840 154670 295896
rect 154726 295840 158148 295896
rect 154665 295838 158148 295840
rect 154665 295835 154731 295838
rect 154573 295626 154639 295629
rect 220721 295626 220787 295629
rect 154573 295624 158148 295626
rect 154573 295568 154578 295624
rect 154634 295568 158148 295624
rect 154573 295566 158148 295568
rect 217948 295624 220787 295626
rect 217948 295568 220726 295624
rect 220782 295568 220787 295624
rect 217948 295566 220787 295568
rect 154573 295563 154639 295566
rect 220721 295563 220787 295566
rect 155401 295354 155467 295357
rect 155401 295352 158148 295354
rect 155401 295296 155406 295352
rect 155462 295296 158148 295352
rect 155401 295294 158148 295296
rect 155401 295291 155467 295294
rect 220261 295218 220327 295221
rect 217948 295216 220327 295218
rect 217948 295160 220266 295216
rect 220322 295160 220327 295216
rect 217948 295158 220327 295160
rect 220261 295155 220327 295158
rect 154757 295082 154823 295085
rect 154757 295080 158148 295082
rect 154757 295024 154762 295080
rect 154818 295024 158148 295080
rect 154757 295022 158148 295024
rect 154757 295019 154823 295022
rect 111793 294946 111859 294949
rect 109910 294944 111859 294946
rect 109910 294888 111798 294944
rect 111854 294888 111859 294944
rect 109910 294886 111859 294888
rect 109910 294712 109970 294886
rect 111793 294883 111859 294886
rect 154665 294810 154731 294813
rect 219893 294810 219959 294813
rect 154665 294808 158148 294810
rect 154665 294752 154670 294808
rect 154726 294752 158148 294808
rect 154665 294750 158148 294752
rect 217948 294808 219959 294810
rect 217948 294752 219898 294808
rect 219954 294752 219959 294808
rect 217948 294750 219959 294752
rect 154665 294747 154731 294750
rect 219893 294747 219959 294750
rect 111885 294538 111951 294541
rect 109910 294536 111951 294538
rect 109910 294480 111890 294536
rect 111946 294480 111951 294536
rect 109910 294478 111951 294480
rect 109910 294032 109970 294478
rect 111885 294475 111951 294478
rect 154849 294538 154915 294541
rect 154849 294536 158148 294538
rect 154849 294480 154854 294536
rect 154910 294480 158148 294536
rect 154849 294478 158148 294480
rect 154849 294475 154915 294478
rect 220721 294402 220787 294405
rect 217948 294400 220787 294402
rect 217948 294344 220726 294400
rect 220782 294344 220787 294400
rect 217948 294342 220787 294344
rect 220721 294339 220787 294342
rect 154573 294266 154639 294269
rect 256693 294266 256759 294269
rect 154573 294264 158148 294266
rect 154573 294208 154578 294264
rect 154634 294208 158148 294264
rect 154573 294206 158148 294208
rect 256693 294264 260084 294266
rect 256693 294208 256698 294264
rect 256754 294208 260084 294264
rect 256693 294206 260084 294208
rect 154573 294203 154639 294206
rect 256693 294203 256759 294206
rect 154573 293994 154639 293997
rect 220445 293994 220511 293997
rect 154573 293992 158148 293994
rect 154573 293936 154578 293992
rect 154634 293936 158148 293992
rect 154573 293934 158148 293936
rect 217948 293992 220511 293994
rect 217948 293936 220450 293992
rect 220506 293936 220511 293992
rect 217948 293934 220511 293936
rect 154573 293931 154639 293934
rect 220445 293931 220511 293934
rect 111793 293722 111859 293725
rect 109910 293720 111859 293722
rect 109910 293664 111798 293720
rect 111854 293664 111859 293720
rect 109910 293662 111859 293664
rect 109910 293352 109970 293662
rect 111793 293659 111859 293662
rect 154573 293722 154639 293725
rect 154573 293720 158148 293722
rect 154573 293664 154578 293720
rect 154634 293664 158148 293720
rect 154573 293662 158148 293664
rect 154573 293659 154639 293662
rect 220629 293586 220695 293589
rect 217948 293584 220695 293586
rect 217948 293528 220634 293584
rect 220690 293528 220695 293584
rect 217948 293526 220695 293528
rect 220629 293523 220695 293526
rect 154665 293450 154731 293453
rect 154665 293448 158148 293450
rect 154665 293392 154670 293448
rect 154726 293392 158148 293448
rect 154665 293390 158148 293392
rect 154665 293387 154731 293390
rect -960 293178 480 293268
rect 3417 293178 3483 293181
rect 111885 293178 111951 293181
rect -960 293176 3483 293178
rect -960 293120 3422 293176
rect 3478 293120 3483 293176
rect -960 293118 3483 293120
rect -960 293028 480 293118
rect 3417 293115 3483 293118
rect 109910 293176 111951 293178
rect 109910 293120 111890 293176
rect 111946 293120 111951 293176
rect 109910 293118 111951 293120
rect 109910 292672 109970 293118
rect 111885 293115 111951 293118
rect 155350 293116 155356 293180
rect 155420 293178 155426 293180
rect 220721 293178 220787 293181
rect 155420 293118 158148 293178
rect 217948 293176 220787 293178
rect 217948 293120 220726 293176
rect 220782 293120 220787 293176
rect 217948 293118 220787 293120
rect 155420 293116 155426 293118
rect 220721 293115 220787 293118
rect 155217 292906 155283 292909
rect 155217 292904 158148 292906
rect 155217 292848 155222 292904
rect 155278 292848 158148 292904
rect 155217 292846 158148 292848
rect 155217 292843 155283 292846
rect 220537 292770 220603 292773
rect 217948 292768 220603 292770
rect 217948 292712 220542 292768
rect 220598 292712 220603 292768
rect 217948 292710 220603 292712
rect 220537 292707 220603 292710
rect 154573 292634 154639 292637
rect 154573 292632 158148 292634
rect 154573 292576 154578 292632
rect 154634 292576 158148 292632
rect 154573 292574 158148 292576
rect 154573 292571 154639 292574
rect 155309 292362 155375 292365
rect 219893 292362 219959 292365
rect 155309 292360 158148 292362
rect 155309 292304 155314 292360
rect 155370 292304 158148 292360
rect 155309 292302 158148 292304
rect 217948 292360 219959 292362
rect 217948 292304 219898 292360
rect 219954 292304 219959 292360
rect 217948 292302 219959 292304
rect 155309 292299 155375 292302
rect 219893 292299 219959 292302
rect 111793 292226 111859 292229
rect 109910 292224 111859 292226
rect 109910 292168 111798 292224
rect 111854 292168 111859 292224
rect 109910 292166 111859 292168
rect 109910 291992 109970 292166
rect 111793 292163 111859 292166
rect 256693 292226 256759 292229
rect 256693 292224 260084 292226
rect 256693 292168 256698 292224
rect 256754 292168 260084 292224
rect 256693 292166 260084 292168
rect 256693 292163 256759 292166
rect 220629 291954 220695 291957
rect 217948 291952 220695 291954
rect 217948 291896 220634 291952
rect 220690 291896 220695 291952
rect 217948 291894 220695 291896
rect 220629 291891 220695 291894
rect 111885 291818 111951 291821
rect 109910 291816 111951 291818
rect 109910 291760 111890 291816
rect 111946 291760 111951 291816
rect 109910 291758 111951 291760
rect 109910 291312 109970 291758
rect 111885 291755 111951 291758
rect 220721 291546 220787 291549
rect 217948 291544 220787 291546
rect 217948 291488 220726 291544
rect 220782 291488 220787 291544
rect 217948 291486 220787 291488
rect 220721 291483 220787 291486
rect 220721 291138 220787 291141
rect 217948 291136 220787 291138
rect 217948 291080 220726 291136
rect 220782 291080 220787 291136
rect 217948 291078 220787 291080
rect 220721 291075 220787 291078
rect 111793 290866 111859 290869
rect 109910 290864 111859 290866
rect 109910 290808 111798 290864
rect 111854 290808 111859 290864
rect 109910 290806 111859 290808
rect 109910 290632 109970 290806
rect 111793 290803 111859 290806
rect 220629 290730 220695 290733
rect 217948 290728 220695 290730
rect 217948 290672 220634 290728
rect 220690 290672 220695 290728
rect 217948 290670 220695 290672
rect 220629 290667 220695 290670
rect 111885 290458 111951 290461
rect 109910 290456 111951 290458
rect 109910 290400 111890 290456
rect 111946 290400 111951 290456
rect 109910 290398 111951 290400
rect 109910 289952 109970 290398
rect 111885 290395 111951 290398
rect 220261 290322 220327 290325
rect 217948 290320 220327 290322
rect 217948 290264 220266 290320
rect 220322 290264 220327 290320
rect 217948 290262 220327 290264
rect 220261 290259 220327 290262
rect 256693 290186 256759 290189
rect 256693 290184 260084 290186
rect 256693 290128 256698 290184
rect 256754 290128 260084 290184
rect 256693 290126 260084 290128
rect 256693 290123 256759 290126
rect 220721 289914 220787 289917
rect 217948 289912 220787 289914
rect 217948 289856 220726 289912
rect 220782 289856 220787 289912
rect 217948 289854 220787 289856
rect 220721 289851 220787 289854
rect 111793 289506 111859 289509
rect 220537 289506 220603 289509
rect 109910 289504 111859 289506
rect 109910 289448 111798 289504
rect 111854 289448 111859 289504
rect 109910 289446 111859 289448
rect 217948 289504 220603 289506
rect 217948 289448 220542 289504
rect 220598 289448 220603 289504
rect 217948 289446 220603 289448
rect 109910 289272 109970 289446
rect 111793 289443 111859 289446
rect 220537 289443 220603 289446
rect 111885 289098 111951 289101
rect 220629 289098 220695 289101
rect 109910 289096 111951 289098
rect 109910 289040 111890 289096
rect 111946 289040 111951 289096
rect 109910 289038 111951 289040
rect 217948 289096 220695 289098
rect 217948 289040 220634 289096
rect 220690 289040 220695 289096
rect 217948 289038 220695 289040
rect 109910 288592 109970 289038
rect 111885 289035 111951 289038
rect 220629 289035 220695 289038
rect 220721 288690 220787 288693
rect 217948 288688 220787 288690
rect 217948 288632 220726 288688
rect 220782 288632 220787 288688
rect 217948 288630 220787 288632
rect 220721 288627 220787 288630
rect 219525 288282 219591 288285
rect 217948 288280 219591 288282
rect 217948 288224 219530 288280
rect 219586 288224 219591 288280
rect 217948 288222 219591 288224
rect 219525 288219 219591 288222
rect 111793 288146 111859 288149
rect 109910 288144 111859 288146
rect 109910 288088 111798 288144
rect 111854 288088 111859 288144
rect 109910 288086 111859 288088
rect 109910 287912 109970 288086
rect 111793 288083 111859 288086
rect 256693 288146 256759 288149
rect 256693 288144 260084 288146
rect 256693 288088 256698 288144
rect 256754 288088 260084 288144
rect 256693 288086 260084 288088
rect 256693 288083 256759 288086
rect 220629 287874 220695 287877
rect 217948 287872 220695 287874
rect 217948 287816 220634 287872
rect 220690 287816 220695 287872
rect 217948 287814 220695 287816
rect 220629 287811 220695 287814
rect 111885 287738 111951 287741
rect 109910 287736 111951 287738
rect 109910 287680 111890 287736
rect 111946 287680 111951 287736
rect 109910 287678 111951 287680
rect 109910 287232 109970 287678
rect 111885 287675 111951 287678
rect 220721 287466 220787 287469
rect 217948 287464 220787 287466
rect 217948 287408 220726 287464
rect 220782 287408 220787 287464
rect 217948 287406 220787 287408
rect 220721 287403 220787 287406
rect 219893 287058 219959 287061
rect 217948 287056 219959 287058
rect 217948 287000 219898 287056
rect 219954 287000 219959 287056
rect 217948 286998 219959 287000
rect 219893 286995 219959 286998
rect 111793 286786 111859 286789
rect 109910 286784 111859 286786
rect 109910 286728 111798 286784
rect 111854 286728 111859 286784
rect 109910 286726 111859 286728
rect 109910 286552 109970 286726
rect 111793 286723 111859 286726
rect 219893 286650 219959 286653
rect 217948 286648 219959 286650
rect 217948 286592 219898 286648
rect 219954 286592 219959 286648
rect 217948 286590 219959 286592
rect 219893 286587 219959 286590
rect 111885 286378 111951 286381
rect 109910 286376 111951 286378
rect 109910 286320 111890 286376
rect 111946 286320 111951 286376
rect 109910 286318 111951 286320
rect 109910 285872 109970 286318
rect 111885 286315 111951 286318
rect 220629 286242 220695 286245
rect 217948 286240 220695 286242
rect 217948 286184 220634 286240
rect 220690 286184 220695 286240
rect 217948 286182 220695 286184
rect 220629 286179 220695 286182
rect 257337 286106 257403 286109
rect 257337 286104 260084 286106
rect 257337 286048 257342 286104
rect 257398 286048 260084 286104
rect 257337 286046 260084 286048
rect 257337 286043 257403 286046
rect 220721 285834 220787 285837
rect 217948 285832 220787 285834
rect 217948 285776 220726 285832
rect 220782 285776 220787 285832
rect 217948 285774 220787 285776
rect 220721 285771 220787 285774
rect 111793 285426 111859 285429
rect 109910 285424 111859 285426
rect 109910 285368 111798 285424
rect 111854 285368 111859 285424
rect 109910 285366 111859 285368
rect 109910 285192 109970 285366
rect 111793 285363 111859 285366
rect 583520 285276 584960 285516
rect 111885 285018 111951 285021
rect 109910 285016 111951 285018
rect 109910 284960 111890 285016
rect 111946 284960 111951 285016
rect 109910 284958 111951 284960
rect 109910 284512 109970 284958
rect 111885 284955 111951 284958
rect 111793 284066 111859 284069
rect 109910 284064 111859 284066
rect 109910 284008 111798 284064
rect 111854 284008 111859 284064
rect 109910 284006 111859 284008
rect 109910 283832 109970 284006
rect 111793 284003 111859 284006
rect 257613 284066 257679 284069
rect 257613 284064 260084 284066
rect 257613 284008 257618 284064
rect 257674 284008 260084 284064
rect 257613 284006 260084 284008
rect 257613 284003 257679 284006
rect 111885 283658 111951 283661
rect 109910 283656 111951 283658
rect 109910 283600 111890 283656
rect 111946 283600 111951 283656
rect 109910 283598 111951 283600
rect 109910 283152 109970 283598
rect 111885 283595 111951 283598
rect 112069 282842 112135 282845
rect 109910 282840 112135 282842
rect 109910 282784 112074 282840
rect 112130 282784 112135 282840
rect 109910 282782 112135 282784
rect 109910 282472 109970 282782
rect 112069 282779 112135 282782
rect 111793 282298 111859 282301
rect 109910 282296 111859 282298
rect 109910 282240 111798 282296
rect 111854 282240 111859 282296
rect 109910 282238 111859 282240
rect 109910 281792 109970 282238
rect 111793 282235 111859 282238
rect 256693 282026 256759 282029
rect 256693 282024 260084 282026
rect 256693 281968 256698 282024
rect 256754 281968 260084 282024
rect 256693 281966 260084 281968
rect 256693 281963 256759 281966
rect 111793 281346 111859 281349
rect 109910 281344 111859 281346
rect 109910 281288 111798 281344
rect 111854 281288 111859 281344
rect 109910 281286 111859 281288
rect 109910 281112 109970 281286
rect 111793 281283 111859 281286
rect 111885 280938 111951 280941
rect 109910 280936 111951 280938
rect 109910 280880 111890 280936
rect 111946 280880 111951 280936
rect 109910 280878 111951 280880
rect 109910 280432 109970 280878
rect 111885 280875 111951 280878
rect -960 279972 480 280212
rect 111793 279986 111859 279989
rect 109910 279984 111859 279986
rect 109910 279928 111798 279984
rect 111854 279928 111859 279984
rect 109910 279926 111859 279928
rect 109910 279752 109970 279926
rect 111793 279923 111859 279926
rect 256693 279986 256759 279989
rect 256693 279984 260084 279986
rect 256693 279928 256698 279984
rect 256754 279928 260084 279984
rect 256693 279926 260084 279928
rect 256693 279923 256759 279926
rect 111885 279578 111951 279581
rect 109910 279576 111951 279578
rect 109910 279520 111890 279576
rect 111946 279520 111951 279576
rect 109910 279518 111951 279520
rect 109910 279072 109970 279518
rect 111885 279515 111951 279518
rect 111793 278490 111859 278493
rect 109910 278488 111859 278490
rect 109910 278432 111798 278488
rect 111854 278432 111859 278488
rect 109910 278430 111859 278432
rect 109910 278392 109970 278430
rect 111793 278427 111859 278430
rect 111885 278218 111951 278221
rect 109910 278216 111951 278218
rect 109910 278160 111890 278216
rect 111946 278160 111951 278216
rect 109910 278158 111951 278160
rect 109910 277712 109970 278158
rect 111885 278155 111951 278158
rect 256693 277946 256759 277949
rect 256693 277944 260084 277946
rect 256693 277888 256698 277944
rect 256754 277888 260084 277944
rect 256693 277886 260084 277888
rect 256693 277883 256759 277886
rect 111793 277266 111859 277269
rect 109910 277264 111859 277266
rect 109910 277208 111798 277264
rect 111854 277208 111859 277264
rect 109910 277206 111859 277208
rect 109910 277032 109970 277206
rect 111793 277203 111859 277206
rect 111885 276858 111951 276861
rect 109910 276856 111951 276858
rect 109910 276800 111890 276856
rect 111946 276800 111951 276856
rect 109910 276798 111951 276800
rect 109910 276352 109970 276798
rect 111885 276795 111951 276798
rect 111793 275906 111859 275909
rect 109910 275904 111859 275906
rect 109910 275848 111798 275904
rect 111854 275848 111859 275904
rect 109910 275846 111859 275848
rect 109910 275672 109970 275846
rect 111793 275843 111859 275846
rect 256693 275906 256759 275909
rect 256693 275904 260084 275906
rect 256693 275848 256698 275904
rect 256754 275848 260084 275904
rect 256693 275846 260084 275848
rect 256693 275843 256759 275846
rect 111885 275498 111951 275501
rect 109910 275496 111951 275498
rect 109910 275440 111890 275496
rect 111946 275440 111951 275496
rect 109910 275438 111951 275440
rect 109910 274992 109970 275438
rect 111885 275435 111951 275438
rect 111793 274410 111859 274413
rect 109910 274408 111859 274410
rect 109910 274352 111798 274408
rect 111854 274352 111859 274408
rect 109910 274350 111859 274352
rect 109910 274312 109970 274350
rect 111793 274347 111859 274350
rect 111885 274138 111951 274141
rect 109910 274136 111951 274138
rect 109910 274080 111890 274136
rect 111946 274080 111951 274136
rect 109910 274078 111951 274080
rect 109910 273632 109970 274078
rect 111885 274075 111951 274078
rect 256693 273866 256759 273869
rect 256693 273864 260084 273866
rect 256693 273808 256698 273864
rect 256754 273808 260084 273864
rect 256693 273806 260084 273808
rect 256693 273803 256759 273806
rect 111793 273050 111859 273053
rect 109910 273048 111859 273050
rect 109910 272992 111798 273048
rect 111854 272992 111859 273048
rect 109910 272990 111859 272992
rect 109910 272952 109970 272990
rect 111793 272987 111859 272990
rect 111885 272778 111951 272781
rect 109910 272776 111951 272778
rect 109910 272720 111890 272776
rect 111946 272720 111951 272776
rect 109910 272718 111951 272720
rect 109910 272272 109970 272718
rect 111885 272715 111951 272718
rect 580165 272234 580231 272237
rect 583520 272234 584960 272324
rect 580165 272232 584960 272234
rect 580165 272176 580170 272232
rect 580226 272176 584960 272232
rect 580165 272174 584960 272176
rect 580165 272171 580231 272174
rect 583520 272084 584960 272174
rect 257429 271826 257495 271829
rect 257429 271824 260084 271826
rect 257429 271768 257434 271824
rect 257490 271768 260084 271824
rect 257429 271766 260084 271768
rect 257429 271763 257495 271766
rect 111793 271690 111859 271693
rect 109910 271688 111859 271690
rect 109910 271632 111798 271688
rect 111854 271632 111859 271688
rect 109910 271630 111859 271632
rect 109910 271592 109970 271630
rect 111793 271627 111859 271630
rect 111885 271418 111951 271421
rect 109910 271416 111951 271418
rect 109910 271360 111890 271416
rect 111946 271360 111951 271416
rect 109910 271358 111951 271360
rect 109910 270912 109970 271358
rect 111885 271355 111951 271358
rect 111793 270330 111859 270333
rect 109910 270328 111859 270330
rect 109910 270272 111798 270328
rect 111854 270272 111859 270328
rect 109910 270270 111859 270272
rect 109910 270232 109970 270270
rect 111793 270267 111859 270270
rect 111885 270058 111951 270061
rect 109910 270056 111951 270058
rect 109910 270000 111890 270056
rect 111946 270000 111951 270056
rect 109910 269998 111951 270000
rect 109910 269552 109970 269998
rect 111885 269995 111951 269998
rect 256693 269786 256759 269789
rect 256693 269784 260084 269786
rect 256693 269728 256698 269784
rect 256754 269728 260084 269784
rect 256693 269726 260084 269728
rect 256693 269723 256759 269726
rect 111793 268970 111859 268973
rect 109910 268968 111859 268970
rect 109910 268912 111798 268968
rect 111854 268912 111859 268968
rect 109910 268910 111859 268912
rect 109910 268872 109970 268910
rect 111793 268907 111859 268910
rect 111885 268698 111951 268701
rect 109910 268696 111951 268698
rect 109910 268640 111890 268696
rect 111946 268640 111951 268696
rect 109910 268638 111951 268640
rect 109910 268192 109970 268638
rect 111885 268635 111951 268638
rect 257797 267746 257863 267749
rect 257797 267744 260084 267746
rect 257797 267688 257802 267744
rect 257858 267688 260084 267744
rect 257797 267686 260084 267688
rect 257797 267683 257863 267686
rect 111793 267610 111859 267613
rect 109910 267608 111859 267610
rect 109910 267552 111798 267608
rect 111854 267552 111859 267608
rect 109910 267550 111859 267552
rect 109910 267512 109970 267550
rect 111793 267547 111859 267550
rect -960 267202 480 267292
rect 3049 267202 3115 267205
rect 111885 267202 111951 267205
rect -960 267200 3115 267202
rect -960 267144 3054 267200
rect 3110 267144 3115 267200
rect -960 267142 3115 267144
rect -960 267052 480 267142
rect 3049 267139 3115 267142
rect 109910 267200 111951 267202
rect 109910 267144 111890 267200
rect 111946 267144 111951 267200
rect 109910 267142 111951 267144
rect 109910 266832 109970 267142
rect 111885 267139 111951 267142
rect 111793 266250 111859 266253
rect 109910 266248 111859 266250
rect 109910 266192 111798 266248
rect 111854 266192 111859 266248
rect 109910 266190 111859 266192
rect 109910 266152 109970 266190
rect 111793 266187 111859 266190
rect 111885 265978 111951 265981
rect 109910 265976 111951 265978
rect 109910 265920 111890 265976
rect 111946 265920 111951 265976
rect 109910 265918 111951 265920
rect 109910 265472 109970 265918
rect 111885 265915 111951 265918
rect 256693 265706 256759 265709
rect 256693 265704 260084 265706
rect 256693 265648 256698 265704
rect 256754 265648 260084 265704
rect 256693 265646 260084 265648
rect 256693 265643 256759 265646
rect 111793 264890 111859 264893
rect 109910 264888 111859 264890
rect 109910 264832 111798 264888
rect 111854 264832 111859 264888
rect 109910 264830 111859 264832
rect 109910 264792 109970 264830
rect 111793 264827 111859 264830
rect 111885 264482 111951 264485
rect 109910 264480 111951 264482
rect 109910 264424 111890 264480
rect 111946 264424 111951 264480
rect 109910 264422 111951 264424
rect 109910 264112 109970 264422
rect 111885 264419 111951 264422
rect 256693 263666 256759 263669
rect 256693 263664 260084 263666
rect 256693 263608 256698 263664
rect 256754 263608 260084 263664
rect 256693 263606 260084 263608
rect 256693 263603 256759 263606
rect 111793 263530 111859 263533
rect 109910 263528 111859 263530
rect 109910 263472 111798 263528
rect 111854 263472 111859 263528
rect 109910 263470 111859 263472
rect 109910 263432 109970 263470
rect 111793 263467 111859 263470
rect 111885 263122 111951 263125
rect 109910 263120 111951 263122
rect 109910 263064 111890 263120
rect 111946 263064 111951 263120
rect 109910 263062 111951 263064
rect 109910 262752 109970 263062
rect 111885 263059 111951 263062
rect 112161 262170 112227 262173
rect 109910 262168 112227 262170
rect 109910 262112 112166 262168
rect 112222 262112 112227 262168
rect 109910 262110 112227 262112
rect 109910 262072 109970 262110
rect 112161 262107 112227 262110
rect 111793 261762 111859 261765
rect 109910 261760 111859 261762
rect 109910 261704 111798 261760
rect 111854 261704 111859 261760
rect 109910 261702 111859 261704
rect 109910 261392 109970 261702
rect 111793 261699 111859 261702
rect 256693 261626 256759 261629
rect 256693 261624 260084 261626
rect 256693 261568 256698 261624
rect 256754 261568 260084 261624
rect 256693 261566 260084 261568
rect 256693 261563 256759 261566
rect 112989 261082 113055 261085
rect 112989 261080 113098 261082
rect 112989 261024 112994 261080
rect 113050 261024 113098 261080
rect 112989 261019 113098 261024
rect 111793 260810 111859 260813
rect 109910 260808 111859 260810
rect 109910 260752 111798 260808
rect 111854 260752 111859 260808
rect 109910 260750 111859 260752
rect 109910 260712 109970 260750
rect 111793 260747 111859 260750
rect 113038 260541 113098 261019
rect 112989 260536 113098 260541
rect 112989 260480 112994 260536
rect 113050 260480 113098 260536
rect 112989 260478 113098 260480
rect 112989 260475 113055 260478
rect 111885 260402 111951 260405
rect 109910 260400 111951 260402
rect 109910 260344 111890 260400
rect 111946 260344 111951 260400
rect 109910 260342 111951 260344
rect 109910 260032 109970 260342
rect 111885 260339 111951 260342
rect 256693 259586 256759 259589
rect 256693 259584 260084 259586
rect 256693 259528 256698 259584
rect 256754 259528 260084 259584
rect 256693 259526 260084 259528
rect 256693 259523 256759 259526
rect 109910 259314 109970 259352
rect 111793 259314 111859 259317
rect 109910 259312 111859 259314
rect 109910 259256 111798 259312
rect 111854 259256 111859 259312
rect 109910 259254 111859 259256
rect 111793 259251 111859 259254
rect 111885 259042 111951 259045
rect 109910 259040 111951 259042
rect 109910 258984 111890 259040
rect 111946 258984 111951 259040
rect 109910 258982 111951 258984
rect 109910 258672 109970 258982
rect 111885 258979 111951 258982
rect 580165 258906 580231 258909
rect 583520 258906 584960 258996
rect 580165 258904 584960 258906
rect 580165 258848 580170 258904
rect 580226 258848 584960 258904
rect 580165 258846 584960 258848
rect 580165 258843 580231 258846
rect 583520 258756 584960 258846
rect 109910 257954 109970 257992
rect 111793 257954 111859 257957
rect 109910 257952 111859 257954
rect 109910 257896 111798 257952
rect 111854 257896 111859 257952
rect 109910 257894 111859 257896
rect 111793 257891 111859 257894
rect 111885 257682 111951 257685
rect 109910 257680 111951 257682
rect 109910 257624 111890 257680
rect 111946 257624 111951 257680
rect 109910 257622 111951 257624
rect 109910 257312 109970 257622
rect 111885 257619 111951 257622
rect 256693 257546 256759 257549
rect 256693 257544 260084 257546
rect 256693 257488 256698 257544
rect 256754 257488 260084 257544
rect 256693 257486 260084 257488
rect 256693 257483 256759 257486
rect 109910 256594 109970 256632
rect 113081 256594 113147 256597
rect 109910 256592 113147 256594
rect 109910 256536 113086 256592
rect 113142 256536 113147 256592
rect 109910 256534 113147 256536
rect 113081 256531 113147 256534
rect 111793 256322 111859 256325
rect 109910 256320 111859 256322
rect 109910 256264 111798 256320
rect 111854 256264 111859 256320
rect 109910 256262 111859 256264
rect 109910 255952 109970 256262
rect 111793 256259 111859 256262
rect 256693 255506 256759 255509
rect 256693 255504 260084 255506
rect 256693 255448 256698 255504
rect 256754 255448 260084 255504
rect 256693 255446 260084 255448
rect 256693 255443 256759 255446
rect 109910 255234 109970 255272
rect 112989 255234 113055 255237
rect 109910 255232 113055 255234
rect 109910 255176 112994 255232
rect 113050 255176 113055 255232
rect 109910 255174 113055 255176
rect 112989 255171 113055 255174
rect 111793 254962 111859 254965
rect 109910 254960 111859 254962
rect 109910 254904 111798 254960
rect 111854 254904 111859 254960
rect 109910 254902 111859 254904
rect 109910 254592 109970 254902
rect 111793 254899 111859 254902
rect -960 254146 480 254236
rect 3509 254146 3575 254149
rect -960 254144 3575 254146
rect -960 254088 3514 254144
rect 3570 254088 3575 254144
rect -960 254086 3575 254088
rect -960 253996 480 254086
rect 3509 254083 3575 254086
rect 109910 253874 109970 253912
rect 111793 253874 111859 253877
rect 109910 253872 111859 253874
rect 109910 253816 111798 253872
rect 111854 253816 111859 253872
rect 109910 253814 111859 253816
rect 111793 253811 111859 253814
rect 111885 253602 111951 253605
rect 109910 253600 111951 253602
rect 109910 253544 111890 253600
rect 111946 253544 111951 253600
rect 109910 253542 111951 253544
rect 109910 253232 109970 253542
rect 111885 253539 111951 253542
rect 256693 253466 256759 253469
rect 256693 253464 260084 253466
rect 256693 253408 256698 253464
rect 256754 253408 260084 253464
rect 256693 253406 260084 253408
rect 256693 253403 256759 253406
rect 111793 253058 111859 253061
rect 109910 253056 111859 253058
rect 109910 253000 111798 253056
rect 111854 253000 111859 253056
rect 109910 252998 111859 253000
rect 109910 252552 109970 252998
rect 111793 252995 111859 252998
rect 111793 252242 111859 252245
rect 109910 252240 111859 252242
rect 109910 252184 111798 252240
rect 111854 252184 111859 252240
rect 109910 252182 111859 252184
rect 109910 251872 109970 252182
rect 111793 252179 111859 252182
rect 112253 251698 112319 251701
rect 109910 251696 112319 251698
rect 109910 251640 112258 251696
rect 112314 251640 112319 251696
rect 109910 251638 112319 251640
rect 109910 251192 109970 251638
rect 112253 251635 112319 251638
rect 256693 251426 256759 251429
rect 256693 251424 260084 251426
rect 256693 251368 256698 251424
rect 256754 251368 260084 251424
rect 256693 251366 260084 251368
rect 256693 251363 256759 251366
rect 111793 250882 111859 250885
rect 109910 250880 111859 250882
rect 109910 250824 111798 250880
rect 111854 250824 111859 250880
rect 109910 250822 111859 250824
rect 109910 250512 109970 250822
rect 111793 250819 111859 250822
rect 111885 250338 111951 250341
rect 109910 250336 111951 250338
rect 109910 250280 111890 250336
rect 111946 250280 111951 250336
rect 109910 250278 111951 250280
rect 109910 249832 109970 250278
rect 111885 250275 111951 250278
rect 111793 249522 111859 249525
rect 109910 249520 111859 249522
rect 109910 249464 111798 249520
rect 111854 249464 111859 249520
rect 109910 249462 111859 249464
rect 109910 249152 109970 249462
rect 111793 249459 111859 249462
rect 256693 249386 256759 249389
rect 256693 249384 260084 249386
rect 256693 249328 256698 249384
rect 256754 249328 260084 249384
rect 256693 249326 260084 249328
rect 256693 249323 256759 249326
rect 112805 248978 112871 248981
rect 109910 248976 112871 248978
rect 109910 248920 112810 248976
rect 112866 248920 112871 248976
rect 109910 248918 112871 248920
rect 109910 248472 109970 248918
rect 112805 248915 112871 248918
rect 111793 248026 111859 248029
rect 109910 248024 111859 248026
rect 109910 247968 111798 248024
rect 111854 247968 111859 248024
rect 109910 247966 111859 247968
rect 109910 247792 109970 247966
rect 111793 247963 111859 247966
rect 111885 247618 111951 247621
rect 109910 247616 111951 247618
rect 109910 247560 111890 247616
rect 111946 247560 111951 247616
rect 109910 247558 111951 247560
rect 109910 247112 109970 247558
rect 111885 247555 111951 247558
rect 256693 247346 256759 247349
rect 256693 247344 260084 247346
rect 256693 247288 256698 247344
rect 256754 247288 260084 247344
rect 256693 247286 260084 247288
rect 256693 247283 256759 247286
rect 111793 246666 111859 246669
rect 109910 246664 111859 246666
rect 109910 246608 111798 246664
rect 111854 246608 111859 246664
rect 109910 246606 111859 246608
rect 109910 246432 109970 246606
rect 111793 246603 111859 246606
rect 111885 246258 111951 246261
rect 109910 246256 111951 246258
rect 109910 246200 111890 246256
rect 111946 246200 111951 246256
rect 109910 246198 111951 246200
rect 109910 245752 109970 246198
rect 111885 246195 111951 246198
rect 580349 245578 580415 245581
rect 583520 245578 584960 245668
rect 580349 245576 584960 245578
rect 580349 245520 580354 245576
rect 580410 245520 584960 245576
rect 580349 245518 584960 245520
rect 580349 245515 580415 245518
rect 583520 245428 584960 245518
rect 111793 245306 111859 245309
rect 109910 245304 111859 245306
rect 109910 245248 111798 245304
rect 111854 245248 111859 245304
rect 109910 245246 111859 245248
rect 109910 245072 109970 245246
rect 111793 245243 111859 245246
rect 256693 245306 256759 245309
rect 256693 245304 260084 245306
rect 256693 245248 256698 245304
rect 256754 245248 260084 245304
rect 256693 245246 260084 245248
rect 256693 245243 256759 245246
rect 111885 244898 111951 244901
rect 109910 244896 111951 244898
rect 109910 244840 111890 244896
rect 111946 244840 111951 244896
rect 109910 244838 111951 244840
rect 109910 244392 109970 244838
rect 111885 244835 111951 244838
rect 111793 243946 111859 243949
rect 109910 243944 111859 243946
rect 109910 243888 111798 243944
rect 111854 243888 111859 243944
rect 109910 243886 111859 243888
rect 109910 243712 109970 243886
rect 111793 243883 111859 243886
rect 112345 243538 112411 243541
rect 109910 243536 112411 243538
rect 109910 243480 112350 243536
rect 112406 243480 112411 243536
rect 109910 243478 112411 243480
rect 109910 243032 109970 243478
rect 112345 243475 112411 243478
rect 256693 243266 256759 243269
rect 256693 243264 260084 243266
rect 256693 243208 256698 243264
rect 256754 243208 260084 243264
rect 256693 243206 260084 243208
rect 256693 243203 256759 243206
rect 111793 242586 111859 242589
rect 109910 242584 111859 242586
rect 109910 242528 111798 242584
rect 111854 242528 111859 242584
rect 109910 242526 111859 242528
rect 109910 242352 109970 242526
rect 111793 242523 111859 242526
rect 111977 242178 112043 242181
rect 109910 242176 112043 242178
rect 109910 242120 111982 242176
rect 112038 242120 112043 242176
rect 109910 242118 112043 242120
rect 109910 241672 109970 242118
rect 111977 242115 112043 242118
rect 111885 241498 111951 241501
rect 109910 241496 111951 241498
rect 109910 241440 111890 241496
rect 111946 241440 111951 241496
rect 109910 241438 111951 241440
rect -960 241090 480 241180
rect 3509 241090 3575 241093
rect -960 241088 3575 241090
rect -960 241032 3514 241088
rect 3570 241032 3575 241088
rect -960 241030 3575 241032
rect -960 240940 480 241030
rect 3509 241027 3575 241030
rect 109910 240992 109970 241438
rect 111885 241435 111951 241438
rect 256693 241226 256759 241229
rect 256693 241224 260084 241226
rect 256693 241168 256698 241224
rect 256754 241168 260084 241224
rect 256693 241166 260084 241168
rect 256693 241163 256759 241166
rect 111793 240818 111859 240821
rect 109910 240816 111859 240818
rect 109910 240760 111798 240816
rect 111854 240760 111859 240816
rect 109910 240758 111859 240760
rect 109910 240312 109970 240758
rect 111793 240755 111859 240758
rect 111793 239866 111859 239869
rect 109910 239864 111859 239866
rect 109910 239808 111798 239864
rect 111854 239808 111859 239864
rect 109910 239806 111859 239808
rect 109910 239632 109970 239806
rect 111793 239803 111859 239806
rect 111885 239458 111951 239461
rect 109910 239456 111951 239458
rect 109910 239400 111890 239456
rect 111946 239400 111951 239456
rect 109910 239398 111951 239400
rect 109910 238952 109970 239398
rect 111885 239395 111951 239398
rect 256693 239186 256759 239189
rect 256693 239184 260084 239186
rect 256693 239128 256698 239184
rect 256754 239128 260084 239184
rect 256693 239126 260084 239128
rect 256693 239123 256759 239126
rect 111793 238506 111859 238509
rect 109910 238504 111859 238506
rect 109910 238448 111798 238504
rect 111854 238448 111859 238504
rect 109910 238446 111859 238448
rect 109910 238272 109970 238446
rect 111793 238443 111859 238446
rect 111885 238098 111951 238101
rect 109910 238096 111951 238098
rect 109910 238040 111890 238096
rect 111946 238040 111951 238096
rect 109910 238038 111951 238040
rect 109910 237592 109970 238038
rect 111885 238035 111951 238038
rect 111793 237146 111859 237149
rect 109910 237144 111859 237146
rect 109910 237088 111798 237144
rect 111854 237088 111859 237144
rect 109910 237086 111859 237088
rect 109910 236912 109970 237086
rect 111793 237083 111859 237086
rect 256693 237146 256759 237149
rect 256693 237144 260084 237146
rect 256693 237088 256698 237144
rect 256754 237088 260084 237144
rect 256693 237086 260084 237088
rect 256693 237083 256759 237086
rect 112345 236738 112411 236741
rect 109910 236736 112411 236738
rect 109910 236680 112350 236736
rect 112406 236680 112411 236736
rect 109910 236678 112411 236680
rect 109910 236232 109970 236678
rect 112345 236675 112411 236678
rect 111793 235786 111859 235789
rect 109910 235784 111859 235786
rect 109910 235728 111798 235784
rect 111854 235728 111859 235784
rect 109910 235726 111859 235728
rect 109910 235552 109970 235726
rect 111793 235723 111859 235726
rect 111885 235378 111951 235381
rect 109910 235376 111951 235378
rect 109910 235320 111890 235376
rect 111946 235320 111951 235376
rect 109910 235318 111951 235320
rect 109910 234872 109970 235318
rect 111885 235315 111951 235318
rect 257337 235106 257403 235109
rect 257337 235104 260084 235106
rect 257337 235048 257342 235104
rect 257398 235048 260084 235104
rect 257337 235046 260084 235048
rect 257337 235043 257403 235046
rect 111793 234426 111859 234429
rect 109910 234424 111859 234426
rect 109910 234368 111798 234424
rect 111854 234368 111859 234424
rect 109910 234366 111859 234368
rect 109910 234192 109970 234366
rect 111793 234363 111859 234366
rect 111885 234018 111951 234021
rect 109910 234016 111951 234018
rect 109910 233960 111890 234016
rect 111946 233960 111951 234016
rect 109910 233958 111951 233960
rect 109910 233512 109970 233958
rect 111885 233955 111951 233958
rect 111793 233202 111859 233205
rect 109910 233200 111859 233202
rect 109910 233144 111798 233200
rect 111854 233144 111859 233200
rect 109910 233142 111859 233144
rect 109910 232832 109970 233142
rect 111793 233139 111859 233142
rect 256693 233066 256759 233069
rect 256693 233064 260084 233066
rect 256693 233008 256698 233064
rect 256754 233008 260084 233064
rect 256693 233006 260084 233008
rect 256693 233003 256759 233006
rect 111793 232522 111859 232525
rect 109910 232520 111859 232522
rect 109910 232464 111798 232520
rect 111854 232464 111859 232520
rect 109910 232462 111859 232464
rect 109910 232152 109970 232462
rect 111793 232459 111859 232462
rect 579613 232386 579679 232389
rect 583520 232386 584960 232476
rect 579613 232384 584960 232386
rect 579613 232328 579618 232384
rect 579674 232328 584960 232384
rect 579613 232326 584960 232328
rect 579613 232323 579679 232326
rect 583520 232236 584960 232326
rect 112897 231842 112963 231845
rect 109910 231840 112963 231842
rect 109910 231784 112902 231840
rect 112958 231784 112963 231840
rect 109910 231782 112963 231784
rect 109910 231472 109970 231782
rect 112897 231779 112963 231782
rect 111793 231298 111859 231301
rect 109910 231296 111859 231298
rect 109910 231240 111798 231296
rect 111854 231240 111859 231296
rect 109910 231238 111859 231240
rect 109910 230792 109970 231238
rect 111793 231235 111859 231238
rect 256325 231026 256391 231029
rect 256325 231024 260084 231026
rect 256325 230968 256330 231024
rect 256386 230968 260084 231024
rect 256325 230966 260084 230968
rect 256325 230963 256391 230966
rect 111793 230346 111859 230349
rect 109910 230344 111859 230346
rect 109910 230288 111798 230344
rect 111854 230288 111859 230344
rect 109910 230286 111859 230288
rect 109910 230112 109970 230286
rect 111793 230283 111859 230286
rect 111885 229938 111951 229941
rect 109910 229936 111951 229938
rect 109910 229880 111890 229936
rect 111946 229880 111951 229936
rect 109910 229878 111951 229880
rect 109910 229432 109970 229878
rect 111885 229875 111951 229878
rect 111793 228986 111859 228989
rect 109910 228984 111859 228986
rect 109910 228928 111798 228984
rect 111854 228928 111859 228984
rect 109910 228926 111859 228928
rect 109910 228752 109970 228926
rect 111793 228923 111859 228926
rect 256693 228986 256759 228989
rect 256693 228984 260084 228986
rect 256693 228928 256698 228984
rect 256754 228928 260084 228984
rect 256693 228926 260084 228928
rect 256693 228923 256759 228926
rect 111885 228578 111951 228581
rect 109910 228576 111951 228578
rect 109910 228520 111890 228576
rect 111946 228520 111951 228576
rect 109910 228518 111951 228520
rect -960 227884 480 228124
rect 109910 228072 109970 228518
rect 111885 228515 111951 228518
rect 111793 227626 111859 227629
rect 109910 227624 111859 227626
rect 109910 227568 111798 227624
rect 111854 227568 111859 227624
rect 109910 227566 111859 227568
rect 109910 227392 109970 227566
rect 111793 227563 111859 227566
rect 111885 227218 111951 227221
rect 109910 227216 111951 227218
rect 109910 227160 111890 227216
rect 111946 227160 111951 227216
rect 109910 227158 111951 227160
rect 109910 226712 109970 227158
rect 111885 227155 111951 227158
rect 256693 226946 256759 226949
rect 256693 226944 260084 226946
rect 256693 226888 256698 226944
rect 256754 226888 260084 226944
rect 256693 226886 260084 226888
rect 256693 226883 256759 226886
rect 112345 226266 112411 226269
rect 109910 226264 112411 226266
rect 109910 226208 112350 226264
rect 112406 226208 112411 226264
rect 109910 226206 112411 226208
rect 109910 226032 109970 226206
rect 112345 226203 112411 226206
rect 111793 225722 111859 225725
rect 109910 225720 111859 225722
rect 109910 225664 111798 225720
rect 111854 225664 111859 225720
rect 109910 225662 111859 225664
rect 109910 225352 109970 225662
rect 111793 225659 111859 225662
rect 256693 224906 256759 224909
rect 256693 224904 260084 224906
rect 256693 224848 256698 224904
rect 256754 224848 260084 224904
rect 256693 224846 260084 224848
rect 256693 224843 256759 224846
rect 111793 224770 111859 224773
rect 109910 224768 111859 224770
rect 109910 224712 111798 224768
rect 111854 224712 111859 224768
rect 109910 224710 111859 224712
rect 109910 224672 109970 224710
rect 111793 224707 111859 224710
rect 111885 224498 111951 224501
rect 109910 224496 111951 224498
rect 109910 224440 111890 224496
rect 111946 224440 111951 224496
rect 109910 224438 111951 224440
rect 109910 223992 109970 224438
rect 111885 224435 111951 224438
rect 111793 223410 111859 223413
rect 109910 223408 111859 223410
rect 109910 223352 111798 223408
rect 111854 223352 111859 223408
rect 109910 223350 111859 223352
rect 109910 223312 109970 223350
rect 111793 223347 111859 223350
rect 111885 223138 111951 223141
rect 109910 223136 111951 223138
rect 109910 223080 111890 223136
rect 111946 223080 111951 223136
rect 109910 223078 111951 223080
rect 109910 222632 109970 223078
rect 111885 223075 111951 223078
rect 256693 222866 256759 222869
rect 256693 222864 260084 222866
rect 256693 222808 256698 222864
rect 256754 222808 260084 222864
rect 256693 222806 260084 222808
rect 256693 222803 256759 222806
rect 111793 222050 111859 222053
rect 109910 222048 111859 222050
rect 109910 221992 111798 222048
rect 111854 221992 111859 222048
rect 109910 221990 111859 221992
rect 109910 221952 109970 221990
rect 111793 221987 111859 221990
rect 111885 221642 111951 221645
rect 109910 221640 111951 221642
rect 109910 221584 111890 221640
rect 111946 221584 111951 221640
rect 109910 221582 111951 221584
rect 109910 221272 109970 221582
rect 111885 221579 111951 221582
rect 256693 220826 256759 220829
rect 256693 220824 260084 220826
rect 256693 220768 256698 220824
rect 256754 220768 260084 220824
rect 256693 220766 260084 220768
rect 256693 220763 256759 220766
rect 111793 220690 111859 220693
rect 109910 220688 111859 220690
rect 109910 220632 111798 220688
rect 111854 220632 111859 220688
rect 109910 220630 111859 220632
rect 109910 220592 109970 220630
rect 111793 220627 111859 220630
rect 111885 220282 111951 220285
rect 109910 220280 111951 220282
rect 109910 220224 111890 220280
rect 111946 220224 111951 220280
rect 109910 220222 111951 220224
rect 109910 219912 109970 220222
rect 111885 220219 111951 220222
rect 112621 219330 112687 219333
rect 109910 219328 112687 219330
rect 109910 219272 112626 219328
rect 112682 219272 112687 219328
rect 109910 219270 112687 219272
rect 109910 219232 109970 219270
rect 112621 219267 112687 219270
rect 112805 219058 112871 219061
rect 109910 219056 112871 219058
rect 109910 219000 112810 219056
rect 112866 219000 112871 219056
rect 109910 218998 112871 219000
rect 109910 218552 109970 218998
rect 112805 218995 112871 218998
rect 580165 219058 580231 219061
rect 583520 219058 584960 219148
rect 580165 219056 584960 219058
rect 580165 219000 580170 219056
rect 580226 219000 584960 219056
rect 580165 218998 584960 219000
rect 580165 218995 580231 218998
rect 583520 218908 584960 218998
rect 256693 218786 256759 218789
rect 256693 218784 260084 218786
rect 256693 218728 256698 218784
rect 256754 218728 260084 218784
rect 256693 218726 260084 218728
rect 256693 218723 256759 218726
rect 111793 217970 111859 217973
rect 109910 217968 111859 217970
rect 109910 217912 111798 217968
rect 111854 217912 111859 217968
rect 109910 217910 111859 217912
rect 109910 217872 109970 217910
rect 111793 217907 111859 217910
rect 111885 217698 111951 217701
rect 109910 217696 111951 217698
rect 109910 217640 111890 217696
rect 111946 217640 111951 217696
rect 109910 217638 111951 217640
rect 109910 217192 109970 217638
rect 111885 217635 111951 217638
rect 256693 216746 256759 216749
rect 256693 216744 260084 216746
rect 256693 216688 256698 216744
rect 256754 216688 260084 216744
rect 256693 216686 260084 216688
rect 256693 216683 256759 216686
rect 112897 216610 112963 216613
rect 109910 216608 112963 216610
rect 109910 216552 112902 216608
rect 112958 216552 112963 216608
rect 109910 216550 112963 216552
rect 109910 216512 109970 216550
rect 112897 216547 112963 216550
rect 111793 216202 111859 216205
rect 109910 216200 111859 216202
rect 109910 216144 111798 216200
rect 111854 216144 111859 216200
rect 109910 216142 111859 216144
rect 109910 215832 109970 216142
rect 111793 216139 111859 216142
rect 111793 215250 111859 215253
rect 109910 215248 111859 215250
rect 109910 215192 111798 215248
rect 111854 215192 111859 215248
rect 109910 215190 111859 215192
rect 109910 215152 109970 215190
rect 111793 215187 111859 215190
rect -960 214978 480 215068
rect 3325 214978 3391 214981
rect -960 214976 3391 214978
rect -960 214920 3330 214976
rect 3386 214920 3391 214976
rect -960 214918 3391 214920
rect -960 214828 480 214918
rect 3325 214915 3391 214918
rect 111885 214842 111951 214845
rect 109910 214840 111951 214842
rect 109910 214784 111890 214840
rect 111946 214784 111951 214840
rect 109910 214782 111951 214784
rect 109910 214472 109970 214782
rect 111885 214779 111951 214782
rect 256693 214706 256759 214709
rect 256693 214704 260084 214706
rect 256693 214648 256698 214704
rect 256754 214648 260084 214704
rect 256693 214646 260084 214648
rect 256693 214643 256759 214646
rect 111793 213890 111859 213893
rect 109910 213888 111859 213890
rect 109910 213832 111798 213888
rect 111854 213832 111859 213888
rect 109910 213830 111859 213832
rect 109910 213792 109970 213830
rect 111793 213827 111859 213830
rect 111885 213482 111951 213485
rect 109910 213480 111951 213482
rect 109910 213424 111890 213480
rect 111946 213424 111951 213480
rect 109910 213422 111951 213424
rect 109910 213112 109970 213422
rect 111885 213419 111951 213422
rect 256693 212666 256759 212669
rect 256693 212664 260084 212666
rect 256693 212608 256698 212664
rect 256754 212608 260084 212664
rect 256693 212606 260084 212608
rect 256693 212603 256759 212606
rect 111793 212530 111859 212533
rect 109910 212528 111859 212530
rect 109910 212472 111798 212528
rect 111854 212472 111859 212528
rect 109910 212470 111859 212472
rect 109910 212432 109970 212470
rect 111793 212467 111859 212470
rect 111885 212122 111951 212125
rect 109910 212120 111951 212122
rect 109910 212064 111890 212120
rect 111946 212064 111951 212120
rect 109910 212062 111951 212064
rect 109910 211752 109970 212062
rect 111885 212059 111951 212062
rect 111793 211170 111859 211173
rect 109910 211168 111859 211170
rect 109910 211112 111798 211168
rect 111854 211112 111859 211168
rect 109910 211110 111859 211112
rect 109910 211072 109970 211110
rect 111793 211107 111859 211110
rect 111885 210762 111951 210765
rect 109910 210760 111951 210762
rect 109910 210704 111890 210760
rect 111946 210704 111951 210760
rect 109910 210702 111951 210704
rect 109910 210392 109970 210702
rect 111885 210699 111951 210702
rect 256693 210626 256759 210629
rect 256693 210624 260084 210626
rect 256693 210568 256698 210624
rect 256754 210568 260084 210624
rect 256693 210566 260084 210568
rect 256693 210563 256759 210566
rect 109910 209674 109970 209712
rect 111793 209674 111859 209677
rect 109910 209672 111859 209674
rect 109910 209616 111798 209672
rect 111854 209616 111859 209672
rect 109910 209614 111859 209616
rect 111793 209611 111859 209614
rect 112437 209402 112503 209405
rect 109910 209400 112503 209402
rect 109910 209344 112442 209400
rect 112498 209344 112503 209400
rect 109910 209342 112503 209344
rect 109910 209032 109970 209342
rect 112437 209339 112503 209342
rect 256233 208586 256299 208589
rect 256233 208584 260084 208586
rect 256233 208528 256238 208584
rect 256294 208528 260084 208584
rect 256233 208526 260084 208528
rect 256233 208523 256299 208526
rect 109910 208314 109970 208352
rect 111793 208314 111859 208317
rect 109910 208312 111859 208314
rect 109910 208256 111798 208312
rect 111854 208256 111859 208312
rect 109910 208254 111859 208256
rect 111793 208251 111859 208254
rect 112345 208178 112411 208181
rect 109910 208176 112411 208178
rect 109910 208120 112350 208176
rect 112406 208120 112411 208176
rect 109910 208118 112411 208120
rect 109910 207672 109970 208118
rect 112345 208115 112411 208118
rect 109910 206954 109970 206992
rect 111793 206954 111859 206957
rect 109910 206952 111859 206954
rect 109910 206896 111798 206952
rect 111854 206896 111859 206952
rect 109910 206894 111859 206896
rect 111793 206891 111859 206894
rect 111885 206682 111951 206685
rect 109910 206680 111951 206682
rect 109910 206624 111890 206680
rect 111946 206624 111951 206680
rect 109910 206622 111951 206624
rect 109910 206312 109970 206622
rect 111885 206619 111951 206622
rect 256693 206546 256759 206549
rect 256693 206544 260084 206546
rect 256693 206488 256698 206544
rect 256754 206488 260084 206544
rect 256693 206486 260084 206488
rect 256693 206483 256759 206486
rect 111977 206138 112043 206141
rect 109910 206136 112043 206138
rect 109910 206080 111982 206136
rect 112038 206080 112043 206136
rect 109910 206078 112043 206080
rect 109910 205632 109970 206078
rect 111977 206075 112043 206078
rect 580441 205730 580507 205733
rect 583520 205730 584960 205820
rect 580441 205728 584960 205730
rect 580441 205672 580446 205728
rect 580502 205672 584960 205728
rect 580441 205670 584960 205672
rect 580441 205667 580507 205670
rect 583520 205580 584960 205670
rect 111793 205050 111859 205053
rect 109910 205048 111859 205050
rect 109910 204992 111798 205048
rect 111854 204992 111859 205048
rect 109910 204990 111859 204992
rect 109910 204952 109970 204990
rect 111793 204987 111859 204990
rect 111885 204778 111951 204781
rect 109910 204776 111951 204778
rect 109910 204720 111890 204776
rect 111946 204720 111951 204776
rect 109910 204718 111951 204720
rect 109910 204272 109970 204718
rect 111885 204715 111951 204718
rect 256693 204506 256759 204509
rect 256693 204504 260084 204506
rect 256693 204448 256698 204504
rect 256754 204448 260084 204504
rect 256693 204446 260084 204448
rect 256693 204443 256759 204446
rect 111793 203690 111859 203693
rect 109910 203688 111859 203690
rect 109910 203632 111798 203688
rect 111854 203632 111859 203688
rect 109910 203630 111859 203632
rect 109910 203592 109970 203630
rect 111793 203627 111859 203630
rect 111885 203418 111951 203421
rect 109910 203416 111951 203418
rect 109910 203360 111890 203416
rect 111946 203360 111951 203416
rect 109910 203358 111951 203360
rect 109910 202912 109970 203358
rect 111885 203355 111951 203358
rect 111793 202602 111859 202605
rect 109910 202600 111859 202602
rect 109910 202544 111798 202600
rect 111854 202544 111859 202600
rect 109910 202542 111859 202544
rect 109910 202232 109970 202542
rect 111793 202539 111859 202542
rect 256693 202466 256759 202469
rect 256693 202464 260084 202466
rect 256693 202408 256698 202464
rect 256754 202408 260084 202464
rect 256693 202406 260084 202408
rect 256693 202403 256759 202406
rect 111885 202058 111951 202061
rect 109910 202056 111951 202058
rect -960 201922 480 202012
rect 109910 202000 111890 202056
rect 111946 202000 111951 202056
rect 109910 201998 111951 202000
rect 3233 201922 3299 201925
rect -960 201920 3299 201922
rect -960 201864 3238 201920
rect 3294 201864 3299 201920
rect -960 201862 3299 201864
rect -960 201772 480 201862
rect 3233 201859 3299 201862
rect 109910 201552 109970 201998
rect 111885 201995 111951 201998
rect 111793 201106 111859 201109
rect 109910 201104 111859 201106
rect 109910 201048 111798 201104
rect 111854 201048 111859 201104
rect 109910 201046 111859 201048
rect 109910 200872 109970 201046
rect 111793 201043 111859 201046
rect 112069 200698 112135 200701
rect 109910 200696 112135 200698
rect 109910 200640 112074 200696
rect 112130 200640 112135 200696
rect 109910 200638 112135 200640
rect 109910 200192 109970 200638
rect 112069 200635 112135 200638
rect 256693 200426 256759 200429
rect 256693 200424 260084 200426
rect 256693 200368 256698 200424
rect 256754 200368 260084 200424
rect 256693 200366 260084 200368
rect 256693 200363 256759 200366
rect 111793 199746 111859 199749
rect 109910 199744 111859 199746
rect 109910 199688 111798 199744
rect 111854 199688 111859 199744
rect 109910 199686 111859 199688
rect 109910 199512 109970 199686
rect 111793 199683 111859 199686
rect 111885 199338 111951 199341
rect 109910 199336 111951 199338
rect 109910 199280 111890 199336
rect 111946 199280 111951 199336
rect 109910 199278 111951 199280
rect 109910 198832 109970 199278
rect 111885 199275 111951 199278
rect 111793 198386 111859 198389
rect 109910 198384 111859 198386
rect 109910 198328 111798 198384
rect 111854 198328 111859 198384
rect 109910 198326 111859 198328
rect 109910 198152 109970 198326
rect 111793 198323 111859 198326
rect 256693 198386 256759 198389
rect 256693 198384 260084 198386
rect 256693 198328 256698 198384
rect 256754 198328 260084 198384
rect 256693 198326 260084 198328
rect 256693 198323 256759 198326
rect 112897 197978 112963 197981
rect 109910 197976 112963 197978
rect 109910 197920 112902 197976
rect 112958 197920 112963 197976
rect 109910 197918 112963 197920
rect 109910 197472 109970 197918
rect 112897 197915 112963 197918
rect 112253 197298 112319 197301
rect 109910 197296 112319 197298
rect 109910 197240 112258 197296
rect 112314 197240 112319 197296
rect 109910 197238 112319 197240
rect 109910 196792 109970 197238
rect 112253 197235 112319 197238
rect 111793 196618 111859 196621
rect 109910 196616 111859 196618
rect 109910 196560 111798 196616
rect 111854 196560 111859 196616
rect 109910 196558 111859 196560
rect 109910 196112 109970 196558
rect 111793 196555 111859 196558
rect 256693 196346 256759 196349
rect 256693 196344 260084 196346
rect 256693 196288 256698 196344
rect 256754 196288 260084 196344
rect 256693 196286 260084 196288
rect 256693 196283 256759 196286
rect 111793 195666 111859 195669
rect 109910 195664 111859 195666
rect 109910 195608 111798 195664
rect 111854 195608 111859 195664
rect 109910 195606 111859 195608
rect 109910 195432 109970 195606
rect 111793 195603 111859 195606
rect 111885 195258 111951 195261
rect 109910 195256 111951 195258
rect 109910 195200 111890 195256
rect 111946 195200 111951 195256
rect 109910 195198 111951 195200
rect 109910 194752 109970 195198
rect 111885 195195 111951 195198
rect 111793 194306 111859 194309
rect 109910 194304 111859 194306
rect 109910 194248 111798 194304
rect 111854 194248 111859 194304
rect 109910 194246 111859 194248
rect 109910 194072 109970 194246
rect 111793 194243 111859 194246
rect 256693 194306 256759 194309
rect 256693 194304 260084 194306
rect 256693 194248 256698 194304
rect 256754 194248 260084 194304
rect 256693 194246 260084 194248
rect 256693 194243 256759 194246
rect 111885 193762 111951 193765
rect 109910 193760 111951 193762
rect 109910 193704 111890 193760
rect 111946 193704 111951 193760
rect 109910 193702 111951 193704
rect 109910 193392 109970 193702
rect 111885 193699 111951 193702
rect 111793 192946 111859 192949
rect 109910 192944 111859 192946
rect 109910 192888 111798 192944
rect 111854 192888 111859 192944
rect 109910 192886 111859 192888
rect 109910 192712 109970 192886
rect 111793 192883 111859 192886
rect 111885 192538 111951 192541
rect 109910 192536 111951 192538
rect 109910 192480 111890 192536
rect 111946 192480 111951 192536
rect 109910 192478 111951 192480
rect 109910 192032 109970 192478
rect 111885 192475 111951 192478
rect 580533 192538 580599 192541
rect 583520 192538 584960 192628
rect 580533 192536 584960 192538
rect 580533 192480 580538 192536
rect 580594 192480 584960 192536
rect 580533 192478 584960 192480
rect 580533 192475 580599 192478
rect 583520 192388 584960 192478
rect 256693 192266 256759 192269
rect 256693 192264 260084 192266
rect 256693 192208 256698 192264
rect 256754 192208 260084 192264
rect 256693 192206 260084 192208
rect 256693 192203 256759 192206
rect 111793 191586 111859 191589
rect 109910 191584 111859 191586
rect 109910 191528 111798 191584
rect 111854 191528 111859 191584
rect 109910 191526 111859 191528
rect 109910 191352 109970 191526
rect 111793 191523 111859 191526
rect 111793 190906 111859 190909
rect 109910 190904 111859 190906
rect 109910 190848 111798 190904
rect 111854 190848 111859 190904
rect 109910 190846 111859 190848
rect 109910 190672 109970 190846
rect 111793 190843 111859 190846
rect 111793 190226 111859 190229
rect 109910 190224 111859 190226
rect 109910 190168 111798 190224
rect 111854 190168 111859 190224
rect 109910 190166 111859 190168
rect 109910 189992 109970 190166
rect 111793 190163 111859 190166
rect 256693 190226 256759 190229
rect 256693 190224 260084 190226
rect 256693 190168 256698 190224
rect 256754 190168 260084 190224
rect 256693 190166 260084 190168
rect 256693 190163 256759 190166
rect 111885 189818 111951 189821
rect 109910 189816 111951 189818
rect 109910 189760 111890 189816
rect 111946 189760 111951 189816
rect 109910 189758 111951 189760
rect 109910 189312 109970 189758
rect 111885 189755 111951 189758
rect -960 188866 480 188956
rect 3601 188866 3667 188869
rect 111793 188866 111859 188869
rect -960 188864 3667 188866
rect -960 188808 3606 188864
rect 3662 188808 3667 188864
rect -960 188806 3667 188808
rect -960 188716 480 188806
rect 3601 188803 3667 188806
rect 109910 188864 111859 188866
rect 109910 188808 111798 188864
rect 111854 188808 111859 188864
rect 109910 188806 111859 188808
rect 109910 188632 109970 188806
rect 111793 188803 111859 188806
rect 111885 188458 111951 188461
rect 109910 188456 111951 188458
rect 109910 188400 111890 188456
rect 111946 188400 111951 188456
rect 109910 188398 111951 188400
rect 109910 187952 109970 188398
rect 111885 188395 111951 188398
rect 256693 188186 256759 188189
rect 256693 188184 260084 188186
rect 256693 188128 256698 188184
rect 256754 188128 260084 188184
rect 256693 188126 260084 188128
rect 256693 188123 256759 188126
rect 111793 187506 111859 187509
rect 109910 187504 111859 187506
rect 109910 187448 111798 187504
rect 111854 187448 111859 187504
rect 109910 187446 111859 187448
rect 109910 187272 109970 187446
rect 111793 187443 111859 187446
rect 111885 187098 111951 187101
rect 109910 187096 111951 187098
rect 109910 187040 111890 187096
rect 111946 187040 111951 187096
rect 109910 187038 111951 187040
rect 109910 186592 109970 187038
rect 111885 187035 111951 187038
rect 112897 186282 112963 186285
rect 109910 186280 112963 186282
rect 109910 186224 112902 186280
rect 112958 186224 112963 186280
rect 109910 186222 112963 186224
rect 109910 185912 109970 186222
rect 112897 186219 112963 186222
rect 256693 186146 256759 186149
rect 256693 186144 260084 186146
rect 256693 186088 256698 186144
rect 256754 186088 260084 186144
rect 256693 186086 260084 186088
rect 256693 186083 256759 186086
rect 111793 185738 111859 185741
rect 109910 185736 111859 185738
rect 109910 185680 111798 185736
rect 111854 185680 111859 185736
rect 109910 185678 111859 185680
rect 109910 185232 109970 185678
rect 111793 185675 111859 185678
rect 111793 184650 111859 184653
rect 109910 184648 111859 184650
rect 109910 184592 111798 184648
rect 111854 184592 111859 184648
rect 109910 184590 111859 184592
rect 109910 184552 109970 184590
rect 111793 184587 111859 184590
rect 111885 184378 111951 184381
rect 109910 184376 111951 184378
rect 109910 184320 111890 184376
rect 111946 184320 111951 184376
rect 109910 184318 111951 184320
rect 109910 183872 109970 184318
rect 111885 184315 111951 184318
rect 256693 184106 256759 184109
rect 256693 184104 260084 184106
rect 256693 184048 256698 184104
rect 256754 184048 260084 184104
rect 256693 184046 260084 184048
rect 256693 184043 256759 184046
rect 112529 183562 112595 183565
rect 109910 183560 112595 183562
rect 109910 183504 112534 183560
rect 112590 183504 112595 183560
rect 109910 183502 112595 183504
rect 109910 183192 109970 183502
rect 112529 183499 112595 183502
rect 111793 183018 111859 183021
rect 109910 183016 111859 183018
rect 109910 182960 111798 183016
rect 111854 182960 111859 183016
rect 109910 182958 111859 182960
rect 109910 182512 109970 182958
rect 111793 182955 111859 182958
rect 111793 182066 111859 182069
rect 109910 182064 111859 182066
rect 109910 182008 111798 182064
rect 111854 182008 111859 182064
rect 109910 182006 111859 182008
rect 109910 181832 109970 182006
rect 111793 182003 111859 182006
rect 256693 182066 256759 182069
rect 256693 182064 260084 182066
rect 256693 182008 256698 182064
rect 256754 182008 260084 182064
rect 256693 182006 260084 182008
rect 256693 182003 256759 182006
rect 111793 181522 111859 181525
rect 109910 181520 111859 181522
rect 109910 181464 111798 181520
rect 111854 181464 111859 181520
rect 109910 181462 111859 181464
rect 109910 181152 109970 181462
rect 111793 181459 111859 181462
rect 111793 180570 111859 180573
rect 109910 180568 111859 180570
rect 109910 180512 111798 180568
rect 111854 180512 111859 180568
rect 109910 180510 111859 180512
rect 109910 180472 109970 180510
rect 111793 180507 111859 180510
rect 111885 180298 111951 180301
rect 109910 180296 111951 180298
rect 109910 180240 111890 180296
rect 111946 180240 111951 180296
rect 109910 180238 111951 180240
rect 109910 179792 109970 180238
rect 111885 180235 111951 180238
rect 256693 180026 256759 180029
rect 256693 180024 260084 180026
rect 256693 179968 256698 180024
rect 256754 179968 260084 180024
rect 256693 179966 260084 179968
rect 256693 179963 256759 179966
rect 111793 179210 111859 179213
rect 109910 179208 111859 179210
rect 109910 179152 111798 179208
rect 111854 179152 111859 179208
rect 109910 179150 111859 179152
rect 109910 179112 109970 179150
rect 111793 179147 111859 179150
rect 580165 179210 580231 179213
rect 583520 179210 584960 179300
rect 580165 179208 584960 179210
rect 580165 179152 580170 179208
rect 580226 179152 584960 179208
rect 580165 179150 584960 179152
rect 580165 179147 580231 179150
rect 583520 179060 584960 179150
rect 111885 178938 111951 178941
rect 109910 178936 111951 178938
rect 109910 178880 111890 178936
rect 111946 178880 111951 178936
rect 109910 178878 111951 178880
rect 109910 178432 109970 178878
rect 111885 178875 111951 178878
rect 112713 177986 112779 177989
rect 109910 177984 112779 177986
rect 109910 177928 112718 177984
rect 112774 177928 112779 177984
rect 109910 177926 112779 177928
rect 109910 177752 109970 177926
rect 112713 177923 112779 177926
rect 256693 177986 256759 177989
rect 256693 177984 260084 177986
rect 256693 177928 256698 177984
rect 256754 177928 260084 177984
rect 256693 177926 260084 177928
rect 256693 177923 256759 177926
rect 112805 177578 112871 177581
rect 109910 177576 112871 177578
rect 109910 177520 112810 177576
rect 112866 177520 112871 177576
rect 109910 177518 112871 177520
rect 109910 177072 109970 177518
rect 112805 177515 112871 177518
rect 111793 176490 111859 176493
rect 109910 176488 111859 176490
rect 109910 176432 111798 176488
rect 111854 176432 111859 176488
rect 109910 176430 111859 176432
rect 109910 176392 109970 176430
rect 111793 176427 111859 176430
rect 111885 176218 111951 176221
rect 109910 176216 111951 176218
rect 109910 176160 111890 176216
rect 111946 176160 111951 176216
rect 109910 176158 111951 176160
rect -960 175796 480 176036
rect 109910 175712 109970 176158
rect 111885 176155 111951 176158
rect 256693 175946 256759 175949
rect 256693 175944 260084 175946
rect 256693 175888 256698 175944
rect 256754 175888 260084 175944
rect 256693 175886 260084 175888
rect 256693 175883 256759 175886
rect 111977 175266 112043 175269
rect 109910 175264 112043 175266
rect 109910 175208 111982 175264
rect 112038 175208 112043 175264
rect 109910 175206 112043 175208
rect 109910 175032 109970 175206
rect 111977 175203 112043 175206
rect 112437 174858 112503 174861
rect 109910 174856 112503 174858
rect 109910 174800 112442 174856
rect 112498 174800 112503 174856
rect 109910 174798 112503 174800
rect 109910 174352 109970 174798
rect 112437 174795 112503 174798
rect 257797 173906 257863 173909
rect 257797 173904 260084 173906
rect 257797 173848 257802 173904
rect 257858 173848 260084 173904
rect 257797 173846 260084 173848
rect 257797 173843 257863 173846
rect 111793 173770 111859 173773
rect 109910 173768 111859 173770
rect 109910 173712 111798 173768
rect 111854 173712 111859 173768
rect 109910 173710 111859 173712
rect 109910 173672 109970 173710
rect 111793 173707 111859 173710
rect 111885 173362 111951 173365
rect 109910 173360 111951 173362
rect 109910 173304 111890 173360
rect 111946 173304 111951 173360
rect 109910 173302 111951 173304
rect 109910 172992 109970 173302
rect 111885 173299 111951 173302
rect 109910 172274 109970 172312
rect 109910 172214 113190 172274
rect 111793 172138 111859 172141
rect 109910 172136 111859 172138
rect 109910 172080 111798 172136
rect 111854 172080 111859 172136
rect 109910 172078 111859 172080
rect 109910 171632 109970 172078
rect 111793 172075 111859 172078
rect 113130 171186 113190 172214
rect 256693 171866 256759 171869
rect 256693 171864 260084 171866
rect 256693 171808 256698 171864
rect 256754 171808 260084 171864
rect 256693 171806 260084 171808
rect 256693 171803 256759 171806
rect 155350 171186 155356 171188
rect 113130 171126 155356 171186
rect 155350 171124 155356 171126
rect 155420 171124 155426 171188
rect 111793 171050 111859 171053
rect 109910 171048 111859 171050
rect 109910 170992 111798 171048
rect 111854 170992 111859 171048
rect 109910 170990 111859 170992
rect 109910 170952 109970 170990
rect 111793 170987 111859 170990
rect 111885 170642 111951 170645
rect 109910 170640 111951 170642
rect 109910 170584 111890 170640
rect 111946 170584 111951 170640
rect 109910 170582 111951 170584
rect 109910 170272 109970 170582
rect 111885 170579 111951 170582
rect 256693 169826 256759 169829
rect 256693 169824 260084 169826
rect 256693 169768 256698 169824
rect 256754 169768 260084 169824
rect 256693 169766 260084 169768
rect 256693 169763 256759 169766
rect 256693 167786 256759 167789
rect 256693 167784 260084 167786
rect 256693 167728 256698 167784
rect 256754 167728 260084 167784
rect 256693 167726 260084 167728
rect 256693 167723 256759 167726
rect 580625 165882 580691 165885
rect 583520 165882 584960 165972
rect 580625 165880 584960 165882
rect 580625 165824 580630 165880
rect 580686 165824 584960 165880
rect 580625 165822 584960 165824
rect 580625 165819 580691 165822
rect 256693 165746 256759 165749
rect 256693 165744 260084 165746
rect 256693 165688 256698 165744
rect 256754 165688 260084 165744
rect 583520 165732 584960 165822
rect 256693 165686 260084 165688
rect 256693 165683 256759 165686
rect 256693 163706 256759 163709
rect 256693 163704 260084 163706
rect 256693 163648 256698 163704
rect 256754 163648 260084 163704
rect 256693 163646 260084 163648
rect 256693 163643 256759 163646
rect -960 162890 480 162980
rect 3325 162890 3391 162893
rect -960 162888 3391 162890
rect -960 162832 3330 162888
rect 3386 162832 3391 162888
rect -960 162830 3391 162832
rect -960 162740 480 162830
rect 3325 162827 3391 162830
rect 256693 161666 256759 161669
rect 256693 161664 260084 161666
rect 256693 161608 256698 161664
rect 256754 161608 260084 161664
rect 256693 161606 260084 161608
rect 256693 161603 256759 161606
rect 256693 159626 256759 159629
rect 256693 159624 260084 159626
rect 256693 159568 256698 159624
rect 256754 159568 260084 159624
rect 256693 159566 260084 159568
rect 256693 159563 256759 159566
rect 257429 157586 257495 157589
rect 257429 157584 260084 157586
rect 257429 157528 257434 157584
rect 257490 157528 260084 157584
rect 257429 157526 260084 157528
rect 257429 157523 257495 157526
rect 256693 155546 256759 155549
rect 256693 155544 260084 155546
rect 256693 155488 256698 155544
rect 256754 155488 260084 155544
rect 256693 155486 260084 155488
rect 256693 155483 256759 155486
rect 256693 153506 256759 153509
rect 256693 153504 260084 153506
rect 256693 153448 256698 153504
rect 256754 153448 260084 153504
rect 256693 153446 260084 153448
rect 256693 153443 256759 153446
rect 579981 152690 580047 152693
rect 583520 152690 584960 152780
rect 579981 152688 584960 152690
rect 579981 152632 579986 152688
rect 580042 152632 584960 152688
rect 579981 152630 584960 152632
rect 579981 152627 580047 152630
rect 583520 152540 584960 152630
rect 256693 151466 256759 151469
rect 256693 151464 260084 151466
rect 256693 151408 256698 151464
rect 256754 151408 260084 151464
rect 256693 151406 260084 151408
rect 256693 151403 256759 151406
rect -960 149834 480 149924
rect 3417 149834 3483 149837
rect -960 149832 3483 149834
rect -960 149776 3422 149832
rect 3478 149776 3483 149832
rect -960 149774 3483 149776
rect -960 149684 480 149774
rect 3417 149771 3483 149774
rect 256693 149426 256759 149429
rect 256693 149424 260084 149426
rect 256693 149368 256698 149424
rect 256754 149368 260084 149424
rect 256693 149366 260084 149368
rect 256693 149363 256759 149366
rect 256693 147386 256759 147389
rect 256693 147384 260084 147386
rect 256693 147328 256698 147384
rect 256754 147328 260084 147384
rect 256693 147326 260084 147328
rect 256693 147323 256759 147326
rect 256693 145346 256759 145349
rect 256693 145344 260084 145346
rect 256693 145288 256698 145344
rect 256754 145288 260084 145344
rect 256693 145286 260084 145288
rect 256693 145283 256759 145286
rect 256693 143306 256759 143309
rect 256693 143304 260084 143306
rect 256693 143248 256698 143304
rect 256754 143248 260084 143304
rect 256693 143246 260084 143248
rect 256693 143243 256759 143246
rect 256693 141266 256759 141269
rect 256693 141264 260084 141266
rect 256693 141208 256698 141264
rect 256754 141208 260084 141264
rect 256693 141206 260084 141208
rect 256693 141203 256759 141206
rect 580165 139362 580231 139365
rect 583520 139362 584960 139452
rect 580165 139360 584960 139362
rect 580165 139304 580170 139360
rect 580226 139304 584960 139360
rect 580165 139302 584960 139304
rect 580165 139299 580231 139302
rect 256693 139226 256759 139229
rect 256693 139224 260084 139226
rect 256693 139168 256698 139224
rect 256754 139168 260084 139224
rect 583520 139212 584960 139302
rect 256693 139166 260084 139168
rect 256693 139163 256759 139166
rect 257521 137186 257587 137189
rect 257521 137184 260084 137186
rect 257521 137128 257526 137184
rect 257582 137128 260084 137184
rect 257521 137126 260084 137128
rect 257521 137123 257587 137126
rect -960 136778 480 136868
rect 3417 136778 3483 136781
rect -960 136776 3483 136778
rect -960 136720 3422 136776
rect 3478 136720 3483 136776
rect -960 136718 3483 136720
rect -960 136628 480 136718
rect 3417 136715 3483 136718
rect 256693 135146 256759 135149
rect 256693 135144 260084 135146
rect 256693 135088 256698 135144
rect 256754 135088 260084 135144
rect 256693 135086 260084 135088
rect 256693 135083 256759 135086
rect 256693 133106 256759 133109
rect 256693 133104 260084 133106
rect 256693 133048 256698 133104
rect 256754 133048 260084 133104
rect 256693 133046 260084 133048
rect 256693 133043 256759 133046
rect 256141 131066 256207 131069
rect 256141 131064 260084 131066
rect 256141 131008 256146 131064
rect 256202 131008 260084 131064
rect 256141 131006 260084 131008
rect 256141 131003 256207 131006
rect 133830 130522 133890 130696
rect 136541 130522 136607 130525
rect 133830 130520 136607 130522
rect 133830 130464 136546 130520
rect 136602 130464 136607 130520
rect 133830 130462 136607 130464
rect 136541 130459 136607 130462
rect 154941 129978 155007 129981
rect 154941 129976 158148 129978
rect 154941 129920 154946 129976
rect 155002 129920 158148 129976
rect 154941 129918 158148 129920
rect 154941 129915 155007 129918
rect 256693 129026 256759 129029
rect 256693 129024 260084 129026
rect 256693 128968 256698 129024
rect 256754 128968 260084 129024
rect 256693 128966 260084 128968
rect 256693 128963 256759 128966
rect 133830 127938 133890 128112
rect 154941 128074 155007 128077
rect 154941 128072 158148 128074
rect 154941 128016 154946 128072
rect 155002 128016 158148 128072
rect 154941 128014 158148 128016
rect 154941 128011 155007 128014
rect 136541 127938 136607 127941
rect 133830 127936 136607 127938
rect 133830 127880 136546 127936
rect 136602 127880 136607 127936
rect 133830 127878 136607 127880
rect 136541 127875 136607 127878
rect 256693 126986 256759 126989
rect 256693 126984 260084 126986
rect 256693 126928 256698 126984
rect 256754 126928 260084 126984
rect 256693 126926 260084 126928
rect 256693 126923 256759 126926
rect 154941 126170 155007 126173
rect 154941 126168 158148 126170
rect 154941 126112 154946 126168
rect 155002 126112 158148 126168
rect 154941 126110 158148 126112
rect 154941 126107 155007 126110
rect 580717 126034 580783 126037
rect 583520 126034 584960 126124
rect 580717 126032 584960 126034
rect 580717 125976 580722 126032
rect 580778 125976 584960 126032
rect 580717 125974 584960 125976
rect 580717 125971 580783 125974
rect 583520 125884 584960 125974
rect 133830 125490 133890 125528
rect 136541 125490 136607 125493
rect 133830 125488 136607 125490
rect 133830 125432 136546 125488
rect 136602 125432 136607 125488
rect 133830 125430 136607 125432
rect 136541 125427 136607 125430
rect 256693 124946 256759 124949
rect 256693 124944 260084 124946
rect 256693 124888 256698 124944
rect 256754 124888 260084 124944
rect 256693 124886 260084 124888
rect 256693 124883 256759 124886
rect 154481 124266 154547 124269
rect 154481 124264 158148 124266
rect 154481 124208 154486 124264
rect 154542 124208 158148 124264
rect 154481 124206 158148 124208
rect 154481 124203 154547 124206
rect -960 123572 480 123812
rect 136173 123586 136239 123589
rect 133830 123584 136239 123586
rect 133830 123528 136178 123584
rect 136234 123528 136239 123584
rect 133830 123526 136239 123528
rect 133830 122944 133890 123526
rect 136173 123523 136239 123526
rect 224166 122844 224172 122908
rect 224236 122906 224242 122908
rect 224236 122846 260084 122906
rect 224236 122844 224242 122846
rect 154941 122362 155007 122365
rect 154941 122360 158148 122362
rect 154941 122304 154946 122360
rect 155002 122304 158148 122360
rect 154941 122302 158148 122304
rect 154941 122299 155007 122302
rect 135253 120866 135319 120869
rect 133830 120864 135319 120866
rect 133830 120808 135258 120864
rect 135314 120808 135319 120864
rect 133830 120806 135319 120808
rect 133830 120360 133890 120806
rect 135253 120803 135319 120806
rect 256693 120866 256759 120869
rect 256693 120864 260084 120866
rect 256693 120808 256698 120864
rect 256754 120808 260084 120864
rect 256693 120806 260084 120808
rect 256693 120803 256759 120806
rect 154573 120458 154639 120461
rect 154573 120456 158148 120458
rect 154573 120400 154578 120456
rect 154634 120400 158148 120456
rect 154573 120398 158148 120400
rect 154573 120395 154639 120398
rect 256693 118826 256759 118829
rect 256693 118824 260084 118826
rect 256693 118768 256698 118824
rect 256754 118768 260084 118824
rect 256693 118766 260084 118768
rect 256693 118763 256759 118766
rect 154573 118554 154639 118557
rect 154573 118552 158148 118554
rect 154573 118496 154578 118552
rect 154634 118496 158148 118552
rect 154573 118494 158148 118496
rect 154573 118491 154639 118494
rect 135437 118282 135503 118285
rect 133830 118280 135503 118282
rect 133830 118224 135442 118280
rect 135498 118224 135503 118280
rect 133830 118222 135503 118224
rect 133830 117776 133890 118222
rect 135437 118219 135503 118222
rect 256693 116786 256759 116789
rect 256693 116784 260084 116786
rect 256693 116728 256698 116784
rect 256754 116728 260084 116784
rect 256693 116726 260084 116728
rect 256693 116723 256759 116726
rect 155401 116650 155467 116653
rect 155401 116648 158148 116650
rect 155401 116592 155406 116648
rect 155462 116592 158148 116648
rect 155401 116590 158148 116592
rect 155401 116587 155467 116590
rect 136541 115562 136607 115565
rect 133830 115560 136607 115562
rect 133830 115504 136546 115560
rect 136602 115504 136607 115560
rect 133830 115502 136607 115504
rect 133830 115192 133890 115502
rect 136541 115499 136607 115502
rect 154757 114746 154823 114749
rect 256693 114746 256759 114749
rect 154757 114744 158148 114746
rect 154757 114688 154762 114744
rect 154818 114688 158148 114744
rect 154757 114686 158148 114688
rect 256693 114744 260084 114746
rect 256693 114688 256698 114744
rect 256754 114688 260084 114744
rect 256693 114686 260084 114688
rect 154757 114683 154823 114686
rect 256693 114683 256759 114686
rect 136541 112842 136607 112845
rect 133830 112840 136607 112842
rect 133830 112784 136546 112840
rect 136602 112784 136607 112840
rect 133830 112782 136607 112784
rect 133830 112608 133890 112782
rect 136541 112779 136607 112782
rect 154941 112842 155007 112845
rect 580165 112842 580231 112845
rect 583520 112842 584960 112932
rect 154941 112840 158148 112842
rect 154941 112784 154946 112840
rect 155002 112784 158148 112840
rect 154941 112782 158148 112784
rect 580165 112840 584960 112842
rect 580165 112784 580170 112840
rect 580226 112784 584960 112840
rect 580165 112782 584960 112784
rect 154941 112779 155007 112782
rect 580165 112779 580231 112782
rect 256693 112706 256759 112709
rect 256693 112704 260084 112706
rect 256693 112648 256698 112704
rect 256754 112648 260084 112704
rect 583520 112692 584960 112782
rect 256693 112646 260084 112648
rect 256693 112643 256759 112646
rect 154849 110938 154915 110941
rect 154849 110936 158148 110938
rect 154849 110880 154854 110936
rect 154910 110880 158148 110936
rect 154849 110878 158148 110880
rect 154849 110875 154915 110878
rect -960 110666 480 110756
rect 3417 110666 3483 110669
rect -960 110664 3483 110666
rect -960 110608 3422 110664
rect 3478 110608 3483 110664
rect -960 110606 3483 110608
rect -960 110516 480 110606
rect 3417 110603 3483 110606
rect 256693 110666 256759 110669
rect 256693 110664 260084 110666
rect 256693 110608 256698 110664
rect 256754 110608 260084 110664
rect 256693 110606 260084 110608
rect 256693 110603 256759 110606
rect 136541 110258 136607 110261
rect 133830 110256 136607 110258
rect 133830 110200 136546 110256
rect 136602 110200 136607 110256
rect 133830 110198 136607 110200
rect 133830 110024 133890 110198
rect 136541 110195 136607 110198
rect 155493 109034 155559 109037
rect 155493 109032 158148 109034
rect 155493 108976 155498 109032
rect 155554 108976 158148 109032
rect 155493 108974 158148 108976
rect 155493 108971 155559 108974
rect 256693 108626 256759 108629
rect 256693 108624 260084 108626
rect 256693 108568 256698 108624
rect 256754 108568 260084 108624
rect 256693 108566 260084 108568
rect 256693 108563 256759 108566
rect 136541 107538 136607 107541
rect 133830 107536 136607 107538
rect 133830 107480 136546 107536
rect 136602 107480 136607 107536
rect 133830 107478 136607 107480
rect 133830 107440 133890 107478
rect 136541 107475 136607 107478
rect 155309 107130 155375 107133
rect 155309 107128 158148 107130
rect 155309 107072 155314 107128
rect 155370 107072 158148 107128
rect 155309 107070 158148 107072
rect 155309 107067 155375 107070
rect 256693 106586 256759 106589
rect 256693 106584 260084 106586
rect 256693 106528 256698 106584
rect 256754 106528 260084 106584
rect 256693 106526 260084 106528
rect 256693 106523 256759 106526
rect 154573 105226 154639 105229
rect 154573 105224 158148 105226
rect 154573 105168 154578 105224
rect 154634 105168 158148 105224
rect 154573 105166 158148 105168
rect 154573 105163 154639 105166
rect 133830 104818 133890 104856
rect 136541 104818 136607 104821
rect 133830 104816 136607 104818
rect 133830 104760 136546 104816
rect 136602 104760 136607 104816
rect 133830 104758 136607 104760
rect 136541 104755 136607 104758
rect 256693 104546 256759 104549
rect 256693 104544 260084 104546
rect 256693 104488 256698 104544
rect 256754 104488 260084 104544
rect 256693 104486 260084 104488
rect 256693 104483 256759 104486
rect 154573 103322 154639 103325
rect 154573 103320 158148 103322
rect 154573 103264 154578 103320
rect 154634 103264 158148 103320
rect 154573 103262 158148 103264
rect 154573 103259 154639 103262
rect 136173 102914 136239 102917
rect 133830 102912 136239 102914
rect 133830 102856 136178 102912
rect 136234 102856 136239 102912
rect 133830 102854 136239 102856
rect 133830 102272 133890 102854
rect 136173 102851 136239 102854
rect 256693 102506 256759 102509
rect 256693 102504 260084 102506
rect 256693 102448 256698 102504
rect 256754 102448 260084 102504
rect 256693 102446 260084 102448
rect 256693 102443 256759 102446
rect 154941 101418 155007 101421
rect 154941 101416 158148 101418
rect 154941 101360 154946 101416
rect 155002 101360 158148 101416
rect 154941 101358 158148 101360
rect 154941 101355 155007 101358
rect 256693 100466 256759 100469
rect 256693 100464 260084 100466
rect 256693 100408 256698 100464
rect 256754 100408 260084 100464
rect 256693 100406 260084 100408
rect 256693 100403 256759 100406
rect 136173 100194 136239 100197
rect 133830 100192 136239 100194
rect 133830 100136 136178 100192
rect 136234 100136 136239 100192
rect 133830 100134 136239 100136
rect 133830 99688 133890 100134
rect 136173 100131 136239 100134
rect 154941 99514 155007 99517
rect 580809 99514 580875 99517
rect 583520 99514 584960 99604
rect 154941 99512 158148 99514
rect 154941 99456 154946 99512
rect 155002 99456 158148 99512
rect 154941 99454 158148 99456
rect 580809 99512 584960 99514
rect 580809 99456 580814 99512
rect 580870 99456 584960 99512
rect 580809 99454 584960 99456
rect 154941 99451 155007 99454
rect 580809 99451 580875 99454
rect 583520 99364 584960 99454
rect 256049 98426 256115 98429
rect 256049 98424 260084 98426
rect 256049 98368 256054 98424
rect 256110 98368 260084 98424
rect 256049 98366 260084 98368
rect 256049 98363 256115 98366
rect 136725 97746 136791 97749
rect 133830 97744 136791 97746
rect -960 97610 480 97700
rect 133830 97688 136730 97744
rect 136786 97688 136791 97744
rect 133830 97686 136791 97688
rect 3417 97610 3483 97613
rect -960 97608 3483 97610
rect -960 97552 3422 97608
rect 3478 97552 3483 97608
rect -960 97550 3483 97552
rect -960 97460 480 97550
rect 3417 97547 3483 97550
rect 133830 97104 133890 97686
rect 136725 97683 136791 97686
rect 154849 97610 154915 97613
rect 154849 97608 158148 97610
rect 154849 97552 154854 97608
rect 154910 97552 158148 97608
rect 154849 97550 158148 97552
rect 154849 97547 154915 97550
rect 256693 96386 256759 96389
rect 256693 96384 260084 96386
rect 256693 96328 256698 96384
rect 256754 96328 260084 96384
rect 256693 96326 260084 96328
rect 256693 96323 256759 96326
rect 154941 95706 155007 95709
rect 154941 95704 158148 95706
rect 154941 95648 154946 95704
rect 155002 95648 158148 95704
rect 154941 95646 158148 95648
rect 154941 95643 155007 95646
rect 136541 95162 136607 95165
rect 133830 95160 136607 95162
rect 133830 95104 136546 95160
rect 136602 95104 136607 95160
rect 133830 95102 136607 95104
rect 133830 94520 133890 95102
rect 136541 95099 136607 95102
rect 256693 94346 256759 94349
rect 256693 94344 260084 94346
rect 256693 94288 256698 94344
rect 256754 94288 260084 94344
rect 256693 94286 260084 94288
rect 256693 94283 256759 94286
rect 154573 93802 154639 93805
rect 154573 93800 158148 93802
rect 154573 93744 154578 93800
rect 154634 93744 158148 93800
rect 154573 93742 158148 93744
rect 154573 93739 154639 93742
rect 136081 92442 136147 92445
rect 133830 92440 136147 92442
rect 133830 92384 136086 92440
rect 136142 92384 136147 92440
rect 133830 92382 136147 92384
rect 133830 91936 133890 92382
rect 136081 92379 136147 92382
rect 256693 92306 256759 92309
rect 256693 92304 260084 92306
rect 256693 92248 256698 92304
rect 256754 92248 260084 92304
rect 256693 92246 260084 92248
rect 256693 92243 256759 92246
rect 154941 91898 155007 91901
rect 154941 91896 158148 91898
rect 154941 91840 154946 91896
rect 155002 91840 158148 91896
rect 154941 91838 158148 91840
rect 154941 91835 155007 91838
rect 256693 90266 256759 90269
rect 256693 90264 260084 90266
rect 256693 90208 256698 90264
rect 256754 90208 260084 90264
rect 256693 90206 260084 90208
rect 256693 90203 256759 90206
rect 154941 89994 155007 89997
rect 154941 89992 158148 89994
rect 154941 89936 154946 89992
rect 155002 89936 158148 89992
rect 154941 89934 158148 89936
rect 154941 89931 155007 89934
rect 136541 89586 136607 89589
rect 133830 89584 136607 89586
rect 133830 89528 136546 89584
rect 136602 89528 136607 89584
rect 133830 89526 136607 89528
rect 133830 89352 133890 89526
rect 136541 89523 136607 89526
rect 256693 88226 256759 88229
rect 256693 88224 260084 88226
rect 256693 88168 256698 88224
rect 256754 88168 260084 88224
rect 256693 88166 260084 88168
rect 256693 88163 256759 88166
rect 154941 88090 155007 88093
rect 154941 88088 158148 88090
rect 154941 88032 154946 88088
rect 155002 88032 158148 88088
rect 154941 88030 158148 88032
rect 154941 88027 155007 88030
rect 135253 86866 135319 86869
rect 133830 86864 135319 86866
rect 133830 86808 135258 86864
rect 135314 86808 135319 86864
rect 133830 86806 135319 86808
rect 133830 86768 133890 86806
rect 135253 86803 135319 86806
rect 154941 86186 155007 86189
rect 256693 86186 256759 86189
rect 580901 86186 580967 86189
rect 583520 86186 584960 86276
rect 154941 86184 158148 86186
rect 154941 86128 154946 86184
rect 155002 86128 158148 86184
rect 154941 86126 158148 86128
rect 256693 86184 260084 86186
rect 256693 86128 256698 86184
rect 256754 86128 260084 86184
rect 256693 86126 260084 86128
rect 580901 86184 584960 86186
rect 580901 86128 580906 86184
rect 580962 86128 584960 86184
rect 580901 86126 584960 86128
rect 154941 86123 155007 86126
rect 256693 86123 256759 86126
rect 580901 86123 580967 86126
rect 583520 86036 584960 86126
rect 135805 84826 135871 84829
rect 133830 84824 135871 84826
rect -960 84690 480 84780
rect 133830 84768 135810 84824
rect 135866 84768 135871 84824
rect 133830 84766 135871 84768
rect 3417 84690 3483 84693
rect -960 84688 3483 84690
rect -960 84632 3422 84688
rect 3478 84632 3483 84688
rect -960 84630 3483 84632
rect -960 84540 480 84630
rect 3417 84627 3483 84630
rect 133830 84184 133890 84766
rect 135805 84763 135871 84766
rect 154941 84282 155007 84285
rect 154941 84280 158148 84282
rect 154941 84224 154946 84280
rect 155002 84224 158148 84280
rect 154941 84222 158148 84224
rect 154941 84219 155007 84222
rect 256693 84146 256759 84149
rect 256693 84144 260084 84146
rect 256693 84088 256698 84144
rect 256754 84088 260084 84144
rect 256693 84086 260084 84088
rect 256693 84083 256759 84086
rect 154941 82378 155007 82381
rect 154941 82376 158148 82378
rect 154941 82320 154946 82376
rect 155002 82320 158148 82376
rect 154941 82318 158148 82320
rect 154941 82315 155007 82318
rect 136541 82242 136607 82245
rect 133830 82240 136607 82242
rect 133830 82184 136546 82240
rect 136602 82184 136607 82240
rect 133830 82182 136607 82184
rect 133830 81600 133890 82182
rect 136541 82179 136607 82182
rect 256693 82106 256759 82109
rect 256693 82104 260084 82106
rect 256693 82048 256698 82104
rect 256754 82048 260084 82104
rect 256693 82046 260084 82048
rect 256693 82043 256759 82046
rect 154757 80474 154823 80477
rect 154757 80472 158148 80474
rect 154757 80416 154762 80472
rect 154818 80416 158148 80472
rect 154757 80414 158148 80416
rect 154757 80411 154823 80414
rect 256693 80066 256759 80069
rect 256693 80064 260084 80066
rect 256693 80008 256698 80064
rect 256754 80008 260084 80064
rect 256693 80006 260084 80008
rect 256693 80003 256759 80006
rect 136081 79658 136147 79661
rect 133830 79656 136147 79658
rect 133830 79600 136086 79656
rect 136142 79600 136147 79656
rect 133830 79598 136147 79600
rect 133830 79016 133890 79598
rect 136081 79595 136147 79598
rect 154941 78570 155007 78573
rect 154941 78568 158148 78570
rect 154941 78512 154946 78568
rect 155002 78512 158148 78568
rect 154941 78510 158148 78512
rect 154941 78507 155007 78510
rect 256693 78026 256759 78029
rect 256693 78024 260084 78026
rect 256693 77968 256698 78024
rect 256754 77968 260084 78024
rect 256693 77966 260084 77968
rect 256693 77963 256759 77966
rect 136541 77074 136607 77077
rect 133830 77072 136607 77074
rect 133830 77016 136546 77072
rect 136602 77016 136607 77072
rect 133830 77014 136607 77016
rect 133830 76432 133890 77014
rect 136541 77011 136607 77014
rect 154941 76666 155007 76669
rect 154941 76664 158148 76666
rect 154941 76608 154946 76664
rect 155002 76608 158148 76664
rect 154941 76606 158148 76608
rect 154941 76603 155007 76606
rect 256693 75986 256759 75989
rect 256693 75984 260084 75986
rect 256693 75928 256698 75984
rect 256754 75928 260084 75984
rect 256693 75926 260084 75928
rect 256693 75923 256759 75926
rect 154941 74762 155007 74765
rect 154941 74760 158148 74762
rect 154941 74704 154946 74760
rect 155002 74704 158148 74760
rect 154941 74702 158148 74704
rect 154941 74699 155007 74702
rect 256693 73946 256759 73949
rect 256693 73944 260084 73946
rect 256693 73888 256698 73944
rect 256754 73888 260084 73944
rect 256693 73886 260084 73888
rect 256693 73883 256759 73886
rect 133830 73810 133890 73848
rect 136541 73810 136607 73813
rect 133830 73808 136607 73810
rect 133830 73752 136546 73808
rect 136602 73752 136607 73808
rect 133830 73750 136607 73752
rect 136541 73747 136607 73750
rect 580165 72994 580231 72997
rect 583520 72994 584960 73084
rect 580165 72992 584960 72994
rect 580165 72936 580170 72992
rect 580226 72936 584960 72992
rect 580165 72934 584960 72936
rect 580165 72931 580231 72934
rect 154573 72858 154639 72861
rect 154573 72856 158148 72858
rect 154573 72800 154578 72856
rect 154634 72800 158148 72856
rect 583520 72844 584960 72934
rect 154573 72798 158148 72800
rect 154573 72795 154639 72798
rect 256693 71906 256759 71909
rect 256693 71904 260084 71906
rect 256693 71848 256698 71904
rect 256754 71848 260084 71904
rect 256693 71846 260084 71848
rect 256693 71843 256759 71846
rect -960 71634 480 71724
rect 3509 71634 3575 71637
rect 135345 71634 135411 71637
rect -960 71632 3575 71634
rect -960 71576 3514 71632
rect 3570 71576 3575 71632
rect -960 71574 3575 71576
rect -960 71484 480 71574
rect 3509 71571 3575 71574
rect 133830 71632 135411 71634
rect 133830 71576 135350 71632
rect 135406 71576 135411 71632
rect 133830 71574 135411 71576
rect 133830 71264 133890 71574
rect 135345 71571 135411 71574
rect 154941 70954 155007 70957
rect 154941 70952 158148 70954
rect 154941 70896 154946 70952
rect 155002 70896 158148 70952
rect 154941 70894 158148 70896
rect 154941 70891 155007 70894
rect 256693 69866 256759 69869
rect 256693 69864 260084 69866
rect 256693 69808 256698 69864
rect 256754 69808 260084 69864
rect 256693 69806 260084 69808
rect 256693 69803 256759 69806
rect 154573 69050 154639 69053
rect 154573 69048 158148 69050
rect 154573 68992 154578 69048
rect 154634 68992 158148 69048
rect 154573 68990 158148 68992
rect 154573 68987 154639 68990
rect 135713 68914 135779 68917
rect 133830 68912 135779 68914
rect 133830 68856 135718 68912
rect 135774 68856 135779 68912
rect 133830 68854 135779 68856
rect 133830 68680 133890 68854
rect 135713 68851 135779 68854
rect 256693 67826 256759 67829
rect 256693 67824 260084 67826
rect 256693 67768 256698 67824
rect 256754 67768 260084 67824
rect 256693 67766 260084 67768
rect 256693 67763 256759 67766
rect 154941 67146 155007 67149
rect 154941 67144 158148 67146
rect 154941 67088 154946 67144
rect 155002 67088 158148 67144
rect 154941 67086 158148 67088
rect 154941 67083 155007 67086
rect 136081 66194 136147 66197
rect 133830 66192 136147 66194
rect 133830 66136 136086 66192
rect 136142 66136 136147 66192
rect 133830 66134 136147 66136
rect 133830 66096 133890 66134
rect 136081 66131 136147 66134
rect 257429 65786 257495 65789
rect 257429 65784 260084 65786
rect 257429 65728 257434 65784
rect 257490 65728 260084 65784
rect 257429 65726 260084 65728
rect 257429 65723 257495 65726
rect 154573 65242 154639 65245
rect 154573 65240 158148 65242
rect 154573 65184 154578 65240
rect 154634 65184 158148 65240
rect 154573 65182 158148 65184
rect 154573 65179 154639 65182
rect 136541 64154 136607 64157
rect 133830 64152 136607 64154
rect 133830 64096 136546 64152
rect 136602 64096 136607 64152
rect 133830 64094 136607 64096
rect 133830 63512 133890 64094
rect 136541 64091 136607 64094
rect 256693 63746 256759 63749
rect 256693 63744 260084 63746
rect 256693 63688 256698 63744
rect 256754 63688 260084 63744
rect 256693 63686 260084 63688
rect 256693 63683 256759 63686
rect 154573 63338 154639 63341
rect 154573 63336 158148 63338
rect 154573 63280 154578 63336
rect 154634 63280 158148 63336
rect 154573 63278 158148 63280
rect 154573 63275 154639 63278
rect 256693 61706 256759 61709
rect 256693 61704 260084 61706
rect 256693 61648 256698 61704
rect 256754 61648 260084 61704
rect 256693 61646 260084 61648
rect 256693 61643 256759 61646
rect 135621 61570 135687 61573
rect 133830 61568 135687 61570
rect 133830 61512 135626 61568
rect 135682 61512 135687 61568
rect 133830 61510 135687 61512
rect 133830 60928 133890 61510
rect 135621 61507 135687 61510
rect 154941 61434 155007 61437
rect 154941 61432 158148 61434
rect 154941 61376 154946 61432
rect 155002 61376 158148 61432
rect 154941 61374 158148 61376
rect 154941 61371 155007 61374
rect 256693 59666 256759 59669
rect 580073 59666 580139 59669
rect 583520 59666 584960 59756
rect 256693 59664 260084 59666
rect 256693 59608 256698 59664
rect 256754 59608 260084 59664
rect 256693 59606 260084 59608
rect 580073 59664 584960 59666
rect 580073 59608 580078 59664
rect 580134 59608 584960 59664
rect 580073 59606 584960 59608
rect 256693 59603 256759 59606
rect 580073 59603 580139 59606
rect 154941 59530 155007 59533
rect 154941 59528 158148 59530
rect 154941 59472 154946 59528
rect 155002 59472 158148 59528
rect 583520 59516 584960 59606
rect 154941 59470 158148 59472
rect 154941 59467 155007 59470
rect 136541 58986 136607 58989
rect 133830 58984 136607 58986
rect 133830 58928 136546 58984
rect 136602 58928 136607 58984
rect 133830 58926 136607 58928
rect -960 58578 480 58668
rect 3601 58578 3667 58581
rect -960 58576 3667 58578
rect -960 58520 3606 58576
rect 3662 58520 3667 58576
rect -960 58518 3667 58520
rect -960 58428 480 58518
rect 3601 58515 3667 58518
rect 133830 58344 133890 58926
rect 136541 58923 136607 58926
rect 154941 57626 155007 57629
rect 256693 57626 256759 57629
rect 154941 57624 158148 57626
rect 154941 57568 154946 57624
rect 155002 57568 158148 57624
rect 154941 57566 158148 57568
rect 256693 57624 260084 57626
rect 256693 57568 256698 57624
rect 256754 57568 260084 57624
rect 256693 57566 260084 57568
rect 154941 57563 155007 57566
rect 256693 57563 256759 57566
rect 135253 56402 135319 56405
rect 133830 56400 135319 56402
rect 133830 56344 135258 56400
rect 135314 56344 135319 56400
rect 133830 56342 135319 56344
rect 133830 55760 133890 56342
rect 135253 56339 135319 56342
rect 154941 55722 155007 55725
rect 154941 55720 158148 55722
rect 154941 55664 154946 55720
rect 155002 55664 158148 55720
rect 154941 55662 158148 55664
rect 154941 55659 155007 55662
rect 256693 55586 256759 55589
rect 256693 55584 260084 55586
rect 256693 55528 256698 55584
rect 256754 55528 260084 55584
rect 256693 55526 260084 55528
rect 256693 55523 256759 55526
rect 154941 53818 155007 53821
rect 154941 53816 158148 53818
rect 154941 53760 154946 53816
rect 155002 53760 158148 53816
rect 154941 53758 158148 53760
rect 154941 53755 155007 53758
rect 136541 53546 136607 53549
rect 133830 53544 136607 53546
rect 133830 53488 136546 53544
rect 136602 53488 136607 53544
rect 133830 53486 136607 53488
rect 133830 53176 133890 53486
rect 136541 53483 136607 53486
rect 257337 53546 257403 53549
rect 257337 53544 260084 53546
rect 257337 53488 257342 53544
rect 257398 53488 260084 53544
rect 257337 53486 260084 53488
rect 257337 53483 257403 53486
rect 208710 52804 208716 52868
rect 208780 52866 208786 52868
rect 216673 52866 216739 52869
rect 208780 52864 216739 52866
rect 208780 52808 216678 52864
rect 216734 52808 216739 52864
rect 208780 52806 216739 52808
rect 208780 52804 208786 52806
rect 216673 52803 216739 52806
rect 173566 52668 173572 52732
rect 173636 52730 173642 52732
rect 251766 52730 251772 52732
rect 173636 52670 251772 52730
rect 173636 52668 173642 52670
rect 251766 52668 251772 52670
rect 251836 52668 251842 52732
rect 169886 52260 169892 52324
rect 169956 52322 169962 52324
rect 194358 52322 194364 52324
rect 169956 52262 178234 52322
rect 169956 52260 169962 52262
rect 157977 52186 158043 52189
rect 157977 52184 176210 52186
rect 157977 52128 157982 52184
rect 158038 52128 176210 52184
rect 157977 52126 176210 52128
rect 157977 52123 158043 52126
rect 161790 51988 161796 52052
rect 161860 52050 161866 52052
rect 161860 51988 161904 52050
rect 163630 51988 163636 52052
rect 163700 52050 163706 52052
rect 169150 52050 169156 52052
rect 163700 51990 163836 52050
rect 163700 51988 163706 51990
rect 161335 51948 161401 51951
rect 161335 51946 161444 51948
rect 160323 51916 160389 51917
rect 160318 51914 160324 51916
rect 160232 51854 160324 51914
rect 160318 51852 160324 51854
rect 160388 51852 160394 51916
rect 160967 51914 161033 51917
rect 160967 51912 161076 51914
rect 160507 51878 160573 51883
rect 160323 51851 160389 51852
rect 160507 51822 160512 51878
rect 160568 51822 160573 51878
rect 160967 51856 160972 51912
rect 161028 51856 161076 51912
rect 161335 51890 161340 51946
rect 161396 51916 161444 51946
rect 161396 51890 161428 51916
rect 161335 51885 161428 51890
rect 160967 51851 161076 51856
rect 161384 51854 161428 51885
rect 161422 51852 161428 51854
rect 161492 51852 161498 51916
rect 161703 51914 161769 51917
rect 161844 51914 161904 51988
rect 161703 51912 161904 51914
rect 161703 51856 161708 51912
rect 161764 51856 161904 51912
rect 161703 51854 161904 51856
rect 161979 51914 162045 51917
rect 162158 51914 162164 51916
rect 161979 51912 162164 51914
rect 161979 51856 161984 51912
rect 162040 51856 162164 51912
rect 161979 51854 162164 51856
rect 161703 51851 161769 51854
rect 161979 51851 162045 51854
rect 162158 51852 162164 51854
rect 162228 51852 162234 51916
rect 162439 51914 162505 51917
rect 162715 51916 162781 51917
rect 162710 51914 162716 51916
rect 162304 51912 162505 51914
rect 162304 51856 162444 51912
rect 162500 51856 162505 51912
rect 162304 51854 162505 51856
rect 162624 51854 162716 51914
rect 160507 51817 160573 51822
rect 160185 51780 160251 51781
rect 160134 51778 160140 51780
rect 160094 51718 160140 51778
rect 160204 51776 160251 51780
rect 160246 51720 160251 51776
rect 160134 51716 160140 51718
rect 160204 51716 160251 51720
rect 160185 51715 160251 51716
rect 159909 51642 159975 51645
rect 160510 51642 160570 51817
rect 159909 51640 160570 51642
rect 159909 51584 159914 51640
rect 159970 51584 160570 51640
rect 159909 51582 160570 51584
rect 160645 51642 160711 51645
rect 161016 51642 161076 51851
rect 161151 51778 161217 51781
rect 161381 51778 161447 51781
rect 161151 51776 161447 51778
rect 161151 51720 161156 51776
rect 161212 51720 161386 51776
rect 161442 51720 161447 51776
rect 161151 51718 161447 51720
rect 161151 51715 161217 51718
rect 161381 51715 161447 51718
rect 160645 51640 161076 51642
rect 160645 51584 160650 51640
rect 160706 51584 161076 51640
rect 160645 51582 161076 51584
rect 159909 51579 159975 51582
rect 160645 51579 160711 51582
rect 161606 51580 161612 51644
rect 161676 51642 161682 51644
rect 161749 51642 161815 51645
rect 161676 51640 161815 51642
rect 161676 51584 161754 51640
rect 161810 51584 161815 51640
rect 161676 51582 161815 51584
rect 161676 51580 161682 51582
rect 161749 51579 161815 51582
rect 162304 51509 162364 51854
rect 162439 51851 162505 51854
rect 162710 51852 162716 51854
rect 162780 51852 162786 51916
rect 163451 51912 163517 51917
rect 163451 51856 163456 51912
rect 163512 51856 163517 51912
rect 162715 51851 162781 51852
rect 163451 51851 163517 51856
rect 163776 51914 163836 51990
rect 168790 51990 169156 52050
rect 165383 51948 165449 51951
rect 165383 51946 165492 51948
rect 163911 51914 163977 51917
rect 163776 51912 163977 51914
rect 163776 51856 163916 51912
rect 163972 51856 163977 51912
rect 163776 51854 163977 51856
rect 163911 51851 163977 51854
rect 164095 51914 164161 51917
rect 164095 51912 164296 51914
rect 164095 51856 164100 51912
rect 164156 51856 164296 51912
rect 164095 51854 164296 51856
rect 164095 51851 164161 51854
rect 162991 51812 163057 51815
rect 162948 51810 163057 51812
rect 162948 51780 162996 51810
rect 162894 51716 162900 51780
rect 162964 51754 162996 51780
rect 163052 51754 163057 51810
rect 162964 51749 163057 51754
rect 162964 51718 163008 51749
rect 162964 51716 162970 51718
rect 163454 51645 163514 51851
rect 163635 51810 163701 51815
rect 163635 51754 163640 51810
rect 163696 51754 163701 51810
rect 163635 51749 163701 51754
rect 164049 51778 164115 51781
rect 164236 51778 164296 51854
rect 164463 51912 164529 51917
rect 164463 51856 164468 51912
rect 164524 51856 164529 51912
rect 164463 51851 164529 51856
rect 164739 51912 164805 51917
rect 164739 51856 164744 51912
rect 164800 51856 164805 51912
rect 165383 51890 165388 51946
rect 165444 51890 165492 51946
rect 165383 51885 165492 51890
rect 165567 51946 165633 51951
rect 165567 51890 165572 51946
rect 165628 51890 165633 51946
rect 165843 51946 165909 51951
rect 166671 51948 166737 51951
rect 167591 51948 167657 51951
rect 167775 51948 167841 51951
rect 165843 51916 165848 51946
rect 165904 51916 165909 51946
rect 166398 51946 166737 51948
rect 165567 51885 165633 51890
rect 164739 51851 164805 51856
rect 164049 51776 164296 51778
rect 163454 51640 163563 51645
rect 163454 51584 163502 51640
rect 163558 51584 163563 51640
rect 163454 51582 163563 51584
rect 163497 51579 163563 51582
rect 162301 51504 162367 51509
rect 162301 51448 162306 51504
rect 162362 51448 162367 51504
rect 162301 51443 162367 51448
rect 162761 51506 162827 51509
rect 163638 51506 163698 51749
rect 164049 51720 164054 51776
rect 164110 51720 164296 51776
rect 164049 51718 164296 51720
rect 164049 51715 164115 51718
rect 162761 51504 163698 51506
rect 162761 51448 162766 51504
rect 162822 51448 163698 51504
rect 162761 51446 163698 51448
rect 162761 51443 162827 51446
rect 163814 51444 163820 51508
rect 163884 51506 163890 51508
rect 164466 51506 164526 51851
rect 163884 51446 164526 51506
rect 163884 51444 163890 51446
rect 164742 51373 164802 51851
rect 164877 51778 164943 51781
rect 165291 51778 165357 51781
rect 164877 51776 165357 51778
rect 164877 51720 164882 51776
rect 164938 51720 165296 51776
rect 165352 51720 165357 51776
rect 164877 51718 165357 51720
rect 164877 51715 164943 51718
rect 165291 51715 165357 51718
rect 165432 51645 165492 51885
rect 165061 51642 165127 51645
rect 165061 51640 165170 51642
rect 165061 51584 165066 51640
rect 165122 51584 165170 51640
rect 165061 51579 165170 51584
rect 165429 51640 165495 51645
rect 165429 51584 165434 51640
rect 165490 51584 165495 51640
rect 165429 51579 165495 51584
rect 164693 51368 164802 51373
rect 164693 51312 164698 51368
rect 164754 51312 164802 51368
rect 164693 51310 164802 51312
rect 165110 51373 165170 51579
rect 165245 51506 165311 51509
rect 165570 51506 165630 51885
rect 165838 51852 165844 51916
rect 165908 51914 165914 51916
rect 166119 51914 166185 51917
rect 165908 51854 165966 51914
rect 166076 51912 166185 51914
rect 166076 51856 166124 51912
rect 166180 51856 166185 51912
rect 165908 51852 165914 51854
rect 166076 51851 166185 51856
rect 166398 51890 166676 51946
rect 166732 51890 166737 51946
rect 167548 51946 167657 51948
rect 167548 51916 167596 51946
rect 166398 51888 166737 51890
rect 166076 51780 166136 51851
rect 166022 51716 166028 51780
rect 166092 51718 166136 51780
rect 166398 51778 166458 51888
rect 166671 51885 166737 51888
rect 166947 51878 167013 51883
rect 166947 51822 166952 51878
rect 167008 51822 167013 51878
rect 167494 51852 167500 51916
rect 167564 51890 167596 51916
rect 167652 51890 167657 51946
rect 167564 51885 167657 51890
rect 167732 51946 167841 51948
rect 167732 51890 167780 51946
rect 167836 51890 167841 51946
rect 167732 51885 167841 51890
rect 168603 51946 168669 51951
rect 168603 51890 168608 51946
rect 168664 51890 168669 51946
rect 168790 51917 168850 51990
rect 169150 51988 169156 51990
rect 169220 51988 169226 52052
rect 174302 52050 174308 52052
rect 174264 51988 174308 52050
rect 174372 51988 174378 52052
rect 175958 52050 175964 52052
rect 174540 51990 175964 52050
rect 169707 51946 169773 51951
rect 168603 51885 168669 51890
rect 168787 51912 168853 51917
rect 169707 51916 169712 51946
rect 169768 51916 169773 51946
rect 167564 51854 167608 51885
rect 167564 51852 167570 51854
rect 166947 51817 167013 51822
rect 166763 51780 166829 51781
rect 166758 51778 166764 51780
rect 166214 51718 166458 51778
rect 166672 51718 166764 51778
rect 166092 51716 166098 51718
rect 165245 51504 165630 51506
rect 165245 51448 165250 51504
rect 165306 51448 165630 51504
rect 165245 51446 165630 51448
rect 166214 51506 166274 51718
rect 166758 51716 166764 51718
rect 166828 51716 166834 51780
rect 166763 51715 166829 51716
rect 166717 51642 166783 51645
rect 166950 51642 167010 51817
rect 167269 51778 167335 51781
rect 167407 51778 167473 51781
rect 167269 51776 167473 51778
rect 167269 51720 167274 51776
rect 167330 51720 167412 51776
rect 167468 51720 167473 51776
rect 167269 51718 167473 51720
rect 167269 51715 167335 51718
rect 167407 51715 167473 51718
rect 167732 51645 167792 51885
rect 167959 51878 168025 51883
rect 167959 51822 167964 51878
rect 168020 51822 168025 51878
rect 167959 51817 168025 51822
rect 166717 51640 167010 51642
rect 166717 51584 166722 51640
rect 166778 51584 167010 51640
rect 166717 51582 167010 51584
rect 167729 51640 167795 51645
rect 167729 51584 167734 51640
rect 167790 51584 167795 51640
rect 166717 51579 166783 51582
rect 167729 51579 167795 51584
rect 166625 51506 166691 51509
rect 166214 51504 166691 51506
rect 166214 51448 166630 51504
rect 166686 51448 166691 51504
rect 166214 51446 166691 51448
rect 165245 51443 165311 51446
rect 166625 51443 166691 51446
rect 167729 51506 167795 51509
rect 167962 51506 168022 51817
rect 168606 51778 168666 51885
rect 168787 51856 168792 51912
rect 168848 51856 168853 51912
rect 168787 51851 168853 51856
rect 169702 51852 169708 51916
rect 169772 51914 169778 51916
rect 170167 51914 170233 51917
rect 170438 51914 170444 51916
rect 169772 51854 169830 51914
rect 170167 51912 170444 51914
rect 170167 51856 170172 51912
rect 170228 51856 170444 51912
rect 170167 51854 170444 51856
rect 169772 51852 169778 51854
rect 170167 51851 170233 51854
rect 170438 51852 170444 51854
rect 170508 51852 170514 51916
rect 170627 51912 170693 51917
rect 171271 51914 171337 51917
rect 171639 51914 171705 51917
rect 170627 51856 170632 51912
rect 170688 51856 170693 51912
rect 170627 51851 170693 51856
rect 171044 51912 171337 51914
rect 171044 51856 171276 51912
rect 171332 51856 171337 51912
rect 171044 51854 171337 51856
rect 167729 51504 168022 51506
rect 167729 51448 167734 51504
rect 167790 51448 168022 51504
rect 167729 51446 168022 51448
rect 168422 51718 168666 51778
rect 168971 51776 169037 51781
rect 170075 51780 170141 51781
rect 168971 51720 168976 51776
rect 169032 51720 169037 51776
rect 167729 51443 167795 51446
rect 165110 51368 165219 51373
rect 165110 51312 165158 51368
rect 165214 51312 165219 51368
rect 165110 51310 165219 51312
rect 164693 51307 164759 51310
rect 165153 51307 165219 51310
rect 165797 51370 165863 51373
rect 168422 51370 168482 51718
rect 168971 51715 169037 51720
rect 170070 51716 170076 51780
rect 170140 51778 170146 51780
rect 170140 51718 170232 51778
rect 170140 51716 170146 51718
rect 170075 51715 170141 51716
rect 168649 51642 168715 51645
rect 168974 51642 169034 51715
rect 170630 51645 170690 51851
rect 170765 51776 170831 51781
rect 170765 51720 170770 51776
rect 170826 51720 170831 51776
rect 170765 51715 170831 51720
rect 168649 51640 169034 51642
rect 168649 51584 168654 51640
rect 168710 51584 169034 51640
rect 168649 51582 169034 51584
rect 170121 51642 170187 51645
rect 170121 51640 170322 51642
rect 170121 51584 170126 51640
rect 170182 51584 170322 51640
rect 170121 51582 170322 51584
rect 168649 51579 168715 51582
rect 170121 51579 170187 51582
rect 168741 51506 168807 51509
rect 168966 51506 168972 51508
rect 168741 51504 168972 51506
rect 168741 51448 168746 51504
rect 168802 51448 168972 51504
rect 168741 51446 168972 51448
rect 168741 51443 168807 51446
rect 168966 51444 168972 51446
rect 169036 51444 169042 51508
rect 169753 51506 169819 51509
rect 169886 51506 169892 51508
rect 169753 51504 169892 51506
rect 169753 51448 169758 51504
rect 169814 51448 169892 51504
rect 169753 51446 169892 51448
rect 169753 51443 169819 51446
rect 169886 51444 169892 51446
rect 169956 51444 169962 51508
rect 165797 51368 168482 51370
rect 165797 51312 165802 51368
rect 165858 51312 168482 51368
rect 165797 51310 168482 51312
rect 169937 51370 170003 51373
rect 170262 51370 170322 51582
rect 170581 51640 170690 51645
rect 170581 51584 170586 51640
rect 170642 51584 170690 51640
rect 170581 51582 170690 51584
rect 170768 51642 170828 51715
rect 170768 51582 170874 51642
rect 170581 51579 170647 51582
rect 170814 51509 170874 51582
rect 170814 51504 170923 51509
rect 170814 51448 170862 51504
rect 170918 51448 170923 51504
rect 170814 51446 170923 51448
rect 171044 51506 171104 51854
rect 171271 51851 171337 51854
rect 171412 51912 171705 51914
rect 171412 51856 171644 51912
rect 171700 51856 171705 51912
rect 173111 51914 173177 51917
rect 173755 51916 173821 51917
rect 173382 51914 173388 51916
rect 173111 51912 173388 51914
rect 171412 51854 171705 51856
rect 171225 51506 171291 51509
rect 171044 51504 171291 51506
rect 171044 51448 171230 51504
rect 171286 51448 171291 51504
rect 171044 51446 171291 51448
rect 170857 51443 170923 51446
rect 171225 51443 171291 51446
rect 171412 51373 171472 51854
rect 171639 51851 171705 51854
rect 172099 51878 172165 51883
rect 172099 51822 172104 51878
rect 172160 51822 172165 51878
rect 172099 51817 172165 51822
rect 172651 51878 172717 51883
rect 172651 51822 172656 51878
rect 172712 51822 172717 51878
rect 173111 51856 173116 51912
rect 173172 51856 173388 51912
rect 173111 51854 173388 51856
rect 173111 51851 173177 51854
rect 173382 51852 173388 51854
rect 173452 51852 173458 51916
rect 173750 51914 173756 51916
rect 173664 51854 173756 51914
rect 173750 51852 173756 51854
rect 173820 51852 173826 51916
rect 173939 51914 174005 51917
rect 174118 51914 174124 51916
rect 173939 51912 174124 51914
rect 173939 51856 173944 51912
rect 174000 51856 174124 51912
rect 173939 51854 174124 51856
rect 173755 51851 173821 51852
rect 173939 51851 174005 51854
rect 174118 51852 174124 51854
rect 174188 51852 174194 51916
rect 172651 51817 172717 51822
rect 171593 51642 171659 51645
rect 171550 51640 171659 51642
rect 171550 51584 171598 51640
rect 171654 51584 171659 51640
rect 171550 51579 171659 51584
rect 169937 51368 170322 51370
rect 169937 51312 169942 51368
rect 169998 51312 170322 51368
rect 169937 51310 170322 51312
rect 171409 51368 171475 51373
rect 171409 51312 171414 51368
rect 171470 51312 171475 51368
rect 165797 51307 165863 51310
rect 169937 51307 170003 51310
rect 171409 51307 171475 51312
rect 171550 51237 171610 51579
rect 172102 51370 172162 51817
rect 172329 51506 172395 51509
rect 172513 51506 172579 51509
rect 172329 51504 172579 51506
rect 172329 51448 172334 51504
rect 172390 51448 172518 51504
rect 172574 51448 172579 51504
rect 172329 51446 172579 51448
rect 172654 51506 172714 51817
rect 174264 51781 174324 51988
rect 174399 51914 174465 51917
rect 174540 51914 174600 51990
rect 175958 51988 175964 51990
rect 176028 51988 176034 52052
rect 176150 51951 176210 52126
rect 176147 51946 176213 51951
rect 177527 51948 177593 51951
rect 174859 51916 174925 51917
rect 174854 51914 174860 51916
rect 174399 51912 174600 51914
rect 174399 51856 174404 51912
rect 174460 51856 174600 51912
rect 174399 51854 174600 51856
rect 174768 51854 174860 51914
rect 174399 51851 174465 51854
rect 174854 51852 174860 51854
rect 174924 51852 174930 51916
rect 176147 51890 176152 51946
rect 176208 51890 176213 51946
rect 177484 51946 177593 51948
rect 176147 51885 176213 51890
rect 176326 51852 176332 51916
rect 176396 51914 176402 51916
rect 177484 51914 177532 51946
rect 176396 51890 177532 51914
rect 177588 51890 177593 51946
rect 177987 51916 178053 51917
rect 177982 51914 177988 51916
rect 176396 51885 177593 51890
rect 176396 51854 177544 51885
rect 177896 51854 177988 51914
rect 176396 51852 176402 51854
rect 177982 51852 177988 51854
rect 178052 51852 178058 51916
rect 178174 51914 178234 52262
rect 193124 52262 194364 52322
rect 181023 51948 181089 51951
rect 180980 51946 181089 51948
rect 178631 51914 178697 51917
rect 178907 51916 178973 51917
rect 178902 51914 178908 51916
rect 178174 51912 178697 51914
rect 178174 51856 178636 51912
rect 178692 51856 178697 51912
rect 178174 51854 178697 51856
rect 178816 51854 178908 51914
rect 174859 51851 174925 51852
rect 177987 51851 178053 51852
rect 178631 51851 178697 51854
rect 178902 51852 178908 51854
rect 178972 51852 178978 51916
rect 179643 51914 179709 51917
rect 180379 51916 180445 51917
rect 180980 51916 181028 51946
rect 180006 51914 180012 51916
rect 179643 51912 180012 51914
rect 179643 51856 179648 51912
rect 179704 51856 180012 51912
rect 179643 51854 180012 51856
rect 178907 51851 178973 51852
rect 179643 51851 179709 51854
rect 180006 51852 180012 51854
rect 180076 51852 180082 51916
rect 180374 51914 180380 51916
rect 180288 51854 180380 51914
rect 180374 51852 180380 51854
rect 180444 51852 180450 51916
rect 180926 51852 180932 51916
rect 180996 51890 181028 51916
rect 181084 51890 181089 51946
rect 181299 51946 181365 51951
rect 181299 51916 181304 51946
rect 181360 51916 181365 51946
rect 182403 51946 182469 51951
rect 180996 51885 181089 51890
rect 180996 51854 181040 51885
rect 180996 51852 181002 51854
rect 181294 51852 181300 51916
rect 181364 51914 181370 51916
rect 181364 51854 181422 51914
rect 182403 51890 182408 51946
rect 182464 51914 182469 51946
rect 182955 51946 183021 51951
rect 182955 51916 182960 51946
rect 183016 51916 183021 51946
rect 192523 51946 192589 51951
rect 182766 51914 182772 51916
rect 182464 51890 182772 51914
rect 182403 51885 182772 51890
rect 182406 51854 182772 51885
rect 181364 51852 181370 51854
rect 182766 51852 182772 51854
rect 182836 51852 182842 51916
rect 182950 51852 182956 51916
rect 183020 51914 183026 51916
rect 183599 51914 183665 51917
rect 183870 51914 183876 51916
rect 183020 51854 183078 51914
rect 183599 51912 183876 51914
rect 183599 51856 183604 51912
rect 183660 51856 183876 51912
rect 183599 51854 183876 51856
rect 183020 51852 183026 51854
rect 180379 51851 180445 51852
rect 183599 51851 183665 51854
rect 183870 51852 183876 51854
rect 183940 51852 183946 51916
rect 184151 51914 184217 51917
rect 184611 51916 184677 51917
rect 184422 51914 184428 51916
rect 184151 51912 184428 51914
rect 184151 51856 184156 51912
rect 184212 51856 184428 51912
rect 184151 51854 184428 51856
rect 184151 51851 184217 51854
rect 184422 51852 184428 51854
rect 184492 51852 184498 51916
rect 184606 51852 184612 51916
rect 184676 51914 184682 51916
rect 184676 51854 184768 51914
rect 184676 51852 184682 51854
rect 185342 51852 185348 51916
rect 185412 51914 185418 51916
rect 185623 51914 185689 51917
rect 187003 51916 187069 51917
rect 186998 51914 187004 51916
rect 185412 51912 185689 51914
rect 185412 51856 185628 51912
rect 185684 51856 185689 51912
rect 185412 51854 185689 51856
rect 186912 51854 187004 51914
rect 185412 51852 185418 51854
rect 184611 51851 184677 51852
rect 185623 51851 185689 51854
rect 186998 51852 187004 51854
rect 187068 51852 187074 51916
rect 188470 51852 188476 51916
rect 188540 51914 188546 51916
rect 188843 51914 188909 51917
rect 188540 51912 188909 51914
rect 188540 51856 188848 51912
rect 188904 51856 188909 51912
rect 188540 51854 188909 51856
rect 188540 51852 188546 51854
rect 187003 51851 187069 51852
rect 188843 51851 188909 51854
rect 189022 51852 189028 51916
rect 189092 51914 189098 51916
rect 192523 51914 192528 51946
rect 189092 51890 192528 51914
rect 192584 51890 192589 51946
rect 189092 51885 192589 51890
rect 189092 51854 192586 51885
rect 189092 51852 189098 51854
rect 192702 51852 192708 51916
rect 192772 51914 192778 51916
rect 192891 51914 192957 51917
rect 192772 51912 192957 51914
rect 192772 51856 192896 51912
rect 192952 51856 192957 51912
rect 192772 51854 192957 51856
rect 193124 51914 193184 52262
rect 194358 52260 194364 52262
rect 194428 52260 194434 52324
rect 194542 52260 194548 52324
rect 194612 52322 194618 52324
rect 194910 52322 194916 52324
rect 194612 52262 194916 52322
rect 194612 52260 194618 52262
rect 194910 52260 194916 52262
rect 194980 52260 194986 52324
rect 208710 52322 208716 52324
rect 204670 52262 208716 52322
rect 193806 52186 193812 52188
rect 193538 52126 193812 52186
rect 193538 51951 193598 52126
rect 193806 52124 193812 52126
rect 193876 52124 193882 52188
rect 194726 52124 194732 52188
rect 194796 52186 194802 52188
rect 194796 52126 195530 52186
rect 194796 52124 194802 52126
rect 194542 51988 194548 52052
rect 194612 52050 194618 52052
rect 194612 51990 194886 52050
rect 194612 51988 194618 51990
rect 193535 51946 193601 51951
rect 193351 51914 193417 51917
rect 193124 51912 193417 51914
rect 193124 51856 193356 51912
rect 193412 51856 193417 51912
rect 193535 51890 193540 51946
rect 193596 51890 193601 51946
rect 194826 51917 194886 51990
rect 195470 51951 195530 52126
rect 196198 51988 196204 52052
rect 196268 52050 196274 52052
rect 204670 52050 204730 52262
rect 208710 52260 208716 52262
rect 208780 52260 208786 52324
rect 204846 52124 204852 52188
rect 204916 52186 204922 52188
rect 204916 52126 205282 52186
rect 204916 52124 204922 52126
rect 196268 51990 196818 52050
rect 196268 51988 196274 51990
rect 195467 51946 195533 51951
rect 193535 51885 193601 51890
rect 193903 51914 193969 51917
rect 194174 51914 194180 51916
rect 193903 51912 194180 51914
rect 193124 51854 193417 51856
rect 192772 51852 192778 51854
rect 192891 51851 192957 51854
rect 193351 51851 193417 51854
rect 193903 51856 193908 51912
rect 193964 51856 194180 51912
rect 193903 51854 194180 51856
rect 193903 51851 193969 51854
rect 194174 51852 194180 51854
rect 194244 51852 194250 51916
rect 194823 51912 194889 51917
rect 195099 51916 195165 51917
rect 195094 51914 195100 51916
rect 194823 51856 194828 51912
rect 194884 51856 194889 51912
rect 194823 51851 194889 51856
rect 195008 51854 195100 51914
rect 195094 51852 195100 51854
rect 195164 51852 195170 51916
rect 195467 51890 195472 51946
rect 195528 51890 195533 51946
rect 195835 51946 195901 51951
rect 195467 51885 195533 51890
rect 195646 51852 195652 51916
rect 195716 51914 195722 51916
rect 195835 51914 195840 51946
rect 195716 51890 195840 51914
rect 195896 51890 195901 51946
rect 195716 51885 195901 51890
rect 195716 51854 195898 51885
rect 195716 51852 195722 51854
rect 196382 51852 196388 51916
rect 196452 51914 196458 51916
rect 196571 51914 196637 51917
rect 196452 51912 196637 51914
rect 196452 51856 196576 51912
rect 196632 51856 196637 51912
rect 196452 51854 196637 51856
rect 196758 51914 196818 51990
rect 201864 51990 204730 52050
rect 201864 51951 201924 51990
rect 205222 51951 205282 52126
rect 205582 52124 205588 52188
rect 205652 52186 205658 52188
rect 218697 52186 218763 52189
rect 205652 52184 218763 52186
rect 205652 52128 218702 52184
rect 218758 52128 218763 52184
rect 205652 52126 218763 52128
rect 205652 52124 205658 52126
rect 218697 52123 218763 52126
rect 207238 51988 207244 52052
rect 207308 52050 207314 52052
rect 207308 51990 208364 52050
rect 207308 51988 207314 51990
rect 198595 51946 198661 51951
rect 197123 51914 197189 51917
rect 196758 51912 197189 51914
rect 196758 51856 197128 51912
rect 197184 51856 197189 51912
rect 196758 51854 197189 51856
rect 196452 51852 196458 51854
rect 195099 51851 195165 51852
rect 196571 51851 196637 51854
rect 197123 51851 197189 51854
rect 198222 51852 198228 51916
rect 198292 51914 198298 51916
rect 198411 51914 198477 51917
rect 198595 51916 198600 51946
rect 198656 51916 198661 51946
rect 201815 51946 201924 51951
rect 198292 51912 198477 51914
rect 198292 51856 198416 51912
rect 198472 51856 198477 51912
rect 198292 51854 198477 51856
rect 198292 51852 198298 51854
rect 198411 51851 198477 51854
rect 198590 51852 198596 51916
rect 198660 51914 198666 51916
rect 198660 51854 198718 51914
rect 198660 51852 198666 51854
rect 200062 51852 200068 51916
rect 200132 51914 200138 51916
rect 201263 51914 201329 51917
rect 200132 51912 201329 51914
rect 200132 51856 201268 51912
rect 201324 51856 201329 51912
rect 201815 51890 201820 51946
rect 201876 51890 201924 51946
rect 205219 51946 205285 51951
rect 201815 51888 201924 51890
rect 201815 51885 201881 51888
rect 200132 51854 201329 51856
rect 200132 51852 200138 51854
rect 201263 51851 201329 51854
rect 202086 51852 202092 51916
rect 202156 51914 202162 51916
rect 202367 51914 202433 51917
rect 202156 51912 202433 51914
rect 202156 51856 202372 51912
rect 202428 51856 202433 51912
rect 202156 51854 202433 51856
rect 202156 51852 202162 51854
rect 202367 51851 202433 51854
rect 203374 51852 203380 51916
rect 203444 51914 203450 51916
rect 204115 51914 204181 51917
rect 203444 51912 204181 51914
rect 203444 51856 204120 51912
rect 204176 51856 204181 51912
rect 203444 51854 204181 51856
rect 203444 51852 203450 51854
rect 204115 51851 204181 51854
rect 204483 51914 204549 51917
rect 205030 51914 205036 51916
rect 204483 51912 205036 51914
rect 204483 51856 204488 51912
rect 204544 51856 205036 51912
rect 204483 51854 205036 51856
rect 204483 51851 204549 51854
rect 205030 51852 205036 51854
rect 205100 51852 205106 51916
rect 205219 51890 205224 51946
rect 205280 51890 205285 51946
rect 205403 51916 205469 51917
rect 205219 51885 205285 51890
rect 205398 51852 205404 51916
rect 205468 51914 205474 51916
rect 205468 51854 205560 51914
rect 205766 51886 205772 51950
rect 205836 51948 205842 51950
rect 206139 51948 206205 51951
rect 205836 51946 206205 51948
rect 205836 51890 206144 51946
rect 206200 51890 206205 51946
rect 206323 51946 206389 51951
rect 206323 51916 206328 51946
rect 206384 51916 206389 51946
rect 206875 51946 206941 51951
rect 205836 51888 206205 51890
rect 205836 51886 205842 51888
rect 206139 51885 206205 51888
rect 205468 51852 205474 51854
rect 206318 51852 206324 51916
rect 206388 51914 206394 51916
rect 206388 51854 206446 51914
rect 206388 51852 206394 51854
rect 206686 51852 206692 51916
rect 206756 51914 206762 51916
rect 206875 51914 206880 51946
rect 206756 51890 206880 51914
rect 206936 51890 206941 51946
rect 207059 51916 207125 51917
rect 206756 51885 206941 51890
rect 206756 51854 206938 51885
rect 206756 51852 206762 51854
rect 207054 51852 207060 51916
rect 207124 51914 207130 51916
rect 207124 51854 207216 51914
rect 207124 51852 207130 51854
rect 207422 51852 207428 51916
rect 207492 51914 207498 51916
rect 208163 51914 208229 51917
rect 207492 51912 208229 51914
rect 207492 51856 208168 51912
rect 208224 51856 208229 51912
rect 207492 51854 208229 51856
rect 207492 51852 207498 51854
rect 205403 51851 205469 51852
rect 207059 51851 207125 51852
rect 208163 51851 208229 51854
rect 173014 51716 173020 51780
rect 173084 51778 173090 51780
rect 173847 51778 173913 51781
rect 173084 51776 173913 51778
rect 173084 51720 173852 51776
rect 173908 51720 173913 51776
rect 173084 51718 173913 51720
rect 173084 51716 173090 51718
rect 173847 51715 173913 51718
rect 174215 51776 174324 51781
rect 174445 51780 174511 51781
rect 174445 51778 174492 51780
rect 174215 51720 174220 51776
rect 174276 51720 174324 51776
rect 174215 51718 174324 51720
rect 174400 51776 174492 51778
rect 174400 51720 174450 51776
rect 174400 51718 174492 51720
rect 174215 51715 174281 51718
rect 174445 51716 174492 51718
rect 174556 51716 174562 51780
rect 174629 51778 174695 51781
rect 175406 51778 175412 51780
rect 174629 51776 175412 51778
rect 174629 51720 174634 51776
rect 174690 51720 175412 51776
rect 174629 51718 175412 51720
rect 174445 51715 174511 51716
rect 174629 51715 174695 51718
rect 175406 51716 175412 51718
rect 175476 51716 175482 51780
rect 175641 51778 175707 51781
rect 176101 51778 176167 51781
rect 175641 51776 176167 51778
rect 175641 51720 175646 51776
rect 175702 51720 176106 51776
rect 176162 51720 176167 51776
rect 175641 51718 176167 51720
rect 175641 51715 175707 51718
rect 176101 51715 176167 51718
rect 178953 51778 179019 51781
rect 205582 51778 205588 51780
rect 178953 51776 205588 51778
rect 178953 51720 178958 51776
rect 179014 51720 205588 51776
rect 178953 51718 205588 51720
rect 178953 51715 179019 51718
rect 205582 51716 205588 51718
rect 205652 51716 205658 51780
rect 206502 51716 206508 51780
rect 206572 51778 206578 51780
rect 207335 51778 207401 51781
rect 207611 51780 207677 51781
rect 207606 51778 207612 51780
rect 206572 51776 207401 51778
rect 206572 51720 207340 51776
rect 207396 51720 207401 51776
rect 206572 51718 207401 51720
rect 207520 51718 207612 51778
rect 206572 51716 206578 51718
rect 207335 51715 207401 51718
rect 207606 51716 207612 51718
rect 207676 51716 207682 51780
rect 208071 51778 208137 51781
rect 208304 51778 208364 51990
rect 209078 51988 209084 52052
rect 209148 52050 209154 52052
rect 209148 51990 209652 52050
rect 209148 51988 209154 51990
rect 209592 51951 209652 51990
rect 209592 51946 209701 51951
rect 208991 51914 209057 51917
rect 209267 51916 209333 51917
rect 209262 51914 209268 51916
rect 208948 51912 209057 51914
rect 208948 51856 208996 51912
rect 209052 51856 209057 51912
rect 208948 51851 209057 51856
rect 209176 51854 209268 51914
rect 209262 51852 209268 51854
rect 209332 51852 209338 51916
rect 209446 51914 209452 51916
rect 209408 51852 209452 51914
rect 209516 51852 209522 51916
rect 209592 51890 209640 51946
rect 209696 51890 209701 51946
rect 211107 51946 211173 51951
rect 209592 51888 209701 51890
rect 209635 51885 209701 51888
rect 210279 51914 210345 51917
rect 210555 51916 210621 51917
rect 210923 51916 210989 51917
rect 210279 51912 210388 51914
rect 210279 51856 210284 51912
rect 210340 51856 210388 51912
rect 209267 51851 209333 51852
rect 208948 51781 209008 51851
rect 208071 51776 208364 51778
rect 208071 51720 208076 51776
rect 208132 51720 208364 51776
rect 208071 51718 208364 51720
rect 208945 51776 209011 51781
rect 208945 51720 208950 51776
rect 209006 51720 209011 51776
rect 207611 51715 207677 51716
rect 208071 51715 208137 51718
rect 208945 51715 209011 51720
rect 209408 51778 209468 51852
rect 210279 51851 210388 51856
rect 210550 51852 210556 51916
rect 210620 51914 210626 51916
rect 210918 51914 210924 51916
rect 210620 51854 210712 51914
rect 210832 51854 210924 51914
rect 210620 51852 210626 51854
rect 210918 51852 210924 51854
rect 210988 51852 210994 51916
rect 211107 51890 211112 51946
rect 211168 51890 211173 51946
rect 212303 51946 212369 51951
rect 211107 51885 211173 51890
rect 210555 51851 210621 51852
rect 210923 51851 210989 51852
rect 209543 51778 209609 51781
rect 209408 51776 209609 51778
rect 209408 51720 209548 51776
rect 209604 51720 209609 51776
rect 209408 51718 209609 51720
rect 209543 51715 209609 51718
rect 210182 51716 210188 51780
rect 210252 51778 210258 51780
rect 210328 51778 210388 51851
rect 210252 51718 210388 51778
rect 210252 51716 210258 51718
rect 210550 51716 210556 51780
rect 210620 51778 210626 51780
rect 211110 51778 211170 51885
rect 212022 51852 212028 51916
rect 212092 51914 212098 51916
rect 212303 51914 212308 51946
rect 212092 51890 212308 51914
rect 212364 51890 212369 51946
rect 214787 51946 214853 51951
rect 212487 51914 212553 51917
rect 212092 51885 212369 51890
rect 212444 51912 212553 51914
rect 212092 51854 212366 51885
rect 212444 51856 212492 51912
rect 212548 51856 212553 51912
rect 212092 51852 212098 51854
rect 212444 51851 212553 51856
rect 213315 51912 213381 51917
rect 213315 51856 213320 51912
rect 213376 51856 213381 51912
rect 213315 51851 213381 51856
rect 213494 51852 213500 51916
rect 213564 51914 213570 51916
rect 213867 51914 213933 51917
rect 213564 51912 213933 51914
rect 213564 51856 213872 51912
rect 213928 51856 213933 51912
rect 213564 51854 213933 51856
rect 213564 51852 213570 51854
rect 213867 51851 213933 51854
rect 214046 51852 214052 51916
rect 214116 51914 214122 51916
rect 214787 51914 214792 51946
rect 214116 51890 214792 51914
rect 214848 51890 214853 51946
rect 215523 51946 215589 51951
rect 215523 51916 215528 51946
rect 215584 51916 215589 51946
rect 214116 51885 214853 51890
rect 214116 51854 214850 51885
rect 214116 51852 214122 51854
rect 215518 51852 215524 51916
rect 215588 51914 215594 51916
rect 215588 51854 215646 51914
rect 215588 51852 215594 51854
rect 211659 51780 211725 51781
rect 212211 51780 212277 51781
rect 212444 51780 212504 51851
rect 211654 51778 211660 51780
rect 210620 51718 211170 51778
rect 211568 51718 211660 51778
rect 210620 51716 210626 51718
rect 211654 51716 211660 51718
rect 211724 51716 211730 51780
rect 212206 51778 212212 51780
rect 212120 51718 212212 51778
rect 212206 51716 212212 51718
rect 212276 51716 212282 51780
rect 212390 51716 212396 51780
rect 212460 51718 212504 51780
rect 213318 51781 213378 51851
rect 213318 51776 213427 51781
rect 213318 51720 213366 51776
rect 213422 51720 213427 51776
rect 213318 51718 213427 51720
rect 212460 51716 212466 51718
rect 211659 51715 211725 51716
rect 212211 51715 212277 51716
rect 213361 51715 213427 51718
rect 213683 51778 213749 51781
rect 213821 51778 213887 51781
rect 213683 51776 213887 51778
rect 213683 51720 213688 51776
rect 213744 51720 213826 51776
rect 213882 51720 213887 51776
rect 213683 51718 213887 51720
rect 213683 51715 213749 51718
rect 213821 51715 213887 51718
rect 214230 51716 214236 51780
rect 214300 51778 214306 51780
rect 214695 51778 214761 51781
rect 214300 51776 214761 51778
rect 214300 51720 214700 51776
rect 214756 51720 214761 51776
rect 214300 51718 214761 51720
rect 214300 51716 214306 51718
rect 214695 51715 214761 51718
rect 173198 51580 173204 51644
rect 173268 51642 173274 51644
rect 221549 51642 221615 51645
rect 173268 51640 221615 51642
rect 173268 51584 221554 51640
rect 221610 51584 221615 51640
rect 173268 51582 221615 51584
rect 173268 51580 173274 51582
rect 221549 51579 221615 51582
rect 172789 51506 172855 51509
rect 172654 51504 172855 51506
rect 172654 51448 172794 51504
rect 172850 51448 172855 51504
rect 172654 51446 172855 51448
rect 172329 51443 172395 51446
rect 172513 51443 172579 51446
rect 172789 51443 172855 51446
rect 173566 51444 173572 51508
rect 173636 51506 173642 51508
rect 173801 51506 173867 51509
rect 177757 51506 177823 51509
rect 173636 51504 173867 51506
rect 173636 51448 173806 51504
rect 173862 51448 173867 51504
rect 173636 51446 173867 51448
rect 173636 51444 173642 51446
rect 173801 51443 173867 51446
rect 173942 51504 177823 51506
rect 173942 51448 177762 51504
rect 177818 51448 177823 51504
rect 173942 51446 177823 51448
rect 172329 51370 172395 51373
rect 172102 51368 172395 51370
rect 172102 51312 172334 51368
rect 172390 51312 172395 51368
rect 172102 51310 172395 51312
rect 172329 51307 172395 51310
rect 173065 51370 173131 51373
rect 173198 51370 173204 51372
rect 173065 51368 173204 51370
rect 173065 51312 173070 51368
rect 173126 51312 173204 51368
rect 173065 51310 173204 51312
rect 173065 51307 173131 51310
rect 173198 51308 173204 51310
rect 173268 51308 173274 51372
rect 171501 51232 171610 51237
rect 171501 51176 171506 51232
rect 171562 51176 171610 51232
rect 171501 51174 171610 51176
rect 171501 51171 171567 51174
rect 159357 51098 159423 51101
rect 162853 51098 162919 51101
rect 159357 51096 162919 51098
rect 159357 51040 159362 51096
rect 159418 51040 162858 51096
rect 162914 51040 162919 51096
rect 159357 51038 162919 51040
rect 159357 51035 159423 51038
rect 162853 51035 162919 51038
rect 170121 51098 170187 51101
rect 173942 51098 174002 51446
rect 177757 51443 177823 51446
rect 178861 51506 178927 51509
rect 232497 51506 232563 51509
rect 178861 51504 232563 51506
rect 178861 51448 178866 51504
rect 178922 51448 232502 51504
rect 232558 51448 232563 51504
rect 178861 51446 232563 51448
rect 178861 51443 178927 51446
rect 232497 51443 232563 51446
rect 256693 51506 256759 51509
rect 256693 51504 260084 51506
rect 256693 51448 256698 51504
rect 256754 51448 260084 51504
rect 256693 51446 260084 51448
rect 256693 51443 256759 51446
rect 174169 51370 174235 51373
rect 240961 51370 241027 51373
rect 174169 51368 241027 51370
rect 174169 51312 174174 51368
rect 174230 51312 240966 51368
rect 241022 51312 241027 51368
rect 174169 51310 241027 51312
rect 174169 51307 174235 51310
rect 240961 51307 241027 51310
rect 174486 51172 174492 51236
rect 174556 51234 174562 51236
rect 179137 51234 179203 51237
rect 240777 51234 240843 51237
rect 174556 51174 178970 51234
rect 174556 51172 174562 51174
rect 170121 51096 174002 51098
rect 170121 51040 170126 51096
rect 170182 51040 174002 51096
rect 170121 51038 174002 51040
rect 170121 51035 170187 51038
rect 174854 51036 174860 51100
rect 174924 51098 174930 51100
rect 175273 51098 175339 51101
rect 174924 51096 175339 51098
rect 174924 51040 175278 51096
rect 175334 51040 175339 51096
rect 174924 51038 175339 51040
rect 174924 51036 174930 51038
rect 175273 51035 175339 51038
rect 175406 51036 175412 51100
rect 175476 51098 175482 51100
rect 178769 51098 178835 51101
rect 175476 51096 178835 51098
rect 175476 51040 178774 51096
rect 178830 51040 178835 51096
rect 175476 51038 178835 51040
rect 178910 51098 178970 51174
rect 179137 51232 240843 51234
rect 179137 51176 179142 51232
rect 179198 51176 240782 51232
rect 240838 51176 240843 51232
rect 179137 51174 240843 51176
rect 179137 51171 179203 51174
rect 240777 51171 240843 51174
rect 253289 51098 253355 51101
rect 178910 51096 253355 51098
rect 178910 51040 253294 51096
rect 253350 51040 253355 51096
rect 178910 51038 253355 51040
rect 175476 51036 175482 51038
rect 178769 51035 178835 51038
rect 253289 51035 253355 51038
rect 135345 50962 135411 50965
rect 133830 50960 135411 50962
rect 133830 50904 135350 50960
rect 135406 50904 135411 50960
rect 133830 50902 135411 50904
rect 133830 50592 133890 50902
rect 135345 50899 135411 50902
rect 173382 50900 173388 50964
rect 173452 50962 173458 50964
rect 249241 50962 249307 50965
rect 173452 50960 249307 50962
rect 173452 50904 249246 50960
rect 249302 50904 249307 50960
rect 173452 50902 249307 50904
rect 173452 50900 173458 50902
rect 249241 50899 249307 50902
rect 170806 50764 170812 50828
rect 170876 50826 170882 50828
rect 171041 50826 171107 50829
rect 170876 50824 171107 50826
rect 170876 50768 171046 50824
rect 171102 50768 171107 50824
rect 170876 50766 171107 50768
rect 170876 50764 170882 50766
rect 171041 50763 171107 50766
rect 174353 50826 174419 50829
rect 249057 50826 249123 50829
rect 174353 50824 249123 50826
rect 174353 50768 174358 50824
rect 174414 50768 249062 50824
rect 249118 50768 249123 50824
rect 174353 50766 249123 50768
rect 174353 50763 174419 50766
rect 249057 50763 249123 50766
rect 173750 50628 173756 50692
rect 173820 50690 173826 50692
rect 239397 50690 239463 50693
rect 173820 50688 239463 50690
rect 173820 50632 239402 50688
rect 239458 50632 239463 50688
rect 173820 50630 239463 50632
rect 173820 50628 173826 50630
rect 239397 50627 239463 50630
rect 172881 50554 172947 50557
rect 234061 50554 234127 50557
rect 172881 50552 234127 50554
rect 172881 50496 172886 50552
rect 172942 50496 234066 50552
rect 234122 50496 234127 50552
rect 172881 50494 234127 50496
rect 172881 50491 172947 50494
rect 234061 50491 234127 50494
rect 175958 50356 175964 50420
rect 176028 50418 176034 50420
rect 233877 50418 233943 50421
rect 176028 50416 233943 50418
rect 176028 50360 233882 50416
rect 233938 50360 233943 50416
rect 176028 50358 233943 50360
rect 176028 50356 176034 50358
rect 233877 50355 233943 50358
rect 169661 50284 169727 50285
rect 169661 50282 169708 50284
rect 169616 50280 169708 50282
rect 169616 50224 169666 50280
rect 169616 50222 169708 50224
rect 169661 50220 169708 50222
rect 169772 50220 169778 50284
rect 170622 50220 170628 50284
rect 170692 50282 170698 50284
rect 170765 50282 170831 50285
rect 170692 50280 170831 50282
rect 170692 50224 170770 50280
rect 170826 50224 170831 50280
rect 170692 50222 170831 50224
rect 170692 50220 170698 50222
rect 169661 50219 169727 50220
rect 170765 50219 170831 50222
rect 173014 50220 173020 50284
rect 173084 50282 173090 50284
rect 221457 50282 221523 50285
rect 173084 50280 221523 50282
rect 173084 50224 221462 50280
rect 221518 50224 221523 50280
rect 173084 50222 221523 50224
rect 173084 50220 173090 50222
rect 221457 50219 221523 50222
rect 158069 50146 158135 50149
rect 176469 50146 176535 50149
rect 158069 50144 176535 50146
rect 158069 50088 158074 50144
rect 158130 50088 176474 50144
rect 176530 50088 176535 50144
rect 158069 50086 176535 50088
rect 158069 50083 158135 50086
rect 176469 50083 176535 50086
rect 177757 50146 177823 50149
rect 178902 50146 178908 50148
rect 177757 50144 178908 50146
rect 177757 50088 177762 50144
rect 177818 50088 178908 50144
rect 177757 50086 178908 50088
rect 177757 50083 177823 50086
rect 178902 50084 178908 50086
rect 178972 50084 178978 50148
rect 186497 50146 186563 50149
rect 186998 50146 187004 50148
rect 186497 50144 187004 50146
rect 186497 50088 186502 50144
rect 186558 50088 187004 50144
rect 186497 50086 187004 50088
rect 186497 50083 186563 50086
rect 186998 50084 187004 50086
rect 187068 50084 187074 50148
rect 191414 50084 191420 50148
rect 191484 50146 191490 50148
rect 191741 50146 191807 50149
rect 191484 50144 191807 50146
rect 191484 50088 191746 50144
rect 191802 50088 191807 50144
rect 191484 50086 191807 50088
rect 191484 50084 191490 50086
rect 191741 50083 191807 50086
rect 193990 50084 193996 50148
rect 194060 50146 194066 50148
rect 194225 50146 194291 50149
rect 194060 50144 194291 50146
rect 194060 50088 194230 50144
rect 194286 50088 194291 50144
rect 194060 50086 194291 50088
rect 194060 50084 194066 50086
rect 194225 50083 194291 50086
rect 203558 50084 203564 50148
rect 203628 50146 203634 50148
rect 204161 50146 204227 50149
rect 203628 50144 204227 50146
rect 203628 50088 204166 50144
rect 204222 50088 204227 50144
rect 203628 50086 204227 50088
rect 203628 50084 203634 50086
rect 204161 50083 204227 50086
rect 204529 50146 204595 50149
rect 205449 50148 205515 50149
rect 205030 50146 205036 50148
rect 204529 50144 205036 50146
rect 204529 50088 204534 50144
rect 204590 50088 205036 50144
rect 204529 50086 205036 50088
rect 204529 50083 204595 50086
rect 205030 50084 205036 50086
rect 205100 50084 205106 50148
rect 205398 50146 205404 50148
rect 205358 50086 205404 50146
rect 205468 50144 205515 50148
rect 205510 50088 205515 50144
rect 205398 50084 205404 50086
rect 205468 50084 205515 50088
rect 206502 50084 206508 50148
rect 206572 50146 206578 50148
rect 206921 50146 206987 50149
rect 206572 50144 206987 50146
rect 206572 50088 206926 50144
rect 206982 50088 206987 50144
rect 206572 50086 206987 50088
rect 206572 50084 206578 50086
rect 205449 50083 205515 50084
rect 206921 50083 206987 50086
rect 207054 50084 207060 50148
rect 207124 50146 207130 50148
rect 207381 50146 207447 50149
rect 207124 50144 207447 50146
rect 207124 50088 207386 50144
rect 207442 50088 207447 50144
rect 207124 50086 207447 50088
rect 207124 50084 207130 50086
rect 207381 50083 207447 50086
rect 207606 50084 207612 50148
rect 207676 50146 207682 50148
rect 208301 50146 208367 50149
rect 209313 50148 209379 50149
rect 207676 50144 208367 50146
rect 207676 50088 208306 50144
rect 208362 50088 208367 50144
rect 207676 50086 208367 50088
rect 207676 50084 207682 50086
rect 208301 50083 208367 50086
rect 209262 50084 209268 50148
rect 209332 50146 209379 50148
rect 209589 50148 209655 50149
rect 209332 50144 209424 50146
rect 209374 50088 209424 50144
rect 209332 50086 209424 50088
rect 209589 50144 209636 50148
rect 209700 50146 209706 50148
rect 209589 50088 209594 50144
rect 209332 50084 209379 50086
rect 209313 50083 209379 50084
rect 209589 50084 209636 50088
rect 209700 50086 209746 50146
rect 209700 50084 209706 50086
rect 210366 50084 210372 50148
rect 210436 50146 210442 50148
rect 211061 50146 211127 50149
rect 210436 50144 211127 50146
rect 210436 50088 211066 50144
rect 211122 50088 211127 50144
rect 210436 50086 211127 50088
rect 210436 50084 210442 50086
rect 209589 50083 209655 50084
rect 211061 50083 211127 50086
rect 211337 50146 211403 50149
rect 258574 50146 258580 50148
rect 211337 50144 258580 50146
rect 211337 50088 211342 50144
rect 211398 50088 258580 50144
rect 211337 50086 258580 50088
rect 211337 50083 211403 50086
rect 258574 50084 258580 50086
rect 258644 50084 258650 50148
rect 173985 50010 174051 50013
rect 174261 50012 174327 50013
rect 174118 50010 174124 50012
rect 173985 50008 174124 50010
rect 173985 49952 173990 50008
rect 174046 49952 174124 50008
rect 173985 49950 174124 49952
rect 173985 49947 174051 49950
rect 174118 49948 174124 49950
rect 174188 49948 174194 50012
rect 174261 50008 174308 50012
rect 174372 50010 174378 50012
rect 177757 50010 177823 50013
rect 177982 50010 177988 50012
rect 174261 49952 174266 50008
rect 174261 49948 174308 49952
rect 174372 49950 174418 50010
rect 177757 50008 177988 50010
rect 177757 49952 177762 50008
rect 177818 49952 177988 50008
rect 177757 49950 177988 49952
rect 174372 49948 174378 49950
rect 174261 49947 174327 49948
rect 177757 49947 177823 49950
rect 177982 49948 177988 49950
rect 178052 49948 178058 50012
rect 189257 50010 189323 50013
rect 190126 50010 190132 50012
rect 189257 50008 190132 50010
rect 189257 49952 189262 50008
rect 189318 49952 190132 50008
rect 189257 49950 190132 49952
rect 189257 49947 189323 49950
rect 190126 49948 190132 49950
rect 190196 49948 190202 50012
rect 191046 49948 191052 50012
rect 191116 50010 191122 50012
rect 191373 50010 191439 50013
rect 191649 50012 191715 50013
rect 191598 50010 191604 50012
rect 191116 50008 191439 50010
rect 191116 49952 191378 50008
rect 191434 49952 191439 50008
rect 191116 49950 191439 49952
rect 191558 49950 191604 50010
rect 191668 50008 191715 50012
rect 191710 49952 191715 50008
rect 191116 49948 191122 49950
rect 191373 49947 191439 49950
rect 191598 49948 191604 49950
rect 191668 49948 191715 49952
rect 191649 49947 191715 49948
rect 193857 50010 193923 50013
rect 194174 50010 194180 50012
rect 193857 50008 194180 50010
rect 193857 49952 193862 50008
rect 193918 49952 194180 50008
rect 193857 49950 194180 49952
rect 193857 49947 193923 49950
rect 194174 49948 194180 49950
rect 194244 49948 194250 50012
rect 205950 49948 205956 50012
rect 206020 50010 206026 50012
rect 206185 50010 206251 50013
rect 206020 50008 206251 50010
rect 206020 49952 206190 50008
rect 206246 49952 206251 50008
rect 206020 49950 206251 49952
rect 206020 49948 206026 49950
rect 206185 49947 206251 49950
rect 206829 50010 206895 50013
rect 206829 50008 208594 50010
rect 206829 49952 206834 50008
rect 206890 49952 208594 50008
rect 206829 49950 208594 49952
rect 206829 49947 206895 49950
rect 191230 49812 191236 49876
rect 191300 49874 191306 49876
rect 191465 49874 191531 49877
rect 204897 49876 204963 49877
rect 191300 49872 191531 49874
rect 191300 49816 191470 49872
rect 191526 49816 191531 49872
rect 191300 49814 191531 49816
rect 191300 49812 191306 49814
rect 191465 49811 191531 49814
rect 204846 49812 204852 49876
rect 204916 49874 204963 49876
rect 204916 49872 205008 49874
rect 204958 49816 205008 49872
rect 204916 49814 205008 49816
rect 204916 49812 204963 49814
rect 207422 49812 207428 49876
rect 207492 49874 207498 49876
rect 208025 49874 208091 49877
rect 207492 49872 208091 49874
rect 207492 49816 208030 49872
rect 208086 49816 208091 49872
rect 207492 49814 208091 49816
rect 208534 49874 208594 49950
rect 209262 49948 209268 50012
rect 209332 50010 209338 50012
rect 209773 50010 209839 50013
rect 209332 50008 209839 50010
rect 209332 49952 209778 50008
rect 209834 49952 209839 50008
rect 209332 49950 209839 49952
rect 209332 49948 209338 49950
rect 209773 49947 209839 49950
rect 213494 49948 213500 50012
rect 213564 50010 213570 50012
rect 213637 50010 213703 50013
rect 213564 50008 213703 50010
rect 213564 49952 213642 50008
rect 213698 49952 213703 50008
rect 213564 49950 213703 49952
rect 213564 49948 213570 49950
rect 213637 49947 213703 49950
rect 216397 49874 216463 49877
rect 208534 49872 216463 49874
rect 208534 49816 216402 49872
rect 216458 49816 216463 49872
rect 208534 49814 216463 49816
rect 207492 49812 207498 49814
rect 204897 49811 204963 49812
rect 208025 49811 208091 49814
rect 216397 49811 216463 49814
rect 182449 49738 182515 49741
rect 183921 49740 183987 49741
rect 182950 49738 182956 49740
rect 182449 49736 182956 49738
rect 182449 49680 182454 49736
rect 182510 49680 182956 49736
rect 182449 49678 182956 49680
rect 182449 49675 182515 49678
rect 182950 49676 182956 49678
rect 183020 49676 183026 49740
rect 183870 49738 183876 49740
rect 183830 49678 183876 49738
rect 183940 49736 183987 49740
rect 183982 49680 183987 49736
rect 183870 49676 183876 49678
rect 183940 49676 183987 49680
rect 194358 49676 194364 49740
rect 194428 49738 194434 49740
rect 195697 49738 195763 49741
rect 196341 49740 196407 49741
rect 202045 49740 202111 49741
rect 196341 49738 196388 49740
rect 194428 49736 195763 49738
rect 194428 49680 195702 49736
rect 195758 49680 195763 49736
rect 194428 49678 195763 49680
rect 196296 49736 196388 49738
rect 196296 49680 196346 49736
rect 196296 49678 196388 49680
rect 194428 49676 194434 49678
rect 183921 49675 183987 49676
rect 195697 49675 195763 49678
rect 196341 49676 196388 49678
rect 196452 49676 196458 49740
rect 202045 49738 202092 49740
rect 202000 49736 202092 49738
rect 202000 49680 202050 49736
rect 202000 49678 202092 49680
rect 202045 49676 202092 49678
rect 202156 49676 202162 49740
rect 206870 49676 206876 49740
rect 206940 49738 206946 49740
rect 209589 49738 209655 49741
rect 206940 49736 209655 49738
rect 206940 49680 209594 49736
rect 209650 49680 209655 49736
rect 206940 49678 209655 49680
rect 206940 49676 206946 49678
rect 196341 49675 196407 49676
rect 202045 49675 202111 49676
rect 209589 49675 209655 49678
rect 209865 49738 209931 49741
rect 210734 49738 210740 49740
rect 209865 49736 210740 49738
rect 209865 49680 209870 49736
rect 209926 49680 210740 49736
rect 209865 49678 210740 49680
rect 209865 49675 209931 49678
rect 210734 49676 210740 49678
rect 210804 49676 210810 49740
rect 213678 49676 213684 49740
rect 213748 49738 213754 49740
rect 214189 49738 214255 49741
rect 213748 49736 214255 49738
rect 213748 49680 214194 49736
rect 214250 49680 214255 49736
rect 213748 49678 214255 49680
rect 213748 49676 213754 49678
rect 214189 49675 214255 49678
rect 157885 49602 157951 49605
rect 176326 49602 176332 49604
rect 157885 49600 176332 49602
rect 157885 49544 157890 49600
rect 157946 49544 176332 49600
rect 157885 49542 176332 49544
rect 157885 49539 157951 49542
rect 176326 49540 176332 49542
rect 176396 49540 176402 49604
rect 177021 49602 177087 49605
rect 229921 49602 229987 49605
rect 177021 49600 229987 49602
rect 177021 49544 177026 49600
rect 177082 49544 229926 49600
rect 229982 49544 229987 49600
rect 177021 49542 229987 49544
rect 177021 49539 177087 49542
rect 229921 49539 229987 49542
rect 165705 49468 165771 49469
rect 165654 49466 165660 49468
rect 165614 49406 165660 49466
rect 165724 49464 165771 49468
rect 165766 49408 165771 49464
rect 165654 49404 165660 49406
rect 165724 49404 165771 49408
rect 165705 49403 165771 49404
rect 165889 49466 165955 49469
rect 166206 49466 166212 49468
rect 165889 49464 166212 49466
rect 165889 49408 165894 49464
rect 165950 49408 166212 49464
rect 165889 49406 166212 49408
rect 165889 49403 165955 49406
rect 166206 49404 166212 49406
rect 166276 49404 166282 49468
rect 172421 49466 172487 49469
rect 221641 49466 221707 49469
rect 172421 49464 221707 49466
rect 172421 49408 172426 49464
rect 172482 49408 221646 49464
rect 221702 49408 221707 49464
rect 172421 49406 221707 49408
rect 172421 49403 172487 49406
rect 221641 49403 221707 49406
rect 256693 49466 256759 49469
rect 256693 49464 260084 49466
rect 256693 49408 256698 49464
rect 256754 49408 260084 49464
rect 256693 49406 260084 49408
rect 256693 49403 256759 49406
rect 140037 49330 140103 49333
rect 177297 49330 177363 49333
rect 140037 49328 177363 49330
rect 140037 49272 140042 49328
rect 140098 49272 177302 49328
rect 177358 49272 177363 49328
rect 140037 49270 177363 49272
rect 140037 49267 140103 49270
rect 177297 49267 177363 49270
rect 177849 49330 177915 49333
rect 226977 49330 227043 49333
rect 177849 49328 227043 49330
rect 177849 49272 177854 49328
rect 177910 49272 226982 49328
rect 227038 49272 227043 49328
rect 177849 49270 227043 49272
rect 177849 49267 177915 49270
rect 226977 49267 227043 49270
rect 152549 49194 152615 49197
rect 177665 49194 177731 49197
rect 152549 49192 177731 49194
rect 152549 49136 152554 49192
rect 152610 49136 177670 49192
rect 177726 49136 177731 49192
rect 152549 49134 177731 49136
rect 152549 49131 152615 49134
rect 177665 49131 177731 49134
rect 177941 49194 178007 49197
rect 219157 49194 219223 49197
rect 177941 49192 219223 49194
rect 177941 49136 177946 49192
rect 178002 49136 219162 49192
rect 219218 49136 219223 49192
rect 177941 49134 219223 49136
rect 177941 49131 178007 49134
rect 219157 49131 219223 49134
rect 158253 49058 158319 49061
rect 177113 49058 177179 49061
rect 158253 49056 177179 49058
rect 158253 49000 158258 49056
rect 158314 49000 177118 49056
rect 177174 49000 177179 49056
rect 158253 48998 177179 49000
rect 158253 48995 158319 48998
rect 177113 48995 177179 48998
rect 182357 49058 182423 49061
rect 182950 49058 182956 49060
rect 182357 49056 182956 49058
rect 182357 49000 182362 49056
rect 182418 49000 182956 49056
rect 182357 48998 182956 49000
rect 182357 48995 182423 48998
rect 182950 48996 182956 48998
rect 183020 48996 183026 49060
rect 187141 49058 187207 49061
rect 209773 49058 209839 49061
rect 215150 49058 215156 49060
rect 187141 49056 205650 49058
rect 187141 49000 187146 49056
rect 187202 49000 205650 49056
rect 187141 48998 205650 49000
rect 187141 48995 187207 48998
rect 153929 48922 153995 48925
rect 161381 48922 161447 48925
rect 153929 48920 161447 48922
rect 153929 48864 153934 48920
rect 153990 48864 161386 48920
rect 161442 48864 161447 48920
rect 153929 48862 161447 48864
rect 153929 48859 153995 48862
rect 161381 48859 161447 48862
rect 161749 48922 161815 48925
rect 161974 48922 161980 48924
rect 161749 48920 161980 48922
rect 161749 48864 161754 48920
rect 161810 48864 161980 48920
rect 161749 48862 161980 48864
rect 161749 48859 161815 48862
rect 161974 48860 161980 48862
rect 162044 48860 162050 48924
rect 162945 48922 163011 48925
rect 163262 48922 163268 48924
rect 162945 48920 163268 48922
rect 162945 48864 162950 48920
rect 163006 48864 163268 48920
rect 162945 48862 163268 48864
rect 162945 48859 163011 48862
rect 163262 48860 163268 48862
rect 163332 48860 163338 48924
rect 170070 48860 170076 48924
rect 170140 48922 170146 48924
rect 172145 48922 172211 48925
rect 170140 48920 172211 48922
rect 170140 48864 172150 48920
rect 172206 48864 172211 48920
rect 170140 48862 172211 48864
rect 170140 48860 170146 48862
rect 172145 48859 172211 48862
rect 177941 48922 178007 48925
rect 198457 48924 198523 48925
rect 177941 48920 195990 48922
rect 177941 48864 177946 48920
rect 178002 48864 195990 48920
rect 177941 48862 195990 48864
rect 177941 48859 178007 48862
rect 163129 48788 163195 48789
rect 163078 48724 163084 48788
rect 163148 48786 163195 48788
rect 163313 48786 163379 48789
rect 163446 48786 163452 48788
rect 163148 48784 163240 48786
rect 163190 48728 163240 48784
rect 163148 48726 163240 48728
rect 163313 48784 163452 48786
rect 163313 48728 163318 48784
rect 163374 48728 163452 48784
rect 163313 48726 163452 48728
rect 163148 48724 163195 48726
rect 163129 48723 163195 48724
rect 163313 48723 163379 48726
rect 163446 48724 163452 48726
rect 163516 48724 163522 48788
rect 170305 48786 170371 48789
rect 170990 48786 170996 48788
rect 170305 48784 170996 48786
rect 170305 48728 170310 48784
rect 170366 48728 170996 48784
rect 170305 48726 170996 48728
rect 170305 48723 170371 48726
rect 170990 48724 170996 48726
rect 171060 48724 171066 48788
rect 182265 48786 182331 48789
rect 184473 48788 184539 48789
rect 183134 48786 183140 48788
rect 182265 48784 183140 48786
rect 182265 48728 182270 48784
rect 182326 48728 183140 48784
rect 182265 48726 183140 48728
rect 182265 48723 182331 48726
rect 183134 48724 183140 48726
rect 183204 48724 183210 48788
rect 184422 48724 184428 48788
rect 184492 48786 184539 48788
rect 184492 48784 184584 48786
rect 184534 48728 184584 48784
rect 184492 48726 184584 48728
rect 184492 48724 184539 48726
rect 186998 48724 187004 48788
rect 187068 48786 187074 48788
rect 187601 48786 187667 48789
rect 187068 48784 187667 48786
rect 187068 48728 187606 48784
rect 187662 48728 187667 48784
rect 187068 48726 187667 48728
rect 187068 48724 187074 48726
rect 184473 48723 184539 48724
rect 187601 48723 187667 48726
rect 192150 48724 192156 48788
rect 192220 48786 192226 48788
rect 192937 48786 193003 48789
rect 192220 48784 193003 48786
rect 192220 48728 192942 48784
rect 192998 48728 193003 48784
rect 192220 48726 193003 48728
rect 195930 48786 195990 48862
rect 198406 48860 198412 48924
rect 198476 48922 198523 48924
rect 198476 48920 198568 48922
rect 198518 48864 198568 48920
rect 198476 48862 198568 48864
rect 198476 48860 198523 48862
rect 202086 48860 202092 48924
rect 202156 48922 202162 48924
rect 202505 48922 202571 48925
rect 202156 48920 202571 48922
rect 202156 48864 202510 48920
rect 202566 48864 202571 48920
rect 202156 48862 202571 48864
rect 202156 48860 202162 48862
rect 198457 48859 198523 48860
rect 202505 48859 202571 48862
rect 203190 48860 203196 48924
rect 203260 48922 203266 48924
rect 203977 48922 204043 48925
rect 203260 48920 204043 48922
rect 203260 48864 203982 48920
rect 204038 48864 204043 48920
rect 203260 48862 204043 48864
rect 205590 48922 205650 48998
rect 209773 49056 210250 49058
rect 209773 49000 209778 49056
rect 209834 49000 210250 49056
rect 209773 48998 210250 49000
rect 209773 48995 209839 48998
rect 209129 48922 209195 48925
rect 210049 48922 210115 48925
rect 205590 48920 209195 48922
rect 205590 48864 209134 48920
rect 209190 48864 209195 48920
rect 205590 48862 209195 48864
rect 203260 48860 203266 48862
rect 203977 48859 204043 48862
rect 209129 48859 209195 48862
rect 209776 48920 210115 48922
rect 209776 48864 210054 48920
rect 210110 48864 210115 48920
rect 209776 48862 210115 48864
rect 210190 48922 210250 48998
rect 211110 48998 215156 49058
rect 211110 48922 211170 48998
rect 215150 48996 215156 48998
rect 215220 48996 215226 49060
rect 210190 48862 211170 48922
rect 209776 48789 209836 48862
rect 210049 48859 210115 48862
rect 213126 48860 213132 48924
rect 213196 48922 213202 48924
rect 213821 48922 213887 48925
rect 213196 48920 213887 48922
rect 213196 48864 213826 48920
rect 213882 48864 213887 48920
rect 213196 48862 213887 48864
rect 213196 48860 213202 48862
rect 213821 48859 213887 48862
rect 214414 48860 214420 48924
rect 214484 48922 214490 48924
rect 215017 48922 215083 48925
rect 214484 48920 215083 48922
rect 214484 48864 215022 48920
rect 215078 48864 215083 48920
rect 214484 48862 215083 48864
rect 214484 48860 214490 48862
rect 215017 48859 215083 48862
rect 195930 48726 205650 48786
rect 192220 48724 192226 48726
rect 192937 48723 193003 48726
rect 164417 48650 164483 48653
rect 165286 48650 165292 48652
rect 164417 48648 165292 48650
rect 164417 48592 164422 48648
rect 164478 48592 165292 48648
rect 164417 48590 165292 48592
rect 164417 48587 164483 48590
rect 165286 48588 165292 48590
rect 165356 48588 165362 48652
rect 170305 48650 170371 48653
rect 170438 48650 170444 48652
rect 170305 48648 170444 48650
rect 170305 48592 170310 48648
rect 170366 48592 170444 48648
rect 170305 48590 170444 48592
rect 170305 48587 170371 48590
rect 170438 48588 170444 48590
rect 170508 48588 170514 48652
rect 176929 48650 176995 48653
rect 176929 48648 186330 48650
rect 176929 48592 176934 48648
rect 176990 48592 186330 48648
rect 176929 48590 186330 48592
rect 176929 48587 176995 48590
rect 142889 48514 142955 48517
rect 177573 48514 177639 48517
rect 142889 48512 177639 48514
rect 142889 48456 142894 48512
rect 142950 48456 177578 48512
rect 177634 48456 177639 48512
rect 142889 48454 177639 48456
rect 142889 48451 142955 48454
rect 177573 48451 177639 48454
rect 180885 48514 180951 48517
rect 182541 48516 182607 48517
rect 184565 48516 184631 48517
rect 181294 48514 181300 48516
rect 180885 48512 181300 48514
rect 180885 48456 180890 48512
rect 180946 48456 181300 48512
rect 180885 48454 181300 48456
rect 180885 48451 180951 48454
rect 181294 48452 181300 48454
rect 181364 48452 181370 48516
rect 182541 48512 182588 48516
rect 182652 48514 182658 48516
rect 184565 48514 184612 48516
rect 182541 48456 182546 48512
rect 182541 48452 182588 48456
rect 182652 48454 182698 48514
rect 184520 48512 184612 48514
rect 184520 48456 184570 48512
rect 184520 48454 184612 48456
rect 182652 48452 182658 48454
rect 184565 48452 184612 48454
rect 184676 48452 184682 48516
rect 185158 48514 185164 48516
rect 184798 48454 185164 48514
rect 182541 48451 182607 48452
rect 184565 48451 184631 48452
rect 184798 48381 184858 48454
rect 185158 48452 185164 48454
rect 185228 48452 185234 48516
rect 185342 48452 185348 48516
rect 185412 48514 185418 48516
rect 186037 48514 186103 48517
rect 185412 48512 186103 48514
rect 185412 48456 186042 48512
rect 186098 48456 186103 48512
rect 185412 48454 186103 48456
rect 185412 48452 185418 48454
rect 186037 48451 186103 48454
rect 134609 48378 134675 48381
rect 178309 48378 178375 48381
rect 134609 48376 178375 48378
rect 134609 48320 134614 48376
rect 134670 48320 178314 48376
rect 178370 48320 178375 48376
rect 134609 48318 178375 48320
rect 134609 48315 134675 48318
rect 178309 48315 178375 48318
rect 181110 48316 181116 48380
rect 181180 48378 181186 48380
rect 181253 48378 181319 48381
rect 181180 48376 181319 48378
rect 181180 48320 181258 48376
rect 181314 48320 181319 48376
rect 181180 48318 181319 48320
rect 181180 48316 181186 48318
rect 181253 48315 181319 48318
rect 184749 48376 184858 48381
rect 184749 48320 184754 48376
rect 184810 48320 184858 48376
rect 184749 48318 184858 48320
rect 184749 48315 184815 48318
rect 185158 48316 185164 48380
rect 185228 48378 185234 48380
rect 186129 48378 186195 48381
rect 185228 48376 186195 48378
rect 185228 48320 186134 48376
rect 186190 48320 186195 48376
rect 185228 48318 186195 48320
rect 186270 48378 186330 48590
rect 187182 48588 187188 48652
rect 187252 48650 187258 48652
rect 187509 48650 187575 48653
rect 187252 48648 187575 48650
rect 187252 48592 187514 48648
rect 187570 48592 187575 48648
rect 187252 48590 187575 48592
rect 187252 48588 187258 48590
rect 187509 48587 187575 48590
rect 188889 48650 188955 48653
rect 189022 48650 189028 48652
rect 188889 48648 189028 48650
rect 188889 48592 188894 48648
rect 188950 48592 189028 48648
rect 188889 48590 189028 48592
rect 188889 48587 188955 48590
rect 189022 48588 189028 48590
rect 189092 48588 189098 48652
rect 192334 48588 192340 48652
rect 192404 48650 192410 48652
rect 193121 48650 193187 48653
rect 192404 48648 193187 48650
rect 192404 48592 193126 48648
rect 193182 48592 193187 48648
rect 192404 48590 193187 48592
rect 192404 48588 192410 48590
rect 193121 48587 193187 48590
rect 196198 48588 196204 48652
rect 196268 48650 196274 48652
rect 197261 48650 197327 48653
rect 196268 48648 197327 48650
rect 196268 48592 197266 48648
rect 197322 48592 197327 48648
rect 196268 48590 197327 48592
rect 196268 48588 196274 48590
rect 197261 48587 197327 48590
rect 198038 48588 198044 48652
rect 198108 48650 198114 48652
rect 198549 48650 198615 48653
rect 198108 48648 198615 48650
rect 198108 48592 198554 48648
rect 198610 48592 198615 48648
rect 198108 48590 198615 48592
rect 198108 48588 198114 48590
rect 198549 48587 198615 48590
rect 199326 48588 199332 48652
rect 199396 48650 199402 48652
rect 199837 48650 199903 48653
rect 199396 48648 199903 48650
rect 199396 48592 199842 48648
rect 199898 48592 199903 48648
rect 199396 48590 199903 48592
rect 199396 48588 199402 48590
rect 199837 48587 199903 48590
rect 202270 48588 202276 48652
rect 202340 48650 202346 48652
rect 202597 48650 202663 48653
rect 202340 48648 202663 48650
rect 202340 48592 202602 48648
rect 202658 48592 202663 48648
rect 202340 48590 202663 48592
rect 202340 48588 202346 48590
rect 202597 48587 202663 48590
rect 187233 48514 187299 48517
rect 187550 48514 187556 48516
rect 187233 48512 187556 48514
rect 187233 48456 187238 48512
rect 187294 48456 187556 48512
rect 187233 48454 187556 48456
rect 187233 48451 187299 48454
rect 187550 48452 187556 48454
rect 187620 48452 187626 48516
rect 192518 48452 192524 48516
rect 192588 48514 192594 48516
rect 193029 48514 193095 48517
rect 192588 48512 193095 48514
rect 192588 48456 193034 48512
rect 193090 48456 193095 48512
rect 192588 48454 193095 48456
rect 192588 48452 192594 48454
rect 193029 48451 193095 48454
rect 199694 48452 199700 48516
rect 199764 48514 199770 48516
rect 199929 48514 199995 48517
rect 199764 48512 199995 48514
rect 199764 48456 199934 48512
rect 199990 48456 199995 48512
rect 199764 48454 199995 48456
rect 199764 48452 199770 48454
rect 199929 48451 199995 48454
rect 202454 48452 202460 48516
rect 202524 48514 202530 48516
rect 202781 48514 202847 48517
rect 202524 48512 202847 48514
rect 202524 48456 202786 48512
rect 202842 48456 202847 48512
rect 202524 48454 202847 48456
rect 205590 48514 205650 48726
rect 209773 48784 209839 48789
rect 209773 48728 209778 48784
rect 209834 48728 209839 48784
rect 209773 48723 209839 48728
rect 210182 48724 210188 48788
rect 210252 48786 210258 48788
rect 210325 48786 210391 48789
rect 210785 48788 210851 48789
rect 210734 48786 210740 48788
rect 210252 48784 210391 48786
rect 210252 48728 210330 48784
rect 210386 48728 210391 48784
rect 210252 48726 210391 48728
rect 210694 48726 210740 48786
rect 210804 48784 210851 48788
rect 210846 48728 210851 48784
rect 210252 48724 210258 48726
rect 210325 48723 210391 48726
rect 210734 48724 210740 48726
rect 210804 48724 210851 48728
rect 211838 48724 211844 48788
rect 211908 48786 211914 48788
rect 212257 48786 212323 48789
rect 211908 48784 212323 48786
rect 211908 48728 212262 48784
rect 212318 48728 212323 48784
rect 211908 48726 212323 48728
rect 211908 48724 211914 48726
rect 210785 48723 210851 48724
rect 212257 48723 212323 48726
rect 214782 48724 214788 48788
rect 214852 48786 214858 48788
rect 215201 48786 215267 48789
rect 214852 48784 215267 48786
rect 214852 48728 215206 48784
rect 215262 48728 215267 48784
rect 214852 48726 215267 48728
rect 214852 48724 214858 48726
rect 215201 48723 215267 48726
rect 215518 48724 215524 48788
rect 215588 48786 215594 48788
rect 215753 48786 215819 48789
rect 229737 48786 229803 48789
rect 215588 48784 215819 48786
rect 215588 48728 215758 48784
rect 215814 48728 215819 48784
rect 215588 48726 215819 48728
rect 215588 48724 215594 48726
rect 215753 48723 215819 48726
rect 224910 48784 229803 48786
rect 224910 48728 229742 48784
rect 229798 48728 229803 48784
rect 224910 48726 229803 48728
rect 208301 48650 208367 48653
rect 224910 48650 224970 48726
rect 229737 48723 229803 48726
rect 208301 48648 224970 48650
rect 208301 48592 208306 48648
rect 208362 48592 224970 48648
rect 208301 48590 224970 48592
rect 208301 48587 208367 48590
rect 218789 48514 218855 48517
rect 205590 48512 218855 48514
rect 205590 48456 218794 48512
rect 218850 48456 218855 48512
rect 205590 48454 218855 48456
rect 202524 48452 202530 48454
rect 202781 48451 202847 48454
rect 218789 48451 218855 48454
rect 187141 48378 187207 48381
rect 187417 48380 187483 48381
rect 187366 48378 187372 48380
rect 186270 48376 187207 48378
rect 186270 48320 187146 48376
rect 187202 48320 187207 48376
rect 186270 48318 187207 48320
rect 187326 48318 187372 48378
rect 187436 48376 187483 48380
rect 187478 48320 187483 48376
rect 185228 48316 185234 48318
rect 186129 48315 186195 48318
rect 187141 48315 187207 48318
rect 187366 48316 187372 48318
rect 187436 48316 187483 48320
rect 188654 48316 188660 48380
rect 188724 48378 188730 48380
rect 188981 48378 189047 48381
rect 188724 48376 189047 48378
rect 188724 48320 188986 48376
rect 189042 48320 189047 48376
rect 188724 48318 189047 48320
rect 188724 48316 188730 48318
rect 187417 48315 187483 48316
rect 188981 48315 189047 48318
rect 189717 48378 189783 48381
rect 190310 48378 190316 48380
rect 189717 48376 190316 48378
rect 189717 48320 189722 48376
rect 189778 48320 190316 48376
rect 189717 48318 190316 48320
rect 189717 48315 189783 48318
rect 190310 48316 190316 48318
rect 190380 48316 190386 48380
rect 199009 48378 199075 48381
rect 199510 48378 199516 48380
rect 199009 48376 199516 48378
rect 199009 48320 199014 48376
rect 199070 48320 199516 48376
rect 199009 48318 199516 48320
rect 199009 48315 199075 48318
rect 199510 48316 199516 48318
rect 199580 48316 199586 48380
rect 199745 48378 199811 48381
rect 201401 48380 201467 48381
rect 202689 48380 202755 48381
rect 203793 48380 203859 48381
rect 199878 48378 199884 48380
rect 199745 48376 199884 48378
rect 199745 48320 199750 48376
rect 199806 48320 199884 48376
rect 199745 48318 199884 48320
rect 199745 48315 199811 48318
rect 199878 48316 199884 48318
rect 199948 48316 199954 48380
rect 201350 48378 201356 48380
rect 201310 48318 201356 48378
rect 201420 48376 201467 48380
rect 202638 48378 202644 48380
rect 201462 48320 201467 48376
rect 201350 48316 201356 48318
rect 201420 48316 201467 48320
rect 202598 48318 202644 48378
rect 202708 48376 202755 48380
rect 203742 48378 203748 48380
rect 202750 48320 202755 48376
rect 202638 48316 202644 48318
rect 202708 48316 202755 48320
rect 203702 48318 203748 48378
rect 203812 48376 203859 48380
rect 203854 48320 203859 48376
rect 203742 48316 203748 48318
rect 203812 48316 203859 48320
rect 205030 48316 205036 48380
rect 205100 48378 205106 48380
rect 205357 48378 205423 48381
rect 205100 48376 205423 48378
rect 205100 48320 205362 48376
rect 205418 48320 205423 48376
rect 205100 48318 205423 48320
rect 205100 48316 205106 48318
rect 201401 48315 201467 48316
rect 202689 48315 202755 48316
rect 203793 48315 203859 48316
rect 205357 48315 205423 48318
rect 206134 48316 206140 48380
rect 206204 48378 206210 48380
rect 206461 48378 206527 48381
rect 214189 48380 214255 48381
rect 214189 48378 214236 48380
rect 206204 48376 206527 48378
rect 206204 48320 206466 48376
rect 206522 48320 206527 48376
rect 206204 48318 206527 48320
rect 214144 48376 214236 48378
rect 214144 48320 214194 48376
rect 214144 48318 214236 48320
rect 206204 48316 206210 48318
rect 206461 48315 206527 48318
rect 214189 48316 214236 48318
rect 214300 48316 214306 48380
rect 214598 48316 214604 48380
rect 214668 48378 214674 48380
rect 214833 48378 214899 48381
rect 214668 48376 214899 48378
rect 214668 48320 214838 48376
rect 214894 48320 214899 48376
rect 214668 48318 214899 48320
rect 214668 48316 214674 48318
rect 214189 48315 214255 48316
rect 214833 48315 214899 48318
rect 215150 48316 215156 48380
rect 215220 48378 215226 48380
rect 218973 48378 219039 48381
rect 215220 48376 219039 48378
rect 215220 48320 218978 48376
rect 219034 48320 219039 48376
rect 215220 48318 219039 48320
rect 215220 48316 215226 48318
rect 218973 48315 219039 48318
rect 173985 48242 174051 48245
rect 246297 48242 246363 48245
rect 173985 48240 246363 48242
rect 173985 48184 173990 48240
rect 174046 48184 246302 48240
rect 246358 48184 246363 48240
rect 173985 48182 246363 48184
rect 173985 48179 174051 48182
rect 246297 48179 246363 48182
rect 168557 48106 168623 48109
rect 169334 48106 169340 48108
rect 168557 48104 169340 48106
rect 168557 48048 168562 48104
rect 168618 48048 169340 48104
rect 168557 48046 169340 48048
rect 168557 48043 168623 48046
rect 169334 48044 169340 48046
rect 169404 48044 169410 48108
rect 174261 48106 174327 48109
rect 243537 48106 243603 48109
rect 174261 48104 243603 48106
rect 174261 48048 174266 48104
rect 174322 48048 243542 48104
rect 243598 48048 243603 48104
rect 174261 48046 243603 48048
rect 174261 48043 174327 48046
rect 243537 48043 243603 48046
rect 133830 47698 133890 48008
rect 179965 47972 180031 47973
rect 180149 47972 180215 47973
rect 179965 47970 180012 47972
rect 179920 47968 180012 47970
rect 179920 47912 179970 47968
rect 179920 47910 180012 47912
rect 179965 47908 180012 47910
rect 180076 47908 180082 47972
rect 180149 47968 180196 47972
rect 180260 47970 180266 47972
rect 180425 47970 180491 47973
rect 180558 47970 180564 47972
rect 180149 47912 180154 47968
rect 180149 47908 180196 47912
rect 180260 47910 180306 47970
rect 180425 47968 180564 47970
rect 180425 47912 180430 47968
rect 180486 47912 180564 47968
rect 180425 47910 180564 47912
rect 180260 47908 180266 47910
rect 179965 47907 180031 47908
rect 180149 47907 180215 47908
rect 180425 47907 180491 47910
rect 180558 47908 180564 47910
rect 180628 47908 180634 47972
rect 181161 47970 181227 47973
rect 181294 47970 181300 47972
rect 181161 47968 181300 47970
rect 181161 47912 181166 47968
rect 181222 47912 181300 47968
rect 181161 47910 181300 47912
rect 181161 47907 181227 47910
rect 181294 47908 181300 47910
rect 181364 47908 181370 47972
rect 214046 47908 214052 47972
rect 214116 47970 214122 47972
rect 214557 47970 214623 47973
rect 214116 47968 214623 47970
rect 214116 47912 214562 47968
rect 214618 47912 214623 47968
rect 214116 47910 214623 47912
rect 214116 47908 214122 47910
rect 214557 47907 214623 47910
rect 214966 47908 214972 47972
rect 215036 47970 215042 47972
rect 215109 47970 215175 47973
rect 215036 47968 215175 47970
rect 215036 47912 215114 47968
rect 215170 47912 215175 47968
rect 215036 47910 215175 47912
rect 215036 47908 215042 47910
rect 215109 47907 215175 47910
rect 136541 47698 136607 47701
rect 133830 47696 136607 47698
rect 133830 47640 136546 47696
rect 136602 47640 136607 47696
rect 133830 47638 136607 47640
rect 136541 47635 136607 47638
rect 167269 47698 167335 47701
rect 167678 47698 167684 47700
rect 167269 47696 167684 47698
rect 167269 47640 167274 47696
rect 167330 47640 167684 47696
rect 167269 47638 167684 47640
rect 167269 47635 167335 47638
rect 167678 47636 167684 47638
rect 167748 47636 167754 47700
rect 195646 47636 195652 47700
rect 195716 47698 195722 47700
rect 195881 47698 195947 47701
rect 195716 47696 195947 47698
rect 195716 47640 195886 47696
rect 195942 47640 195947 47696
rect 195716 47638 195947 47640
rect 195716 47636 195722 47638
rect 195881 47635 195947 47638
rect 133321 47562 133387 47565
rect 167361 47564 167427 47565
rect 163814 47562 163820 47564
rect 133321 47560 163820 47562
rect 133321 47504 133326 47560
rect 133382 47504 163820 47560
rect 133321 47502 163820 47504
rect 133321 47499 133387 47502
rect 163814 47500 163820 47502
rect 163884 47500 163890 47564
rect 167310 47562 167316 47564
rect 167270 47502 167316 47562
rect 167380 47560 167427 47564
rect 167422 47504 167427 47560
rect 167310 47500 167316 47502
rect 167380 47500 167427 47504
rect 167361 47499 167427 47500
rect 173157 47562 173223 47565
rect 182173 47562 182239 47565
rect 194409 47564 194475 47565
rect 194358 47562 194364 47564
rect 173157 47560 182239 47562
rect 173157 47504 173162 47560
rect 173218 47504 182178 47560
rect 182234 47504 182239 47560
rect 173157 47502 182239 47504
rect 194318 47502 194364 47562
rect 194428 47560 194475 47564
rect 194470 47504 194475 47560
rect 173157 47499 173223 47502
rect 182173 47499 182239 47502
rect 194358 47500 194364 47502
rect 194428 47500 194475 47504
rect 194409 47499 194475 47500
rect 194685 47562 194751 47565
rect 195094 47562 195100 47564
rect 194685 47560 195100 47562
rect 194685 47504 194690 47560
rect 194746 47504 195100 47560
rect 194685 47502 195100 47504
rect 194685 47499 194751 47502
rect 195094 47500 195100 47502
rect 195164 47500 195170 47564
rect 195605 47562 195671 47565
rect 195830 47562 195836 47564
rect 195605 47560 195836 47562
rect 195605 47504 195610 47560
rect 195666 47504 195836 47560
rect 195605 47502 195836 47504
rect 195605 47499 195671 47502
rect 195830 47500 195836 47502
rect 195900 47500 195906 47564
rect 207606 47500 207612 47564
rect 207676 47562 207682 47564
rect 217317 47562 217383 47565
rect 207676 47560 217383 47562
rect 207676 47504 217322 47560
rect 217378 47504 217383 47560
rect 207676 47502 217383 47504
rect 207676 47500 207682 47502
rect 217317 47499 217383 47502
rect 166717 47428 166783 47429
rect 167085 47428 167151 47429
rect 166717 47426 166764 47428
rect 166672 47424 166764 47426
rect 166672 47368 166722 47424
rect 166672 47366 166764 47368
rect 166717 47364 166764 47366
rect 166828 47364 166834 47428
rect 167085 47424 167132 47428
rect 167196 47426 167202 47428
rect 193581 47426 193647 47429
rect 193806 47426 193812 47428
rect 167085 47368 167090 47424
rect 167085 47364 167132 47368
rect 167196 47366 167242 47426
rect 193581 47424 193812 47426
rect 193581 47368 193586 47424
rect 193642 47368 193812 47424
rect 193581 47366 193812 47368
rect 167196 47364 167202 47366
rect 166717 47363 166783 47364
rect 167085 47363 167151 47364
rect 193581 47363 193647 47366
rect 193806 47364 193812 47366
rect 193876 47364 193882 47428
rect 194174 47364 194180 47428
rect 194244 47426 194250 47428
rect 194317 47426 194383 47429
rect 194244 47424 194383 47426
rect 194244 47368 194322 47424
rect 194378 47368 194383 47424
rect 194244 47366 194383 47368
rect 194244 47364 194250 47366
rect 194317 47363 194383 47366
rect 194726 47364 194732 47428
rect 194796 47426 194802 47428
rect 194869 47426 194935 47429
rect 194796 47424 194935 47426
rect 194796 47368 194874 47424
rect 194930 47368 194935 47424
rect 194796 47366 194935 47368
rect 194796 47364 194802 47366
rect 194869 47363 194935 47366
rect 195278 47364 195284 47428
rect 195348 47426 195354 47428
rect 195789 47426 195855 47429
rect 195348 47424 195855 47426
rect 195348 47368 195794 47424
rect 195850 47368 195855 47424
rect 195348 47366 195855 47368
rect 195348 47364 195354 47366
rect 195789 47363 195855 47366
rect 194910 47228 194916 47292
rect 194980 47290 194986 47292
rect 195605 47290 195671 47293
rect 194980 47288 195671 47290
rect 194980 47232 195610 47288
rect 195666 47232 195671 47288
rect 194980 47230 195671 47232
rect 194980 47228 194986 47230
rect 195605 47227 195671 47230
rect 163405 46882 163471 46885
rect 163630 46882 163636 46884
rect 163405 46880 163636 46882
rect 163405 46824 163410 46880
rect 163466 46824 163636 46880
rect 163405 46822 163636 46824
rect 163405 46819 163471 46822
rect 163630 46820 163636 46822
rect 163700 46820 163706 46884
rect 201953 46746 202019 46749
rect 201910 46744 202019 46746
rect 201910 46688 201958 46744
rect 202014 46688 202019 46744
rect 201910 46683 202019 46688
rect 201910 46477 201970 46683
rect 201861 46472 201970 46477
rect 201861 46416 201866 46472
rect 201922 46416 201970 46472
rect 201861 46414 201970 46416
rect 201861 46411 201927 46414
rect 137277 46338 137343 46341
rect 162158 46338 162164 46340
rect 137277 46336 162164 46338
rect 137277 46280 137282 46336
rect 137338 46280 162164 46336
rect 137277 46278 162164 46280
rect 137277 46275 137343 46278
rect 162158 46276 162164 46278
rect 162228 46276 162234 46340
rect 189022 46276 189028 46340
rect 189092 46338 189098 46340
rect 231853 46338 231919 46341
rect 189092 46336 231919 46338
rect 189092 46280 231858 46336
rect 231914 46280 231919 46336
rect 189092 46278 231919 46280
rect 189092 46276 189098 46278
rect 231853 46275 231919 46278
rect 580809 46338 580875 46341
rect 583520 46338 584960 46428
rect 580809 46336 584960 46338
rect 580809 46280 580814 46336
rect 580870 46280 584960 46336
rect 580809 46278 584960 46280
rect 580809 46275 580875 46278
rect 134793 46202 134859 46205
rect 167177 46202 167243 46205
rect 134793 46200 167243 46202
rect 134793 46144 134798 46200
rect 134854 46144 167182 46200
rect 167238 46144 167243 46200
rect 134793 46142 167243 46144
rect 134793 46139 134859 46142
rect 167177 46139 167243 46142
rect 174537 46202 174603 46205
rect 183645 46202 183711 46205
rect 174537 46200 183711 46202
rect 174537 46144 174542 46200
rect 174598 46144 183650 46200
rect 183706 46144 183711 46200
rect 174537 46142 183711 46144
rect 174537 46139 174603 46142
rect 183645 46139 183711 46142
rect 201493 46202 201559 46205
rect 201861 46202 201927 46205
rect 201493 46200 201927 46202
rect 201493 46144 201498 46200
rect 201554 46144 201866 46200
rect 201922 46144 201927 46200
rect 201493 46142 201927 46144
rect 201493 46139 201559 46142
rect 201861 46139 201927 46142
rect 206870 46140 206876 46204
rect 206940 46202 206946 46204
rect 260097 46202 260163 46205
rect 206940 46200 260163 46202
rect 206940 46144 260102 46200
rect 260158 46144 260163 46200
rect 583520 46188 584960 46278
rect 206940 46142 260163 46144
rect 206940 46140 206946 46142
rect 260097 46139 260163 46142
rect 160737 46066 160803 46069
rect 161422 46066 161428 46068
rect 160737 46064 161428 46066
rect 160737 46008 160742 46064
rect 160798 46008 161428 46064
rect 160737 46006 161428 46008
rect 160737 46003 160803 46006
rect 161422 46004 161428 46006
rect 161492 46004 161498 46068
rect 162025 45930 162091 45933
rect 162710 45930 162716 45932
rect 162025 45928 162716 45930
rect 162025 45872 162030 45928
rect 162086 45872 162716 45928
rect 162025 45870 162716 45872
rect 162025 45867 162091 45870
rect 162710 45868 162716 45870
rect 162780 45868 162786 45932
rect 167494 45732 167500 45796
rect 167564 45794 167570 45796
rect 167821 45794 167887 45797
rect 167564 45792 167887 45794
rect 167564 45736 167826 45792
rect 167882 45736 167887 45792
rect 167564 45734 167887 45736
rect 167564 45732 167570 45734
rect 167821 45731 167887 45734
rect 211245 45794 211311 45797
rect 211654 45794 211660 45796
rect 211245 45792 211660 45794
rect 211245 45736 211250 45792
rect 211306 45736 211660 45792
rect 211245 45734 211660 45736
rect 211245 45731 211311 45734
rect 211654 45732 211660 45734
rect 211724 45732 211730 45796
rect -960 45522 480 45612
rect 3693 45522 3759 45525
rect 135621 45522 135687 45525
rect -960 45520 3759 45522
rect -960 45464 3698 45520
rect 3754 45464 3759 45520
rect -960 45462 3759 45464
rect -960 45372 480 45462
rect 3693 45459 3759 45462
rect 133830 45520 135687 45522
rect 133830 45464 135626 45520
rect 135682 45464 135687 45520
rect 133830 45462 135687 45464
rect 133830 45424 133890 45462
rect 135621 45459 135687 45462
rect 186998 45460 187004 45524
rect 187068 45522 187074 45524
rect 189809 45522 189875 45525
rect 187068 45520 189875 45522
rect 187068 45464 189814 45520
rect 189870 45464 189875 45520
rect 187068 45462 189875 45464
rect 187068 45460 187074 45462
rect 189809 45459 189875 45462
rect 146293 44978 146359 44981
rect 182950 44978 182956 44980
rect 146293 44976 182956 44978
rect 146293 44920 146298 44976
rect 146354 44920 182956 44976
rect 146293 44918 182956 44920
rect 146293 44915 146359 44918
rect 182950 44916 182956 44918
rect 183020 44916 183026 44980
rect 135897 44842 135963 44845
rect 181069 44842 181135 44845
rect 135897 44840 181135 44842
rect 135897 44784 135902 44840
rect 135958 44784 181074 44840
rect 181130 44784 181135 44840
rect 135897 44782 181135 44784
rect 135897 44779 135963 44782
rect 181069 44779 181135 44782
rect 185342 44372 185348 44436
rect 185412 44434 185418 44436
rect 190085 44434 190151 44437
rect 185412 44432 190151 44434
rect 185412 44376 190090 44432
rect 190146 44376 190151 44432
rect 185412 44374 190151 44376
rect 185412 44372 185418 44374
rect 190085 44371 190151 44374
rect 136541 43482 136607 43485
rect 133830 43480 136607 43482
rect 133830 43424 136546 43480
rect 136602 43424 136607 43480
rect 133830 43422 136607 43424
rect 133830 42840 133890 43422
rect 136541 43419 136607 43422
rect 144913 43482 144979 43485
rect 183134 43482 183140 43484
rect 144913 43480 183140 43482
rect 144913 43424 144918 43480
rect 144974 43424 183140 43480
rect 144913 43422 183140 43424
rect 144913 43419 144979 43422
rect 183134 43420 183140 43422
rect 183204 43420 183210 43484
rect 190126 43420 190132 43484
rect 190196 43482 190202 43484
rect 247033 43482 247099 43485
rect 190196 43480 247099 43482
rect 190196 43424 247038 43480
rect 247094 43424 247099 43480
rect 190196 43422 247099 43424
rect 190196 43420 190202 43422
rect 247033 43419 247099 43422
rect 188470 42060 188476 42124
rect 188540 42122 188546 42124
rect 230473 42122 230539 42125
rect 188540 42120 230539 42122
rect 188540 42064 230478 42120
rect 230534 42064 230539 42120
rect 188540 42062 230539 42064
rect 188540 42060 188546 42062
rect 230473 42059 230539 42062
rect 170622 41924 170628 41988
rect 170692 41986 170698 41988
rect 580625 41986 580691 41989
rect 170692 41984 580691 41986
rect 170692 41928 580630 41984
rect 580686 41928 580691 41984
rect 170692 41926 580691 41928
rect 170692 41924 170698 41926
rect 580625 41923 580691 41926
rect 200021 41444 200087 41445
rect 166942 41380 166948 41444
rect 167012 41442 167018 41444
rect 167678 41442 167684 41444
rect 167012 41382 167684 41442
rect 167012 41380 167018 41382
rect 167678 41380 167684 41382
rect 167748 41380 167754 41444
rect 200021 41442 200068 41444
rect 199976 41440 200068 41442
rect 199976 41384 200026 41440
rect 199976 41382 200068 41384
rect 200021 41380 200068 41382
rect 200132 41380 200138 41444
rect 200021 41379 200087 41380
rect 170806 41244 170812 41308
rect 170876 41306 170882 41308
rect 552657 41306 552723 41309
rect 170876 41304 552723 41306
rect 170876 41248 552662 41304
rect 552718 41248 552723 41304
rect 170876 41246 552723 41248
rect 170876 41244 170882 41246
rect 552657 41243 552723 41246
rect 170990 41108 170996 41172
rect 171060 41170 171066 41172
rect 550081 41170 550147 41173
rect 171060 41168 550147 41170
rect 171060 41112 550086 41168
rect 550142 41112 550147 41168
rect 171060 41110 550147 41112
rect 171060 41108 171066 41110
rect 550081 41107 550147 41110
rect 136081 40898 136147 40901
rect 133830 40896 136147 40898
rect 133830 40840 136086 40896
rect 136142 40840 136147 40896
rect 133830 40838 136147 40840
rect 133830 40256 133890 40838
rect 136081 40835 136147 40838
rect 136541 37906 136607 37909
rect 133830 37904 136607 37906
rect 133830 37848 136546 37904
rect 136602 37848 136607 37904
rect 133830 37846 136607 37848
rect 133830 37672 133890 37846
rect 136541 37843 136607 37846
rect 147673 37906 147739 37909
rect 182766 37906 182772 37908
rect 147673 37904 182772 37906
rect 147673 37848 147678 37904
rect 147734 37848 182772 37904
rect 147673 37846 182772 37848
rect 147673 37843 147739 37846
rect 182766 37844 182772 37846
rect 182836 37844 182842 37908
rect 195278 37844 195284 37908
rect 195348 37906 195354 37908
rect 318793 37906 318859 37909
rect 195348 37904 318859 37906
rect 195348 37848 318798 37904
rect 318854 37848 318859 37904
rect 195348 37846 318859 37848
rect 195348 37844 195354 37846
rect 318793 37843 318859 37846
rect 191046 36484 191052 36548
rect 191116 36546 191122 36548
rect 266353 36546 266419 36549
rect 191116 36544 266419 36546
rect 191116 36488 266358 36544
rect 266414 36488 266419 36544
rect 191116 36486 266419 36488
rect 191116 36484 191122 36486
rect 266353 36483 266419 36486
rect 200021 36004 200087 36005
rect 200021 36002 200068 36004
rect 199976 36000 200068 36002
rect 200132 36002 200138 36004
rect 199976 35944 200026 36000
rect 199976 35942 200068 35944
rect 200021 35940 200068 35942
rect 200132 35942 200214 36002
rect 200132 35940 200138 35942
rect 200021 35939 200087 35940
rect 192150 35532 192156 35596
rect 192220 35594 192226 35596
rect 285673 35594 285739 35597
rect 192220 35592 285739 35594
rect 192220 35536 285678 35592
rect 285734 35536 285739 35592
rect 192220 35534 285739 35536
rect 192220 35532 192226 35534
rect 285673 35531 285739 35534
rect 136541 35458 136607 35461
rect 133830 35456 136607 35458
rect 133830 35400 136546 35456
rect 136602 35400 136607 35456
rect 133830 35398 136607 35400
rect 133830 35088 133890 35398
rect 136541 35395 136607 35398
rect 200062 35396 200068 35460
rect 200132 35458 200138 35460
rect 390553 35458 390619 35461
rect 200132 35456 390619 35458
rect 200132 35400 390558 35456
rect 390614 35400 390619 35456
rect 200132 35398 390619 35400
rect 200132 35396 200138 35398
rect 390553 35395 390619 35398
rect 209078 35260 209084 35324
rect 209148 35322 209154 35324
rect 498193 35322 498259 35325
rect 209148 35320 498259 35322
rect 209148 35264 498198 35320
rect 498254 35264 498259 35320
rect 209148 35262 498259 35264
rect 209148 35260 209154 35262
rect 498193 35259 498259 35262
rect 149053 35186 149119 35189
rect 182582 35186 182588 35188
rect 149053 35184 182588 35186
rect 149053 35128 149058 35184
rect 149114 35128 182588 35184
rect 149053 35126 182588 35128
rect 149053 35123 149119 35126
rect 182582 35124 182588 35126
rect 182652 35124 182658 35188
rect 213126 35124 213132 35188
rect 213196 35186 213202 35188
rect 549253 35186 549319 35189
rect 213196 35184 549319 35186
rect 213196 35128 549258 35184
rect 549314 35128 549319 35184
rect 213196 35126 549319 35128
rect 213196 35124 213202 35126
rect 549253 35123 549319 35126
rect 193990 34172 193996 34236
rect 194060 34234 194066 34236
rect 303613 34234 303679 34237
rect 194060 34232 303679 34234
rect 194060 34176 303618 34232
rect 303674 34176 303679 34232
rect 194060 34174 303679 34176
rect 194060 34172 194066 34174
rect 303613 34171 303679 34174
rect 202086 34036 202092 34100
rect 202156 34098 202162 34100
rect 407113 34098 407179 34101
rect 202156 34096 407179 34098
rect 202156 34040 407118 34096
rect 407174 34040 407179 34096
rect 202156 34038 407179 34040
rect 202156 34036 202162 34038
rect 407113 34035 407179 34038
rect 210366 33900 210372 33964
rect 210436 33962 210442 33964
rect 514753 33962 514819 33965
rect 210436 33960 514819 33962
rect 210436 33904 514758 33960
rect 514814 33904 514819 33960
rect 210436 33902 514819 33904
rect 210436 33900 210442 33902
rect 514753 33899 514819 33902
rect 211838 33764 211844 33828
rect 211908 33826 211914 33828
rect 532693 33826 532759 33829
rect 211908 33824 532759 33826
rect 211908 33768 532698 33824
rect 532754 33768 532759 33824
rect 211908 33766 532759 33768
rect 211908 33764 211914 33766
rect 532693 33763 532759 33766
rect 580349 33146 580415 33149
rect 583520 33146 584960 33236
rect 580349 33144 584960 33146
rect 580349 33088 580354 33144
rect 580410 33088 584960 33144
rect 580349 33086 584960 33088
rect 580349 33083 580415 33086
rect 136541 33010 136607 33013
rect 133830 33008 136607 33010
rect 133830 32952 136546 33008
rect 136602 32952 136607 33008
rect 583520 32996 584960 33086
rect 133830 32950 136607 32952
rect -960 32466 480 32556
rect 133830 32504 133890 32950
rect 136541 32947 136607 32950
rect 198038 32676 198044 32740
rect 198108 32738 198114 32740
rect 357525 32738 357591 32741
rect 198108 32736 357591 32738
rect 198108 32680 357530 32736
rect 357586 32680 357591 32736
rect 198108 32678 357591 32680
rect 198108 32676 198114 32678
rect 357525 32675 357591 32678
rect 213494 32540 213500 32604
rect 213564 32602 213570 32604
rect 550633 32602 550699 32605
rect 213564 32600 550699 32602
rect 213564 32544 550638 32600
rect 550694 32544 550699 32600
rect 213564 32542 550699 32544
rect 213564 32540 213570 32542
rect 550633 32539 550699 32542
rect 3785 32466 3851 32469
rect -960 32464 3851 32466
rect -960 32408 3790 32464
rect 3846 32408 3851 32464
rect -960 32406 3851 32408
rect -960 32316 480 32406
rect 3785 32403 3851 32406
rect 213310 32404 213316 32468
rect 213380 32466 213386 32468
rect 552013 32466 552079 32469
rect 213380 32464 552079 32466
rect 213380 32408 552018 32464
rect 552074 32408 552079 32464
rect 213380 32406 552079 32408
rect 213380 32404 213386 32406
rect 552013 32403 552079 32406
rect 199326 31044 199332 31108
rect 199396 31106 199402 31108
rect 371233 31106 371299 31109
rect 199396 31104 371299 31106
rect 199396 31048 371238 31104
rect 371294 31048 371299 31104
rect 199396 31046 371299 31048
rect 199396 31044 199402 31046
rect 371233 31043 371299 31046
rect 212022 30908 212028 30972
rect 212092 30970 212098 30972
rect 531313 30970 531379 30973
rect 212092 30968 531379 30970
rect 212092 30912 531318 30968
rect 531374 30912 531379 30968
rect 212092 30910 531379 30912
rect 212092 30908 212098 30910
rect 531313 30907 531379 30910
rect 133830 29474 133890 29920
rect 195462 29820 195468 29884
rect 195532 29882 195538 29884
rect 320173 29882 320239 29885
rect 195532 29880 320239 29882
rect 195532 29824 320178 29880
rect 320234 29824 320239 29880
rect 195532 29822 320239 29824
rect 195532 29820 195538 29822
rect 320173 29819 320239 29822
rect 196198 29684 196204 29748
rect 196268 29746 196274 29748
rect 338113 29746 338179 29749
rect 196268 29744 338179 29746
rect 196268 29688 338118 29744
rect 338174 29688 338179 29744
rect 196268 29686 338179 29688
rect 196268 29684 196274 29686
rect 338113 29683 338179 29686
rect 203190 29548 203196 29612
rect 203260 29610 203266 29612
rect 423673 29610 423739 29613
rect 203260 29608 423739 29610
rect 203260 29552 423678 29608
rect 423734 29552 423739 29608
rect 203260 29550 423739 29552
rect 203260 29548 203266 29550
rect 423673 29547 423739 29550
rect 135437 29474 135503 29477
rect 133830 29472 135503 29474
rect 133830 29416 135442 29472
rect 135498 29416 135503 29472
rect 133830 29414 135503 29416
rect 135437 29411 135503 29414
rect 199510 28460 199516 28524
rect 199580 28522 199586 28524
rect 373993 28522 374059 28525
rect 199580 28520 374059 28522
rect 199580 28464 373998 28520
rect 374054 28464 374059 28520
rect 199580 28462 374059 28464
rect 199580 28460 199586 28462
rect 373993 28459 374059 28462
rect 210734 28324 210740 28388
rect 210804 28386 210810 28388
rect 513373 28386 513439 28389
rect 210804 28384 513439 28386
rect 210804 28328 513378 28384
rect 513434 28328 513439 28384
rect 210804 28326 513439 28328
rect 210804 28324 210810 28326
rect 513373 28323 513439 28326
rect 210550 28188 210556 28252
rect 210620 28250 210626 28252
rect 516133 28250 516199 28253
rect 210620 28248 516199 28250
rect 210620 28192 516138 28248
rect 516194 28192 516199 28248
rect 210620 28190 516199 28192
rect 210620 28188 210626 28190
rect 516133 28187 516199 28190
rect 136541 27570 136607 27573
rect 133830 27568 136607 27570
rect 133830 27512 136546 27568
rect 136602 27512 136607 27568
rect 133830 27510 136607 27512
rect 133830 27336 133890 27510
rect 136541 27507 136607 27510
rect 205030 26964 205036 27028
rect 205100 27026 205106 27028
rect 445753 27026 445819 27029
rect 205100 27024 445819 27026
rect 205100 26968 445758 27024
rect 445814 26968 445819 27024
rect 205100 26966 445819 26968
rect 205100 26964 205106 26966
rect 445753 26963 445819 26966
rect 209262 26828 209268 26892
rect 209332 26890 209338 26892
rect 498285 26890 498351 26893
rect 209332 26888 498351 26890
rect 209332 26832 498290 26888
rect 498346 26832 498351 26888
rect 209332 26830 498351 26832
rect 209332 26828 209338 26830
rect 498285 26827 498351 26830
rect 214598 25604 214604 25668
rect 214668 25666 214674 25668
rect 569953 25666 570019 25669
rect 214668 25664 570019 25666
rect 214668 25608 569958 25664
rect 570014 25608 570019 25664
rect 214668 25606 570019 25608
rect 214668 25604 214674 25606
rect 569953 25603 570019 25606
rect 180190 25468 180196 25532
rect 180260 25530 180266 25532
rect 580993 25530 581059 25533
rect 180260 25528 581059 25530
rect 180260 25472 580998 25528
rect 581054 25472 581059 25528
rect 180260 25470 581059 25472
rect 180260 25468 180266 25470
rect 580993 25467 581059 25470
rect 22737 24850 22803 24853
rect 177665 24850 177731 24853
rect 22737 24848 177731 24850
rect 22737 24792 22742 24848
rect 22798 24792 177670 24848
rect 177726 24792 177731 24848
rect 22737 24790 177731 24792
rect 22737 24787 22803 24790
rect 177665 24787 177731 24790
rect 192334 24380 192340 24444
rect 192404 24442 192410 24444
rect 284293 24442 284359 24445
rect 192404 24440 284359 24442
rect 192404 24384 284298 24440
rect 284354 24384 284359 24440
rect 192404 24382 284359 24384
rect 192404 24380 192410 24382
rect 284293 24379 284359 24382
rect 209446 24244 209452 24308
rect 209516 24306 209522 24308
rect 496813 24306 496879 24309
rect 209516 24304 496879 24306
rect 209516 24248 496818 24304
rect 496874 24248 496879 24304
rect 209516 24246 496879 24248
rect 209516 24244 209522 24246
rect 496813 24243 496879 24246
rect 18597 24170 18663 24173
rect 160737 24170 160803 24173
rect 18597 24168 160803 24170
rect 18597 24112 18602 24168
rect 18658 24112 160742 24168
rect 160798 24112 160803 24168
rect 18597 24110 160803 24112
rect 18597 24107 18663 24110
rect 160737 24107 160803 24110
rect 214782 24108 214788 24172
rect 214852 24170 214858 24172
rect 568573 24170 568639 24173
rect 214852 24168 568639 24170
rect 214852 24112 568578 24168
rect 568634 24112 568639 24168
rect 214852 24110 568639 24112
rect 214852 24108 214858 24110
rect 568573 24107 568639 24110
rect 19333 22674 19399 22677
rect 161974 22674 161980 22676
rect 19333 22672 161980 22674
rect 19333 22616 19338 22672
rect 19394 22616 161980 22672
rect 19333 22614 161980 22616
rect 19333 22611 19399 22614
rect 161974 22612 161980 22614
rect 162044 22612 162050 22676
rect 196382 21796 196388 21860
rect 196452 21858 196458 21860
rect 336733 21858 336799 21861
rect 196452 21856 336799 21858
rect 196452 21800 336738 21856
rect 336794 21800 336799 21856
rect 196452 21798 336799 21800
rect 196452 21796 196458 21798
rect 336733 21795 336799 21798
rect 198222 21660 198228 21724
rect 198292 21722 198298 21724
rect 353293 21722 353359 21725
rect 198292 21720 353359 21722
rect 198292 21664 353298 21720
rect 353354 21664 353359 21720
rect 198292 21662 353359 21664
rect 198292 21660 198298 21662
rect 353293 21659 353359 21662
rect 199694 21524 199700 21588
rect 199764 21586 199770 21588
rect 374085 21586 374151 21589
rect 199764 21584 374151 21586
rect 199764 21528 374090 21584
rect 374146 21528 374151 21584
rect 199764 21526 374151 21528
rect 199764 21524 199770 21526
rect 374085 21523 374151 21526
rect 93853 21450 93919 21453
rect 167310 21450 167316 21452
rect 93853 21448 167316 21450
rect 93853 21392 93858 21448
rect 93914 21392 167316 21448
rect 93853 21390 167316 21392
rect 93853 21387 93919 21390
rect 167310 21388 167316 21390
rect 167380 21388 167386 21452
rect 185158 21388 185164 21452
rect 185228 21450 185234 21452
rect 196065 21450 196131 21453
rect 185228 21448 196131 21450
rect 185228 21392 196070 21448
rect 196126 21392 196131 21448
rect 185228 21390 196131 21392
rect 185228 21388 185234 21390
rect 196065 21387 196131 21390
rect 203374 21388 203380 21452
rect 203444 21450 203450 21452
rect 426433 21450 426499 21453
rect 203444 21448 426499 21450
rect 203444 21392 426438 21448
rect 426494 21392 426499 21448
rect 203444 21390 426499 21392
rect 203444 21388 203450 21390
rect 426433 21387 426499 21390
rect 1393 21314 1459 21317
rect 160318 21314 160324 21316
rect 1393 21312 160324 21314
rect 1393 21256 1398 21312
rect 1454 21256 160324 21312
rect 1393 21254 160324 21256
rect 1393 21251 1459 21254
rect 160318 21252 160324 21254
rect 160388 21252 160394 21316
rect 180374 21252 180380 21316
rect 180444 21314 180450 21316
rect 581085 21314 581151 21317
rect 180444 21312 581151 21314
rect 180444 21256 581090 21312
rect 581146 21256 581151 21312
rect 180444 21254 581151 21256
rect 180444 21252 180450 21254
rect 581085 21251 581151 21254
rect 202270 20028 202276 20092
rect 202340 20090 202346 20092
rect 407205 20090 407271 20093
rect 202340 20088 407271 20090
rect 202340 20032 407210 20088
rect 407266 20032 407271 20088
rect 202340 20030 407271 20032
rect 202340 20028 202346 20030
rect 407205 20027 407271 20030
rect 205214 19892 205220 19956
rect 205284 19954 205290 19956
rect 442993 19954 443059 19957
rect 205284 19952 443059 19954
rect 205284 19896 442998 19952
rect 443054 19896 443059 19952
rect 205284 19894 443059 19896
rect 205284 19892 205290 19894
rect 442993 19891 443059 19894
rect 580257 19818 580323 19821
rect 583520 19818 584960 19908
rect 580257 19816 584960 19818
rect 580257 19760 580262 19816
rect 580318 19760 584960 19816
rect 580257 19758 584960 19760
rect 580257 19755 580323 19758
rect 583520 19668 584960 19758
rect -960 19410 480 19500
rect 3417 19410 3483 19413
rect -960 19408 3483 19410
rect -960 19352 3422 19408
rect 3478 19352 3483 19408
rect -960 19350 3483 19352
rect -960 19260 480 19350
rect 3417 19347 3483 19350
rect 131113 18866 131179 18869
rect 181110 18866 181116 18868
rect 131113 18864 181116 18866
rect 131113 18808 131118 18864
rect 131174 18808 181116 18864
rect 131113 18806 181116 18808
rect 131113 18803 131179 18806
rect 181110 18804 181116 18806
rect 181180 18804 181186 18868
rect 129733 18730 129799 18733
rect 180926 18730 180932 18732
rect 129733 18728 180932 18730
rect 129733 18672 129738 18728
rect 129794 18672 180932 18728
rect 129733 18670 180932 18672
rect 129733 18667 129799 18670
rect 180926 18668 180932 18670
rect 180996 18668 181002 18732
rect 20713 18594 20779 18597
rect 161790 18594 161796 18596
rect 20713 18592 161796 18594
rect 20713 18536 20718 18592
rect 20774 18536 161796 18592
rect 20713 18534 161796 18536
rect 20713 18531 20779 18534
rect 161790 18532 161796 18534
rect 161860 18532 161866 18596
rect 194174 18532 194180 18596
rect 194244 18594 194250 18596
rect 300853 18594 300919 18597
rect 194244 18592 300919 18594
rect 194244 18536 300858 18592
rect 300914 18536 300919 18592
rect 194244 18534 300919 18536
rect 194244 18532 194250 18534
rect 300853 18531 300919 18534
rect 187182 17716 187188 17780
rect 187252 17778 187258 17780
rect 211797 17778 211863 17781
rect 187252 17776 211863 17778
rect 187252 17720 211802 17776
rect 211858 17720 211863 17776
rect 187252 17718 211863 17720
rect 187252 17716 187258 17718
rect 211797 17715 211863 17718
rect 192518 17580 192524 17644
rect 192588 17642 192594 17644
rect 284385 17642 284451 17645
rect 192588 17640 284451 17642
rect 192588 17584 284390 17640
rect 284446 17584 284451 17640
rect 192588 17582 284451 17584
rect 192588 17580 192594 17582
rect 284385 17579 284451 17582
rect 206502 17444 206508 17508
rect 206572 17506 206578 17508
rect 463693 17506 463759 17509
rect 206572 17504 463759 17506
rect 206572 17448 463698 17504
rect 463754 17448 463759 17504
rect 206572 17446 463759 17448
rect 206572 17444 206578 17446
rect 463693 17443 463759 17446
rect 127065 17370 127131 17373
rect 181294 17370 181300 17372
rect 127065 17368 181300 17370
rect 127065 17312 127070 17368
rect 127126 17312 181300 17368
rect 127065 17310 181300 17312
rect 127065 17307 127131 17310
rect 181294 17308 181300 17310
rect 181364 17308 181370 17372
rect 207238 17308 207244 17372
rect 207308 17370 207314 17372
rect 477493 17370 477559 17373
rect 207308 17368 477559 17370
rect 207308 17312 477498 17368
rect 477554 17312 477559 17368
rect 207308 17310 477559 17312
rect 207308 17308 207314 17310
rect 477493 17307 477559 17310
rect 75913 17234 75979 17237
rect 166206 17234 166212 17236
rect 75913 17232 166212 17234
rect 75913 17176 75918 17232
rect 75974 17176 166212 17232
rect 75913 17174 166212 17176
rect 75913 17171 75979 17174
rect 166206 17172 166212 17174
rect 166276 17172 166282 17236
rect 187366 17172 187372 17236
rect 187436 17234 187442 17236
rect 210417 17234 210483 17237
rect 187436 17232 210483 17234
rect 187436 17176 210422 17232
rect 210478 17176 210483 17232
rect 187436 17174 210483 17176
rect 187436 17172 187442 17174
rect 210417 17171 210483 17174
rect 210918 17172 210924 17236
rect 210988 17234 210994 17236
rect 514845 17234 514911 17237
rect 210988 17232 514911 17234
rect 210988 17176 514850 17232
rect 514906 17176 514911 17232
rect 210988 17174 514911 17176
rect 210988 17172 210994 17174
rect 514845 17171 514911 17174
rect 198406 15948 198412 16012
rect 198476 16010 198482 16012
rect 355225 16010 355291 16013
rect 198476 16008 355291 16010
rect 198476 15952 355230 16008
rect 355286 15952 355291 16008
rect 198476 15950 355291 15952
rect 198476 15948 198482 15950
rect 355225 15947 355291 15950
rect 41873 15874 41939 15877
rect 163446 15874 163452 15876
rect 41873 15872 163452 15874
rect 41873 15816 41878 15872
rect 41934 15816 163452 15872
rect 41873 15814 163452 15816
rect 41873 15811 41939 15814
rect 163446 15812 163452 15814
rect 163516 15812 163522 15876
rect 203558 15812 203564 15876
rect 203628 15874 203634 15876
rect 428457 15874 428523 15877
rect 203628 15872 428523 15874
rect 203628 15816 428462 15872
rect 428518 15816 428523 15872
rect 203628 15814 428523 15816
rect 203628 15812 203634 15814
rect 428457 15811 428523 15814
rect 180558 14724 180564 14788
rect 180628 14786 180634 14788
rect 271137 14786 271203 14789
rect 180628 14784 271203 14786
rect 180628 14728 271142 14784
rect 271198 14728 271203 14784
rect 180628 14726 271203 14728
rect 180628 14724 180634 14726
rect 271137 14723 271203 14726
rect 91553 14650 91619 14653
rect 167126 14650 167132 14652
rect 91553 14648 167132 14650
rect 91553 14592 91558 14648
rect 91614 14592 167132 14648
rect 91553 14590 167132 14592
rect 91553 14587 91619 14590
rect 167126 14588 167132 14590
rect 167196 14588 167202 14652
rect 195646 14588 195652 14652
rect 195716 14650 195722 14652
rect 322105 14650 322171 14653
rect 195716 14648 322171 14650
rect 195716 14592 322110 14648
rect 322166 14592 322171 14648
rect 195716 14590 322171 14592
rect 195716 14588 195722 14590
rect 322105 14587 322171 14590
rect 77293 14514 77359 14517
rect 166022 14514 166028 14516
rect 77293 14512 166028 14514
rect 77293 14456 77298 14512
rect 77354 14456 166028 14512
rect 77293 14454 166028 14456
rect 77293 14451 77359 14454
rect 166022 14452 166028 14454
rect 166092 14452 166098 14516
rect 202454 14452 202460 14516
rect 202524 14514 202530 14516
rect 410793 14514 410859 14517
rect 202524 14512 410859 14514
rect 202524 14456 410798 14512
rect 410854 14456 410859 14512
rect 202524 14454 410859 14456
rect 202524 14452 202530 14454
rect 410793 14451 410859 14454
rect 191230 13500 191236 13564
rect 191300 13562 191306 13564
rect 264973 13562 265039 13565
rect 191300 13560 265039 13562
rect 191300 13504 264978 13560
rect 265034 13504 265039 13560
rect 191300 13502 265039 13504
rect 191300 13500 191306 13502
rect 264973 13499 265039 13502
rect 191414 13364 191420 13428
rect 191484 13426 191490 13428
rect 268377 13426 268443 13429
rect 191484 13424 268443 13426
rect 191484 13368 268382 13424
rect 268438 13368 268443 13424
rect 191484 13366 268443 13368
rect 191484 13364 191490 13366
rect 268377 13363 268443 13366
rect 192702 13228 192708 13292
rect 192772 13290 192778 13292
rect 283097 13290 283163 13293
rect 192772 13288 283163 13290
rect 192772 13232 283102 13288
rect 283158 13232 283163 13288
rect 192772 13230 283163 13232
rect 192772 13228 192778 13230
rect 283097 13227 283163 13230
rect 94681 13154 94747 13157
rect 166942 13154 166948 13156
rect 94681 13152 166948 13154
rect 94681 13096 94686 13152
rect 94742 13096 166948 13152
rect 94681 13094 166948 13096
rect 94681 13091 94747 13094
rect 166942 13092 166948 13094
rect 167012 13092 167018 13156
rect 195830 13092 195836 13156
rect 195900 13154 195906 13156
rect 318057 13154 318123 13157
rect 195900 13152 318123 13154
rect 195900 13096 318062 13152
rect 318118 13096 318123 13152
rect 195900 13094 318123 13096
rect 195900 13092 195906 13094
rect 318057 13091 318123 13094
rect 74993 13018 75059 13021
rect 165838 13018 165844 13020
rect 74993 13016 165844 13018
rect 74993 12960 74998 13016
rect 75054 12960 165844 13016
rect 74993 12958 165844 12960
rect 74993 12955 75059 12958
rect 165838 12956 165844 12958
rect 165908 12956 165914 13020
rect 201350 12956 201356 13020
rect 201420 13018 201426 13020
rect 392577 13018 392643 13021
rect 201420 13016 392643 13018
rect 201420 12960 392582 13016
rect 392638 12960 392643 13016
rect 201420 12958 392643 12960
rect 201420 12956 201426 12958
rect 392577 12955 392643 12958
rect 206686 12004 206692 12068
rect 206756 12066 206762 12068
rect 462313 12066 462379 12069
rect 206756 12064 462379 12066
rect 206756 12008 462318 12064
rect 462374 12008 462379 12064
rect 206756 12006 462379 12008
rect 206756 12004 206762 12006
rect 462313 12003 462379 12006
rect 212206 11868 212212 11932
rect 212276 11930 212282 11932
rect 531405 11930 531471 11933
rect 212276 11928 531471 11930
rect 212276 11872 531410 11928
rect 531466 11872 531471 11928
rect 212276 11870 531471 11872
rect 212276 11868 212282 11870
rect 531405 11867 531471 11870
rect 212390 11732 212396 11796
rect 212460 11794 212466 11796
rect 534441 11794 534507 11797
rect 212460 11792 534507 11794
rect 212460 11736 534446 11792
rect 534502 11736 534507 11792
rect 212460 11734 534507 11736
rect 212460 11732 212466 11734
rect 534441 11731 534507 11734
rect 3601 11658 3667 11661
rect 160134 11658 160140 11660
rect 3601 11656 160140 11658
rect 3601 11600 3606 11656
rect 3662 11600 160140 11656
rect 3601 11598 160140 11600
rect 3601 11595 3667 11598
rect 160134 11596 160140 11598
rect 160204 11596 160210 11660
rect 214966 11596 214972 11660
rect 215036 11658 215042 11660
rect 567561 11658 567627 11661
rect 215036 11656 567627 11658
rect 215036 11600 567566 11656
rect 567622 11600 567627 11656
rect 215036 11598 567627 11600
rect 215036 11596 215042 11598
rect 567561 11595 567627 11598
rect 36721 10298 36787 10301
rect 163262 10298 163268 10300
rect 36721 10296 163268 10298
rect 36721 10240 36726 10296
rect 36782 10240 163268 10296
rect 36721 10238 163268 10240
rect 36721 10235 36787 10238
rect 163262 10236 163268 10238
rect 163332 10236 163338 10300
rect 209630 10236 209636 10300
rect 209700 10298 209706 10300
rect 495433 10298 495499 10301
rect 209700 10296 495499 10298
rect 209700 10240 495438 10296
rect 495494 10240 495499 10296
rect 209700 10238 495499 10240
rect 209700 10236 209706 10238
rect 495433 10235 495499 10238
rect 112805 9210 112871 9213
rect 169150 9210 169156 9212
rect 112805 9208 169156 9210
rect 112805 9152 112810 9208
rect 112866 9152 169156 9208
rect 112805 9150 169156 9152
rect 112805 9147 112871 9150
rect 169150 9148 169156 9150
rect 169220 9148 169226 9212
rect 109309 9074 109375 9077
rect 169334 9074 169340 9076
rect 109309 9072 169340 9074
rect 109309 9016 109314 9072
rect 109370 9016 169340 9072
rect 109309 9014 169340 9016
rect 109309 9011 109375 9014
rect 169334 9012 169340 9014
rect 169404 9012 169410 9076
rect 205398 9012 205404 9076
rect 205468 9074 205474 9076
rect 445017 9074 445083 9077
rect 205468 9072 445083 9074
rect 205468 9016 445022 9072
rect 445078 9016 445083 9072
rect 205468 9014 445083 9016
rect 205468 9012 205474 9014
rect 445017 9011 445083 9014
rect 23013 8938 23079 8941
rect 161606 8938 161612 8940
rect 23013 8936 161612 8938
rect 23013 8880 23018 8936
rect 23074 8880 161612 8936
rect 23013 8878 161612 8880
rect 23013 8875 23079 8878
rect 161606 8876 161612 8878
rect 161676 8876 161682 8940
rect 213678 8876 213684 8940
rect 213748 8938 213754 8940
rect 549069 8938 549135 8941
rect 213748 8936 549135 8938
rect 213748 8880 549074 8936
rect 549130 8880 549135 8936
rect 213748 8878 549135 8880
rect 213748 8876 213754 8878
rect 549069 8875 549135 8878
rect 190310 6836 190316 6900
rect 190380 6898 190386 6900
rect 251265 6898 251331 6901
rect 190380 6896 251331 6898
rect 190380 6840 251270 6896
rect 251326 6840 251331 6896
rect 190380 6838 251331 6840
rect 190380 6836 190386 6838
rect 251265 6835 251331 6838
rect 194358 6700 194364 6764
rect 194428 6762 194434 6764
rect 303153 6762 303219 6765
rect 194428 6760 303219 6762
rect 194428 6704 303158 6760
rect 303214 6704 303219 6760
rect 194428 6702 303219 6704
rect 194428 6700 194434 6702
rect 303153 6699 303219 6702
rect -960 6490 480 6580
rect 198590 6564 198596 6628
rect 198660 6626 198666 6628
rect 356329 6626 356395 6629
rect 198660 6624 356395 6626
rect 198660 6568 356334 6624
rect 356390 6568 356395 6624
rect 198660 6566 356395 6568
rect 198660 6564 198666 6566
rect 356329 6563 356395 6566
rect 580165 6626 580231 6629
rect 583520 6626 584960 6716
rect 580165 6624 584960 6626
rect 580165 6568 580170 6624
rect 580226 6568 584960 6624
rect 580165 6566 584960 6568
rect 580165 6563 580231 6566
rect 3417 6490 3483 6493
rect -960 6488 3483 6490
rect -960 6432 3422 6488
rect 3478 6432 3483 6488
rect -960 6430 3483 6432
rect -960 6340 480 6430
rect 3417 6427 3483 6430
rect 199878 6428 199884 6492
rect 199948 6490 199954 6492
rect 370589 6490 370655 6493
rect 199948 6488 370655 6490
rect 199948 6432 370594 6488
rect 370650 6432 370655 6488
rect 583520 6476 584960 6566
rect 199948 6430 370655 6432
rect 199948 6428 199954 6430
rect 370589 6427 370655 6430
rect 40677 6354 40743 6357
rect 163078 6354 163084 6356
rect 40677 6352 163084 6354
rect 40677 6296 40682 6352
rect 40738 6296 163084 6352
rect 40677 6294 163084 6296
rect 40677 6291 40743 6294
rect 163078 6292 163084 6294
rect 163148 6292 163154 6356
rect 202638 6292 202644 6356
rect 202708 6354 202714 6356
rect 409597 6354 409663 6357
rect 202708 6352 409663 6354
rect 202708 6296 409602 6352
rect 409658 6296 409663 6352
rect 202708 6294 409663 6296
rect 202708 6292 202714 6294
rect 409597 6291 409663 6294
rect 38377 6218 38443 6221
rect 162894 6218 162900 6220
rect 38377 6216 162900 6218
rect 38377 6160 38382 6216
rect 38438 6160 162900 6216
rect 38377 6158 162900 6160
rect 38377 6155 38443 6158
rect 162894 6156 162900 6158
rect 162964 6156 162970 6220
rect 163681 6218 163747 6221
rect 183686 6218 183692 6220
rect 163681 6216 183692 6218
rect 163681 6160 163686 6216
rect 163742 6160 183692 6216
rect 163681 6158 183692 6160
rect 163681 6155 163747 6158
rect 183686 6156 183692 6158
rect 183756 6156 183762 6220
rect 207422 6156 207428 6220
rect 207492 6218 207498 6220
rect 481725 6218 481791 6221
rect 207492 6216 481791 6218
rect 207492 6160 481730 6216
rect 481786 6160 481791 6216
rect 207492 6158 481791 6160
rect 207492 6156 207498 6158
rect 481725 6155 481791 6158
rect 188654 6020 188660 6084
rect 188724 6082 188730 6084
rect 233417 6082 233483 6085
rect 188724 6080 233483 6082
rect 188724 6024 233422 6080
rect 233478 6024 233483 6080
rect 188724 6022 233483 6024
rect 188724 6020 188730 6022
rect 233417 6019 233483 6022
rect 111609 5130 111675 5133
rect 168966 5130 168972 5132
rect 111609 5128 168972 5130
rect 111609 5072 111614 5128
rect 111670 5072 168972 5128
rect 111609 5070 168972 5072
rect 111609 5067 111675 5070
rect 168966 5068 168972 5070
rect 169036 5068 169042 5132
rect 73797 4994 73863 4997
rect 165654 4994 165660 4996
rect 73797 4992 165660 4994
rect 73797 4936 73802 4992
rect 73858 4936 165660 4992
rect 73797 4934 165660 4936
rect 73797 4931 73863 4934
rect 165654 4932 165660 4934
rect 165724 4932 165730 4996
rect 203742 4932 203748 4996
rect 203812 4994 203818 4996
rect 423765 4994 423831 4997
rect 203812 4992 423831 4994
rect 203812 4936 423770 4992
rect 423826 4936 423831 4992
rect 203812 4934 423831 4936
rect 203812 4932 203818 4934
rect 423765 4931 423831 4934
rect 56041 4858 56107 4861
rect 165286 4858 165292 4860
rect 56041 4856 165292 4858
rect 56041 4800 56046 4856
rect 56102 4800 165292 4856
rect 56041 4798 165292 4800
rect 56041 4795 56107 4798
rect 165286 4796 165292 4798
rect 165356 4796 165362 4860
rect 167177 4858 167243 4861
rect 183870 4858 183876 4860
rect 167177 4856 183876 4858
rect 167177 4800 167182 4856
rect 167238 4800 183876 4856
rect 167177 4798 183876 4800
rect 167177 4795 167243 4798
rect 183870 4796 183876 4798
rect 183940 4796 183946 4860
rect 187550 4796 187556 4860
rect 187620 4858 187626 4860
rect 207013 4858 207079 4861
rect 187620 4856 207079 4858
rect 187620 4800 207018 4856
rect 207074 4800 207079 4856
rect 187620 4798 207079 4800
rect 187620 4796 187626 4798
rect 207013 4795 207079 4798
rect 214414 4796 214420 4860
rect 214484 4858 214490 4860
rect 566825 4858 566891 4861
rect 214484 4856 566891 4858
rect 214484 4800 566830 4856
rect 566886 4800 566891 4856
rect 214484 4798 566891 4800
rect 214484 4796 214490 4798
rect 566825 4795 566891 4798
rect 190545 4042 190611 4045
rect 260649 4042 260715 4045
rect 190545 4040 260715 4042
rect 190545 3984 190550 4040
rect 190606 3984 260654 4040
rect 260710 3984 260715 4040
rect 190545 3982 260715 3984
rect 190545 3979 190611 3982
rect 260649 3979 260715 3982
rect 190729 3906 190795 3909
rect 264145 3906 264211 3909
rect 190729 3904 264211 3906
rect 190729 3848 190734 3904
rect 190790 3848 264150 3904
rect 264206 3848 264211 3904
rect 190729 3846 264211 3848
rect 190729 3843 190795 3846
rect 264145 3843 264211 3846
rect 191598 3708 191604 3772
rect 191668 3770 191674 3772
rect 267733 3770 267799 3773
rect 191668 3768 267799 3770
rect 191668 3712 267738 3768
rect 267794 3712 267799 3768
rect 191668 3710 267799 3712
rect 191668 3708 191674 3710
rect 267733 3707 267799 3710
rect 188838 3572 188844 3636
rect 188908 3634 188914 3636
rect 278313 3634 278379 3637
rect 188908 3632 278379 3634
rect 188908 3576 278318 3632
rect 278374 3576 278379 3632
rect 188908 3574 278379 3576
rect 188908 3572 188914 3574
rect 278313 3571 278379 3574
rect 258574 3436 258580 3500
rect 258644 3498 258650 3500
rect 519537 3498 519603 3501
rect 258644 3496 519603 3498
rect 258644 3440 519542 3496
rect 519598 3440 519603 3496
rect 258644 3438 519603 3440
rect 258644 3436 258650 3438
rect 519537 3435 519603 3438
rect 206318 3300 206324 3364
rect 206388 3362 206394 3364
rect 468661 3362 468727 3365
rect 206388 3360 468727 3362
rect 206388 3304 468666 3360
rect 468722 3304 468727 3360
rect 206388 3302 468727 3304
rect 206388 3300 206394 3302
rect 468661 3299 468727 3302
<< via3 >>
rect 251772 670652 251836 670716
rect 224172 300324 224236 300388
rect 155356 293116 155420 293180
rect 155356 171124 155420 171188
rect 224172 122844 224236 122908
rect 208716 52804 208780 52868
rect 173572 52668 173636 52732
rect 251772 52668 251836 52732
rect 169892 52260 169956 52324
rect 161796 51988 161860 52052
rect 163636 51988 163700 52052
rect 160324 51912 160388 51916
rect 160324 51856 160328 51912
rect 160328 51856 160384 51912
rect 160384 51856 160388 51912
rect 160324 51852 160388 51856
rect 161428 51852 161492 51916
rect 162164 51852 162228 51916
rect 162716 51912 162780 51916
rect 162716 51856 162720 51912
rect 162720 51856 162776 51912
rect 162776 51856 162780 51912
rect 160140 51776 160204 51780
rect 160140 51720 160190 51776
rect 160190 51720 160204 51776
rect 160140 51716 160204 51720
rect 161612 51580 161676 51644
rect 162716 51852 162780 51856
rect 162900 51716 162964 51780
rect 163820 51444 163884 51508
rect 165844 51890 165848 51916
rect 165848 51890 165904 51916
rect 165904 51890 165908 51916
rect 165844 51852 165908 51890
rect 166028 51716 166092 51780
rect 167500 51852 167564 51916
rect 169156 51988 169220 52052
rect 174308 51988 174372 52052
rect 166764 51776 166828 51780
rect 166764 51720 166768 51776
rect 166768 51720 166824 51776
rect 166824 51720 166828 51776
rect 166764 51716 166828 51720
rect 169708 51890 169712 51916
rect 169712 51890 169768 51916
rect 169768 51890 169772 51916
rect 169708 51852 169772 51890
rect 170444 51852 170508 51916
rect 170076 51776 170140 51780
rect 170076 51720 170080 51776
rect 170080 51720 170136 51776
rect 170136 51720 170140 51776
rect 170076 51716 170140 51720
rect 168972 51444 169036 51508
rect 169892 51444 169956 51508
rect 173388 51852 173452 51916
rect 173756 51912 173820 51916
rect 173756 51856 173760 51912
rect 173760 51856 173816 51912
rect 173816 51856 173820 51912
rect 173756 51852 173820 51856
rect 174124 51852 174188 51916
rect 175964 51988 176028 52052
rect 174860 51912 174924 51916
rect 174860 51856 174864 51912
rect 174864 51856 174920 51912
rect 174920 51856 174924 51912
rect 174860 51852 174924 51856
rect 176332 51852 176396 51916
rect 177988 51912 178052 51916
rect 177988 51856 177992 51912
rect 177992 51856 178048 51912
rect 178048 51856 178052 51912
rect 177988 51852 178052 51856
rect 178908 51912 178972 51916
rect 178908 51856 178912 51912
rect 178912 51856 178968 51912
rect 178968 51856 178972 51912
rect 178908 51852 178972 51856
rect 180012 51852 180076 51916
rect 180380 51912 180444 51916
rect 180380 51856 180384 51912
rect 180384 51856 180440 51912
rect 180440 51856 180444 51912
rect 180380 51852 180444 51856
rect 180932 51852 180996 51916
rect 181300 51890 181304 51916
rect 181304 51890 181360 51916
rect 181360 51890 181364 51916
rect 181300 51852 181364 51890
rect 182772 51852 182836 51916
rect 182956 51890 182960 51916
rect 182960 51890 183016 51916
rect 183016 51890 183020 51916
rect 182956 51852 183020 51890
rect 183876 51852 183940 51916
rect 184428 51852 184492 51916
rect 184612 51912 184676 51916
rect 184612 51856 184616 51912
rect 184616 51856 184672 51912
rect 184672 51856 184676 51912
rect 184612 51852 184676 51856
rect 185348 51852 185412 51916
rect 187004 51912 187068 51916
rect 187004 51856 187008 51912
rect 187008 51856 187064 51912
rect 187064 51856 187068 51912
rect 187004 51852 187068 51856
rect 188476 51852 188540 51916
rect 189028 51852 189092 51916
rect 192708 51852 192772 51916
rect 194364 52260 194428 52324
rect 194548 52260 194612 52324
rect 194916 52260 194980 52324
rect 193812 52124 193876 52188
rect 194732 52124 194796 52188
rect 194548 51988 194612 52052
rect 196204 51988 196268 52052
rect 208716 52260 208780 52324
rect 204852 52124 204916 52188
rect 194180 51852 194244 51916
rect 195100 51912 195164 51916
rect 195100 51856 195104 51912
rect 195104 51856 195160 51912
rect 195160 51856 195164 51912
rect 195100 51852 195164 51856
rect 195652 51852 195716 51916
rect 196388 51852 196452 51916
rect 205588 52124 205652 52188
rect 207244 51988 207308 52052
rect 198228 51852 198292 51916
rect 198596 51890 198600 51916
rect 198600 51890 198656 51916
rect 198656 51890 198660 51916
rect 198596 51852 198660 51890
rect 200068 51852 200132 51916
rect 202092 51852 202156 51916
rect 203380 51852 203444 51916
rect 205036 51852 205100 51916
rect 205404 51912 205468 51916
rect 205404 51856 205408 51912
rect 205408 51856 205464 51912
rect 205464 51856 205468 51912
rect 205404 51852 205468 51856
rect 205772 51886 205836 51950
rect 206324 51890 206328 51916
rect 206328 51890 206384 51916
rect 206384 51890 206388 51916
rect 206324 51852 206388 51890
rect 206692 51852 206756 51916
rect 207060 51912 207124 51916
rect 207060 51856 207064 51912
rect 207064 51856 207120 51912
rect 207120 51856 207124 51912
rect 207060 51852 207124 51856
rect 207428 51852 207492 51916
rect 173020 51716 173084 51780
rect 174492 51776 174556 51780
rect 174492 51720 174506 51776
rect 174506 51720 174556 51776
rect 174492 51716 174556 51720
rect 175412 51716 175476 51780
rect 205588 51716 205652 51780
rect 206508 51716 206572 51780
rect 207612 51776 207676 51780
rect 207612 51720 207616 51776
rect 207616 51720 207672 51776
rect 207672 51720 207676 51776
rect 207612 51716 207676 51720
rect 209084 51988 209148 52052
rect 209268 51912 209332 51916
rect 209268 51856 209272 51912
rect 209272 51856 209328 51912
rect 209328 51856 209332 51912
rect 209268 51852 209332 51856
rect 209452 51852 209516 51916
rect 210556 51912 210620 51916
rect 210556 51856 210560 51912
rect 210560 51856 210616 51912
rect 210616 51856 210620 51912
rect 210556 51852 210620 51856
rect 210924 51912 210988 51916
rect 210924 51856 210928 51912
rect 210928 51856 210984 51912
rect 210984 51856 210988 51912
rect 210924 51852 210988 51856
rect 210188 51716 210252 51780
rect 210556 51716 210620 51780
rect 212028 51852 212092 51916
rect 213500 51852 213564 51916
rect 214052 51852 214116 51916
rect 215524 51890 215528 51916
rect 215528 51890 215584 51916
rect 215584 51890 215588 51916
rect 215524 51852 215588 51890
rect 211660 51776 211724 51780
rect 211660 51720 211664 51776
rect 211664 51720 211720 51776
rect 211720 51720 211724 51776
rect 211660 51716 211724 51720
rect 212212 51776 212276 51780
rect 212212 51720 212216 51776
rect 212216 51720 212272 51776
rect 212272 51720 212276 51776
rect 212212 51716 212276 51720
rect 212396 51716 212460 51780
rect 214236 51716 214300 51780
rect 173204 51580 173268 51644
rect 173572 51444 173636 51508
rect 173204 51308 173268 51372
rect 174492 51172 174556 51236
rect 174860 51036 174924 51100
rect 175412 51036 175476 51100
rect 173388 50900 173452 50964
rect 170812 50764 170876 50828
rect 173756 50628 173820 50692
rect 175964 50356 176028 50420
rect 169708 50280 169772 50284
rect 169708 50224 169722 50280
rect 169722 50224 169772 50280
rect 169708 50220 169772 50224
rect 170628 50220 170692 50284
rect 173020 50220 173084 50284
rect 178908 50084 178972 50148
rect 187004 50084 187068 50148
rect 191420 50084 191484 50148
rect 193996 50084 194060 50148
rect 203564 50084 203628 50148
rect 205036 50084 205100 50148
rect 205404 50144 205468 50148
rect 205404 50088 205454 50144
rect 205454 50088 205468 50144
rect 205404 50084 205468 50088
rect 206508 50084 206572 50148
rect 207060 50084 207124 50148
rect 207612 50084 207676 50148
rect 209268 50144 209332 50148
rect 209268 50088 209318 50144
rect 209318 50088 209332 50144
rect 209268 50084 209332 50088
rect 209636 50144 209700 50148
rect 209636 50088 209650 50144
rect 209650 50088 209700 50144
rect 209636 50084 209700 50088
rect 210372 50084 210436 50148
rect 258580 50084 258644 50148
rect 174124 49948 174188 50012
rect 174308 50008 174372 50012
rect 174308 49952 174322 50008
rect 174322 49952 174372 50008
rect 174308 49948 174372 49952
rect 177988 49948 178052 50012
rect 190132 49948 190196 50012
rect 191052 49948 191116 50012
rect 191604 50008 191668 50012
rect 191604 49952 191654 50008
rect 191654 49952 191668 50008
rect 191604 49948 191668 49952
rect 194180 49948 194244 50012
rect 205956 49948 206020 50012
rect 191236 49812 191300 49876
rect 204852 49872 204916 49876
rect 204852 49816 204902 49872
rect 204902 49816 204916 49872
rect 204852 49812 204916 49816
rect 207428 49812 207492 49876
rect 209268 49948 209332 50012
rect 213500 49948 213564 50012
rect 182956 49676 183020 49740
rect 183876 49736 183940 49740
rect 183876 49680 183926 49736
rect 183926 49680 183940 49736
rect 183876 49676 183940 49680
rect 194364 49676 194428 49740
rect 196388 49736 196452 49740
rect 196388 49680 196402 49736
rect 196402 49680 196452 49736
rect 196388 49676 196452 49680
rect 202092 49736 202156 49740
rect 202092 49680 202106 49736
rect 202106 49680 202156 49736
rect 202092 49676 202156 49680
rect 206876 49676 206940 49740
rect 210740 49676 210804 49740
rect 213684 49676 213748 49740
rect 176332 49540 176396 49604
rect 165660 49464 165724 49468
rect 165660 49408 165710 49464
rect 165710 49408 165724 49464
rect 165660 49404 165724 49408
rect 166212 49404 166276 49468
rect 182956 48996 183020 49060
rect 161980 48860 162044 48924
rect 163268 48860 163332 48924
rect 170076 48860 170140 48924
rect 163084 48784 163148 48788
rect 163084 48728 163134 48784
rect 163134 48728 163148 48784
rect 163084 48724 163148 48728
rect 163452 48724 163516 48788
rect 170996 48724 171060 48788
rect 183140 48724 183204 48788
rect 184428 48784 184492 48788
rect 184428 48728 184478 48784
rect 184478 48728 184492 48784
rect 184428 48724 184492 48728
rect 187004 48724 187068 48788
rect 192156 48724 192220 48788
rect 198412 48920 198476 48924
rect 198412 48864 198462 48920
rect 198462 48864 198476 48920
rect 198412 48860 198476 48864
rect 202092 48860 202156 48924
rect 203196 48860 203260 48924
rect 215156 48996 215220 49060
rect 213132 48860 213196 48924
rect 214420 48860 214484 48924
rect 165292 48588 165356 48652
rect 170444 48588 170508 48652
rect 181300 48452 181364 48516
rect 182588 48512 182652 48516
rect 182588 48456 182602 48512
rect 182602 48456 182652 48512
rect 182588 48452 182652 48456
rect 184612 48512 184676 48516
rect 184612 48456 184626 48512
rect 184626 48456 184676 48512
rect 184612 48452 184676 48456
rect 185164 48452 185228 48516
rect 185348 48452 185412 48516
rect 181116 48316 181180 48380
rect 185164 48316 185228 48380
rect 187188 48588 187252 48652
rect 189028 48588 189092 48652
rect 192340 48588 192404 48652
rect 196204 48588 196268 48652
rect 198044 48588 198108 48652
rect 199332 48588 199396 48652
rect 202276 48588 202340 48652
rect 187556 48452 187620 48516
rect 192524 48452 192588 48516
rect 199700 48452 199764 48516
rect 202460 48452 202524 48516
rect 210188 48724 210252 48788
rect 210740 48784 210804 48788
rect 210740 48728 210790 48784
rect 210790 48728 210804 48784
rect 210740 48724 210804 48728
rect 211844 48724 211908 48788
rect 214788 48724 214852 48788
rect 215524 48724 215588 48788
rect 187372 48376 187436 48380
rect 187372 48320 187422 48376
rect 187422 48320 187436 48376
rect 187372 48316 187436 48320
rect 188660 48316 188724 48380
rect 190316 48316 190380 48380
rect 199516 48316 199580 48380
rect 199884 48316 199948 48380
rect 201356 48376 201420 48380
rect 201356 48320 201406 48376
rect 201406 48320 201420 48376
rect 201356 48316 201420 48320
rect 202644 48376 202708 48380
rect 202644 48320 202694 48376
rect 202694 48320 202708 48376
rect 202644 48316 202708 48320
rect 203748 48376 203812 48380
rect 203748 48320 203798 48376
rect 203798 48320 203812 48376
rect 203748 48316 203812 48320
rect 205036 48316 205100 48380
rect 206140 48316 206204 48380
rect 214236 48376 214300 48380
rect 214236 48320 214250 48376
rect 214250 48320 214300 48376
rect 214236 48316 214300 48320
rect 214604 48316 214668 48380
rect 215156 48316 215220 48380
rect 169340 48044 169404 48108
rect 180012 47968 180076 47972
rect 180012 47912 180026 47968
rect 180026 47912 180076 47968
rect 180012 47908 180076 47912
rect 180196 47968 180260 47972
rect 180196 47912 180210 47968
rect 180210 47912 180260 47968
rect 180196 47908 180260 47912
rect 180564 47908 180628 47972
rect 181300 47908 181364 47972
rect 214052 47908 214116 47972
rect 214972 47908 215036 47972
rect 167684 47636 167748 47700
rect 195652 47636 195716 47700
rect 163820 47500 163884 47564
rect 167316 47560 167380 47564
rect 167316 47504 167366 47560
rect 167366 47504 167380 47560
rect 167316 47500 167380 47504
rect 194364 47560 194428 47564
rect 194364 47504 194414 47560
rect 194414 47504 194428 47560
rect 194364 47500 194428 47504
rect 195100 47500 195164 47564
rect 195836 47500 195900 47564
rect 207612 47500 207676 47564
rect 166764 47424 166828 47428
rect 166764 47368 166778 47424
rect 166778 47368 166828 47424
rect 166764 47364 166828 47368
rect 167132 47424 167196 47428
rect 167132 47368 167146 47424
rect 167146 47368 167196 47424
rect 167132 47364 167196 47368
rect 193812 47364 193876 47428
rect 194180 47364 194244 47428
rect 194732 47364 194796 47428
rect 195284 47364 195348 47428
rect 194916 47228 194980 47292
rect 163636 46820 163700 46884
rect 162164 46276 162228 46340
rect 189028 46276 189092 46340
rect 206876 46140 206940 46204
rect 161428 46004 161492 46068
rect 162716 45868 162780 45932
rect 167500 45732 167564 45796
rect 211660 45732 211724 45796
rect 187004 45460 187068 45524
rect 182956 44916 183020 44980
rect 185348 44372 185412 44436
rect 183140 43420 183204 43484
rect 190132 43420 190196 43484
rect 188476 42060 188540 42124
rect 170628 41924 170692 41988
rect 166948 41380 167012 41444
rect 167684 41380 167748 41444
rect 200068 41440 200132 41444
rect 200068 41384 200082 41440
rect 200082 41384 200132 41440
rect 200068 41380 200132 41384
rect 170812 41244 170876 41308
rect 170996 41108 171060 41172
rect 182772 37844 182836 37908
rect 195284 37844 195348 37908
rect 191052 36484 191116 36548
rect 200068 36000 200132 36004
rect 200068 35944 200082 36000
rect 200082 35944 200132 36000
rect 200068 35940 200132 35944
rect 192156 35532 192220 35596
rect 200068 35396 200132 35460
rect 209084 35260 209148 35324
rect 182588 35124 182652 35188
rect 213132 35124 213196 35188
rect 193996 34172 194060 34236
rect 202092 34036 202156 34100
rect 210372 33900 210436 33964
rect 211844 33764 211908 33828
rect 198044 32676 198108 32740
rect 213500 32540 213564 32604
rect 213316 32404 213380 32468
rect 199332 31044 199396 31108
rect 212028 30908 212092 30972
rect 195468 29820 195532 29884
rect 196204 29684 196268 29748
rect 203196 29548 203260 29612
rect 199516 28460 199580 28524
rect 210740 28324 210804 28388
rect 210556 28188 210620 28252
rect 205036 26964 205100 27028
rect 209268 26828 209332 26892
rect 214604 25604 214668 25668
rect 180196 25468 180260 25532
rect 192340 24380 192404 24444
rect 209452 24244 209516 24308
rect 214788 24108 214852 24172
rect 161980 22612 162044 22676
rect 196388 21796 196452 21860
rect 198228 21660 198292 21724
rect 199700 21524 199764 21588
rect 167316 21388 167380 21452
rect 185164 21388 185228 21452
rect 203380 21388 203444 21452
rect 160324 21252 160388 21316
rect 180380 21252 180444 21316
rect 202276 20028 202340 20092
rect 205220 19892 205284 19956
rect 181116 18804 181180 18868
rect 180932 18668 180996 18732
rect 161796 18532 161860 18596
rect 194180 18532 194244 18596
rect 187188 17716 187252 17780
rect 192524 17580 192588 17644
rect 206508 17444 206572 17508
rect 181300 17308 181364 17372
rect 207244 17308 207308 17372
rect 166212 17172 166276 17236
rect 187372 17172 187436 17236
rect 210924 17172 210988 17236
rect 198412 15948 198476 16012
rect 163452 15812 163516 15876
rect 203564 15812 203628 15876
rect 180564 14724 180628 14788
rect 167132 14588 167196 14652
rect 195652 14588 195716 14652
rect 166028 14452 166092 14516
rect 202460 14452 202524 14516
rect 191236 13500 191300 13564
rect 191420 13364 191484 13428
rect 192708 13228 192772 13292
rect 166948 13092 167012 13156
rect 195836 13092 195900 13156
rect 165844 12956 165908 13020
rect 201356 12956 201420 13020
rect 206692 12004 206756 12068
rect 212212 11868 212276 11932
rect 212396 11732 212460 11796
rect 160140 11596 160204 11660
rect 214972 11596 215036 11660
rect 163268 10236 163332 10300
rect 209636 10236 209700 10300
rect 169156 9148 169220 9212
rect 169340 9012 169404 9076
rect 205404 9012 205468 9076
rect 161612 8876 161676 8940
rect 213684 8876 213748 8940
rect 190316 6836 190380 6900
rect 194364 6700 194428 6764
rect 198596 6564 198660 6628
rect 199884 6428 199948 6492
rect 163084 6292 163148 6356
rect 202644 6292 202708 6356
rect 162900 6156 162964 6220
rect 183692 6156 183756 6220
rect 207428 6156 207492 6220
rect 188660 6020 188724 6084
rect 168972 5068 169036 5132
rect 165660 4932 165724 4996
rect 203748 4932 203812 4996
rect 165292 4796 165356 4860
rect 183876 4796 183940 4860
rect 187556 4796 187620 4860
rect 214420 4796 214484 4860
rect 191604 3708 191668 3772
rect 188844 3572 188908 3636
rect 258580 3436 258644 3500
rect 206324 3300 206388 3364
<< metal4 >>
rect -8726 711558 -8106 711590
rect -8726 711322 -8694 711558
rect -8458 711322 -8374 711558
rect -8138 711322 -8106 711558
rect -8726 711238 -8106 711322
rect -8726 711002 -8694 711238
rect -8458 711002 -8374 711238
rect -8138 711002 -8106 711238
rect -8726 677494 -8106 711002
rect -8726 677258 -8694 677494
rect -8458 677258 -8374 677494
rect -8138 677258 -8106 677494
rect -8726 677174 -8106 677258
rect -8726 676938 -8694 677174
rect -8458 676938 -8374 677174
rect -8138 676938 -8106 677174
rect -8726 641494 -8106 676938
rect -8726 641258 -8694 641494
rect -8458 641258 -8374 641494
rect -8138 641258 -8106 641494
rect -8726 641174 -8106 641258
rect -8726 640938 -8694 641174
rect -8458 640938 -8374 641174
rect -8138 640938 -8106 641174
rect -8726 605494 -8106 640938
rect -8726 605258 -8694 605494
rect -8458 605258 -8374 605494
rect -8138 605258 -8106 605494
rect -8726 605174 -8106 605258
rect -8726 604938 -8694 605174
rect -8458 604938 -8374 605174
rect -8138 604938 -8106 605174
rect -8726 569494 -8106 604938
rect -8726 569258 -8694 569494
rect -8458 569258 -8374 569494
rect -8138 569258 -8106 569494
rect -8726 569174 -8106 569258
rect -8726 568938 -8694 569174
rect -8458 568938 -8374 569174
rect -8138 568938 -8106 569174
rect -8726 533494 -8106 568938
rect -8726 533258 -8694 533494
rect -8458 533258 -8374 533494
rect -8138 533258 -8106 533494
rect -8726 533174 -8106 533258
rect -8726 532938 -8694 533174
rect -8458 532938 -8374 533174
rect -8138 532938 -8106 533174
rect -8726 497494 -8106 532938
rect -8726 497258 -8694 497494
rect -8458 497258 -8374 497494
rect -8138 497258 -8106 497494
rect -8726 497174 -8106 497258
rect -8726 496938 -8694 497174
rect -8458 496938 -8374 497174
rect -8138 496938 -8106 497174
rect -8726 461494 -8106 496938
rect -8726 461258 -8694 461494
rect -8458 461258 -8374 461494
rect -8138 461258 -8106 461494
rect -8726 461174 -8106 461258
rect -8726 460938 -8694 461174
rect -8458 460938 -8374 461174
rect -8138 460938 -8106 461174
rect -8726 425494 -8106 460938
rect -8726 425258 -8694 425494
rect -8458 425258 -8374 425494
rect -8138 425258 -8106 425494
rect -8726 425174 -8106 425258
rect -8726 424938 -8694 425174
rect -8458 424938 -8374 425174
rect -8138 424938 -8106 425174
rect -8726 389494 -8106 424938
rect -8726 389258 -8694 389494
rect -8458 389258 -8374 389494
rect -8138 389258 -8106 389494
rect -8726 389174 -8106 389258
rect -8726 388938 -8694 389174
rect -8458 388938 -8374 389174
rect -8138 388938 -8106 389174
rect -8726 353494 -8106 388938
rect -8726 353258 -8694 353494
rect -8458 353258 -8374 353494
rect -8138 353258 -8106 353494
rect -8726 353174 -8106 353258
rect -8726 352938 -8694 353174
rect -8458 352938 -8374 353174
rect -8138 352938 -8106 353174
rect -8726 317494 -8106 352938
rect -8726 317258 -8694 317494
rect -8458 317258 -8374 317494
rect -8138 317258 -8106 317494
rect -8726 317174 -8106 317258
rect -8726 316938 -8694 317174
rect -8458 316938 -8374 317174
rect -8138 316938 -8106 317174
rect -8726 281494 -8106 316938
rect -8726 281258 -8694 281494
rect -8458 281258 -8374 281494
rect -8138 281258 -8106 281494
rect -8726 281174 -8106 281258
rect -8726 280938 -8694 281174
rect -8458 280938 -8374 281174
rect -8138 280938 -8106 281174
rect -8726 245494 -8106 280938
rect -8726 245258 -8694 245494
rect -8458 245258 -8374 245494
rect -8138 245258 -8106 245494
rect -8726 245174 -8106 245258
rect -8726 244938 -8694 245174
rect -8458 244938 -8374 245174
rect -8138 244938 -8106 245174
rect -8726 209494 -8106 244938
rect -8726 209258 -8694 209494
rect -8458 209258 -8374 209494
rect -8138 209258 -8106 209494
rect -8726 209174 -8106 209258
rect -8726 208938 -8694 209174
rect -8458 208938 -8374 209174
rect -8138 208938 -8106 209174
rect -8726 173494 -8106 208938
rect -8726 173258 -8694 173494
rect -8458 173258 -8374 173494
rect -8138 173258 -8106 173494
rect -8726 173174 -8106 173258
rect -8726 172938 -8694 173174
rect -8458 172938 -8374 173174
rect -8138 172938 -8106 173174
rect -8726 137494 -8106 172938
rect -8726 137258 -8694 137494
rect -8458 137258 -8374 137494
rect -8138 137258 -8106 137494
rect -8726 137174 -8106 137258
rect -8726 136938 -8694 137174
rect -8458 136938 -8374 137174
rect -8138 136938 -8106 137174
rect -8726 101494 -8106 136938
rect -8726 101258 -8694 101494
rect -8458 101258 -8374 101494
rect -8138 101258 -8106 101494
rect -8726 101174 -8106 101258
rect -8726 100938 -8694 101174
rect -8458 100938 -8374 101174
rect -8138 100938 -8106 101174
rect -8726 65494 -8106 100938
rect -8726 65258 -8694 65494
rect -8458 65258 -8374 65494
rect -8138 65258 -8106 65494
rect -8726 65174 -8106 65258
rect -8726 64938 -8694 65174
rect -8458 64938 -8374 65174
rect -8138 64938 -8106 65174
rect -8726 29494 -8106 64938
rect -8726 29258 -8694 29494
rect -8458 29258 -8374 29494
rect -8138 29258 -8106 29494
rect -8726 29174 -8106 29258
rect -8726 28938 -8694 29174
rect -8458 28938 -8374 29174
rect -8138 28938 -8106 29174
rect -8726 -7066 -8106 28938
rect -7766 710598 -7146 710630
rect -7766 710362 -7734 710598
rect -7498 710362 -7414 710598
rect -7178 710362 -7146 710598
rect -7766 710278 -7146 710362
rect -7766 710042 -7734 710278
rect -7498 710042 -7414 710278
rect -7178 710042 -7146 710278
rect -7766 673774 -7146 710042
rect -7766 673538 -7734 673774
rect -7498 673538 -7414 673774
rect -7178 673538 -7146 673774
rect -7766 673454 -7146 673538
rect -7766 673218 -7734 673454
rect -7498 673218 -7414 673454
rect -7178 673218 -7146 673454
rect -7766 637774 -7146 673218
rect -7766 637538 -7734 637774
rect -7498 637538 -7414 637774
rect -7178 637538 -7146 637774
rect -7766 637454 -7146 637538
rect -7766 637218 -7734 637454
rect -7498 637218 -7414 637454
rect -7178 637218 -7146 637454
rect -7766 601774 -7146 637218
rect -7766 601538 -7734 601774
rect -7498 601538 -7414 601774
rect -7178 601538 -7146 601774
rect -7766 601454 -7146 601538
rect -7766 601218 -7734 601454
rect -7498 601218 -7414 601454
rect -7178 601218 -7146 601454
rect -7766 565774 -7146 601218
rect -7766 565538 -7734 565774
rect -7498 565538 -7414 565774
rect -7178 565538 -7146 565774
rect -7766 565454 -7146 565538
rect -7766 565218 -7734 565454
rect -7498 565218 -7414 565454
rect -7178 565218 -7146 565454
rect -7766 529774 -7146 565218
rect -7766 529538 -7734 529774
rect -7498 529538 -7414 529774
rect -7178 529538 -7146 529774
rect -7766 529454 -7146 529538
rect -7766 529218 -7734 529454
rect -7498 529218 -7414 529454
rect -7178 529218 -7146 529454
rect -7766 493774 -7146 529218
rect -7766 493538 -7734 493774
rect -7498 493538 -7414 493774
rect -7178 493538 -7146 493774
rect -7766 493454 -7146 493538
rect -7766 493218 -7734 493454
rect -7498 493218 -7414 493454
rect -7178 493218 -7146 493454
rect -7766 457774 -7146 493218
rect -7766 457538 -7734 457774
rect -7498 457538 -7414 457774
rect -7178 457538 -7146 457774
rect -7766 457454 -7146 457538
rect -7766 457218 -7734 457454
rect -7498 457218 -7414 457454
rect -7178 457218 -7146 457454
rect -7766 421774 -7146 457218
rect -7766 421538 -7734 421774
rect -7498 421538 -7414 421774
rect -7178 421538 -7146 421774
rect -7766 421454 -7146 421538
rect -7766 421218 -7734 421454
rect -7498 421218 -7414 421454
rect -7178 421218 -7146 421454
rect -7766 385774 -7146 421218
rect -7766 385538 -7734 385774
rect -7498 385538 -7414 385774
rect -7178 385538 -7146 385774
rect -7766 385454 -7146 385538
rect -7766 385218 -7734 385454
rect -7498 385218 -7414 385454
rect -7178 385218 -7146 385454
rect -7766 349774 -7146 385218
rect -7766 349538 -7734 349774
rect -7498 349538 -7414 349774
rect -7178 349538 -7146 349774
rect -7766 349454 -7146 349538
rect -7766 349218 -7734 349454
rect -7498 349218 -7414 349454
rect -7178 349218 -7146 349454
rect -7766 313774 -7146 349218
rect -7766 313538 -7734 313774
rect -7498 313538 -7414 313774
rect -7178 313538 -7146 313774
rect -7766 313454 -7146 313538
rect -7766 313218 -7734 313454
rect -7498 313218 -7414 313454
rect -7178 313218 -7146 313454
rect -7766 277774 -7146 313218
rect -7766 277538 -7734 277774
rect -7498 277538 -7414 277774
rect -7178 277538 -7146 277774
rect -7766 277454 -7146 277538
rect -7766 277218 -7734 277454
rect -7498 277218 -7414 277454
rect -7178 277218 -7146 277454
rect -7766 241774 -7146 277218
rect -7766 241538 -7734 241774
rect -7498 241538 -7414 241774
rect -7178 241538 -7146 241774
rect -7766 241454 -7146 241538
rect -7766 241218 -7734 241454
rect -7498 241218 -7414 241454
rect -7178 241218 -7146 241454
rect -7766 205774 -7146 241218
rect -7766 205538 -7734 205774
rect -7498 205538 -7414 205774
rect -7178 205538 -7146 205774
rect -7766 205454 -7146 205538
rect -7766 205218 -7734 205454
rect -7498 205218 -7414 205454
rect -7178 205218 -7146 205454
rect -7766 169774 -7146 205218
rect -7766 169538 -7734 169774
rect -7498 169538 -7414 169774
rect -7178 169538 -7146 169774
rect -7766 169454 -7146 169538
rect -7766 169218 -7734 169454
rect -7498 169218 -7414 169454
rect -7178 169218 -7146 169454
rect -7766 133774 -7146 169218
rect -7766 133538 -7734 133774
rect -7498 133538 -7414 133774
rect -7178 133538 -7146 133774
rect -7766 133454 -7146 133538
rect -7766 133218 -7734 133454
rect -7498 133218 -7414 133454
rect -7178 133218 -7146 133454
rect -7766 97774 -7146 133218
rect -7766 97538 -7734 97774
rect -7498 97538 -7414 97774
rect -7178 97538 -7146 97774
rect -7766 97454 -7146 97538
rect -7766 97218 -7734 97454
rect -7498 97218 -7414 97454
rect -7178 97218 -7146 97454
rect -7766 61774 -7146 97218
rect -7766 61538 -7734 61774
rect -7498 61538 -7414 61774
rect -7178 61538 -7146 61774
rect -7766 61454 -7146 61538
rect -7766 61218 -7734 61454
rect -7498 61218 -7414 61454
rect -7178 61218 -7146 61454
rect -7766 25774 -7146 61218
rect -7766 25538 -7734 25774
rect -7498 25538 -7414 25774
rect -7178 25538 -7146 25774
rect -7766 25454 -7146 25538
rect -7766 25218 -7734 25454
rect -7498 25218 -7414 25454
rect -7178 25218 -7146 25454
rect -7766 -6106 -7146 25218
rect -6806 709638 -6186 709670
rect -6806 709402 -6774 709638
rect -6538 709402 -6454 709638
rect -6218 709402 -6186 709638
rect -6806 709318 -6186 709402
rect -6806 709082 -6774 709318
rect -6538 709082 -6454 709318
rect -6218 709082 -6186 709318
rect -6806 670054 -6186 709082
rect -6806 669818 -6774 670054
rect -6538 669818 -6454 670054
rect -6218 669818 -6186 670054
rect -6806 669734 -6186 669818
rect -6806 669498 -6774 669734
rect -6538 669498 -6454 669734
rect -6218 669498 -6186 669734
rect -6806 634054 -6186 669498
rect -6806 633818 -6774 634054
rect -6538 633818 -6454 634054
rect -6218 633818 -6186 634054
rect -6806 633734 -6186 633818
rect -6806 633498 -6774 633734
rect -6538 633498 -6454 633734
rect -6218 633498 -6186 633734
rect -6806 598054 -6186 633498
rect -6806 597818 -6774 598054
rect -6538 597818 -6454 598054
rect -6218 597818 -6186 598054
rect -6806 597734 -6186 597818
rect -6806 597498 -6774 597734
rect -6538 597498 -6454 597734
rect -6218 597498 -6186 597734
rect -6806 562054 -6186 597498
rect -6806 561818 -6774 562054
rect -6538 561818 -6454 562054
rect -6218 561818 -6186 562054
rect -6806 561734 -6186 561818
rect -6806 561498 -6774 561734
rect -6538 561498 -6454 561734
rect -6218 561498 -6186 561734
rect -6806 526054 -6186 561498
rect -6806 525818 -6774 526054
rect -6538 525818 -6454 526054
rect -6218 525818 -6186 526054
rect -6806 525734 -6186 525818
rect -6806 525498 -6774 525734
rect -6538 525498 -6454 525734
rect -6218 525498 -6186 525734
rect -6806 490054 -6186 525498
rect -6806 489818 -6774 490054
rect -6538 489818 -6454 490054
rect -6218 489818 -6186 490054
rect -6806 489734 -6186 489818
rect -6806 489498 -6774 489734
rect -6538 489498 -6454 489734
rect -6218 489498 -6186 489734
rect -6806 454054 -6186 489498
rect -6806 453818 -6774 454054
rect -6538 453818 -6454 454054
rect -6218 453818 -6186 454054
rect -6806 453734 -6186 453818
rect -6806 453498 -6774 453734
rect -6538 453498 -6454 453734
rect -6218 453498 -6186 453734
rect -6806 418054 -6186 453498
rect -6806 417818 -6774 418054
rect -6538 417818 -6454 418054
rect -6218 417818 -6186 418054
rect -6806 417734 -6186 417818
rect -6806 417498 -6774 417734
rect -6538 417498 -6454 417734
rect -6218 417498 -6186 417734
rect -6806 382054 -6186 417498
rect -6806 381818 -6774 382054
rect -6538 381818 -6454 382054
rect -6218 381818 -6186 382054
rect -6806 381734 -6186 381818
rect -6806 381498 -6774 381734
rect -6538 381498 -6454 381734
rect -6218 381498 -6186 381734
rect -6806 346054 -6186 381498
rect -6806 345818 -6774 346054
rect -6538 345818 -6454 346054
rect -6218 345818 -6186 346054
rect -6806 345734 -6186 345818
rect -6806 345498 -6774 345734
rect -6538 345498 -6454 345734
rect -6218 345498 -6186 345734
rect -6806 310054 -6186 345498
rect -6806 309818 -6774 310054
rect -6538 309818 -6454 310054
rect -6218 309818 -6186 310054
rect -6806 309734 -6186 309818
rect -6806 309498 -6774 309734
rect -6538 309498 -6454 309734
rect -6218 309498 -6186 309734
rect -6806 274054 -6186 309498
rect -6806 273818 -6774 274054
rect -6538 273818 -6454 274054
rect -6218 273818 -6186 274054
rect -6806 273734 -6186 273818
rect -6806 273498 -6774 273734
rect -6538 273498 -6454 273734
rect -6218 273498 -6186 273734
rect -6806 238054 -6186 273498
rect -6806 237818 -6774 238054
rect -6538 237818 -6454 238054
rect -6218 237818 -6186 238054
rect -6806 237734 -6186 237818
rect -6806 237498 -6774 237734
rect -6538 237498 -6454 237734
rect -6218 237498 -6186 237734
rect -6806 202054 -6186 237498
rect -6806 201818 -6774 202054
rect -6538 201818 -6454 202054
rect -6218 201818 -6186 202054
rect -6806 201734 -6186 201818
rect -6806 201498 -6774 201734
rect -6538 201498 -6454 201734
rect -6218 201498 -6186 201734
rect -6806 166054 -6186 201498
rect -6806 165818 -6774 166054
rect -6538 165818 -6454 166054
rect -6218 165818 -6186 166054
rect -6806 165734 -6186 165818
rect -6806 165498 -6774 165734
rect -6538 165498 -6454 165734
rect -6218 165498 -6186 165734
rect -6806 130054 -6186 165498
rect -6806 129818 -6774 130054
rect -6538 129818 -6454 130054
rect -6218 129818 -6186 130054
rect -6806 129734 -6186 129818
rect -6806 129498 -6774 129734
rect -6538 129498 -6454 129734
rect -6218 129498 -6186 129734
rect -6806 94054 -6186 129498
rect -6806 93818 -6774 94054
rect -6538 93818 -6454 94054
rect -6218 93818 -6186 94054
rect -6806 93734 -6186 93818
rect -6806 93498 -6774 93734
rect -6538 93498 -6454 93734
rect -6218 93498 -6186 93734
rect -6806 58054 -6186 93498
rect -6806 57818 -6774 58054
rect -6538 57818 -6454 58054
rect -6218 57818 -6186 58054
rect -6806 57734 -6186 57818
rect -6806 57498 -6774 57734
rect -6538 57498 -6454 57734
rect -6218 57498 -6186 57734
rect -6806 22054 -6186 57498
rect -6806 21818 -6774 22054
rect -6538 21818 -6454 22054
rect -6218 21818 -6186 22054
rect -6806 21734 -6186 21818
rect -6806 21498 -6774 21734
rect -6538 21498 -6454 21734
rect -6218 21498 -6186 21734
rect -6806 -5146 -6186 21498
rect -5846 708678 -5226 708710
rect -5846 708442 -5814 708678
rect -5578 708442 -5494 708678
rect -5258 708442 -5226 708678
rect -5846 708358 -5226 708442
rect -5846 708122 -5814 708358
rect -5578 708122 -5494 708358
rect -5258 708122 -5226 708358
rect -5846 666334 -5226 708122
rect -5846 666098 -5814 666334
rect -5578 666098 -5494 666334
rect -5258 666098 -5226 666334
rect -5846 666014 -5226 666098
rect -5846 665778 -5814 666014
rect -5578 665778 -5494 666014
rect -5258 665778 -5226 666014
rect -5846 630334 -5226 665778
rect -5846 630098 -5814 630334
rect -5578 630098 -5494 630334
rect -5258 630098 -5226 630334
rect -5846 630014 -5226 630098
rect -5846 629778 -5814 630014
rect -5578 629778 -5494 630014
rect -5258 629778 -5226 630014
rect -5846 594334 -5226 629778
rect -5846 594098 -5814 594334
rect -5578 594098 -5494 594334
rect -5258 594098 -5226 594334
rect -5846 594014 -5226 594098
rect -5846 593778 -5814 594014
rect -5578 593778 -5494 594014
rect -5258 593778 -5226 594014
rect -5846 558334 -5226 593778
rect -5846 558098 -5814 558334
rect -5578 558098 -5494 558334
rect -5258 558098 -5226 558334
rect -5846 558014 -5226 558098
rect -5846 557778 -5814 558014
rect -5578 557778 -5494 558014
rect -5258 557778 -5226 558014
rect -5846 522334 -5226 557778
rect -5846 522098 -5814 522334
rect -5578 522098 -5494 522334
rect -5258 522098 -5226 522334
rect -5846 522014 -5226 522098
rect -5846 521778 -5814 522014
rect -5578 521778 -5494 522014
rect -5258 521778 -5226 522014
rect -5846 486334 -5226 521778
rect -5846 486098 -5814 486334
rect -5578 486098 -5494 486334
rect -5258 486098 -5226 486334
rect -5846 486014 -5226 486098
rect -5846 485778 -5814 486014
rect -5578 485778 -5494 486014
rect -5258 485778 -5226 486014
rect -5846 450334 -5226 485778
rect -5846 450098 -5814 450334
rect -5578 450098 -5494 450334
rect -5258 450098 -5226 450334
rect -5846 450014 -5226 450098
rect -5846 449778 -5814 450014
rect -5578 449778 -5494 450014
rect -5258 449778 -5226 450014
rect -5846 414334 -5226 449778
rect -5846 414098 -5814 414334
rect -5578 414098 -5494 414334
rect -5258 414098 -5226 414334
rect -5846 414014 -5226 414098
rect -5846 413778 -5814 414014
rect -5578 413778 -5494 414014
rect -5258 413778 -5226 414014
rect -5846 378334 -5226 413778
rect -5846 378098 -5814 378334
rect -5578 378098 -5494 378334
rect -5258 378098 -5226 378334
rect -5846 378014 -5226 378098
rect -5846 377778 -5814 378014
rect -5578 377778 -5494 378014
rect -5258 377778 -5226 378014
rect -5846 342334 -5226 377778
rect -5846 342098 -5814 342334
rect -5578 342098 -5494 342334
rect -5258 342098 -5226 342334
rect -5846 342014 -5226 342098
rect -5846 341778 -5814 342014
rect -5578 341778 -5494 342014
rect -5258 341778 -5226 342014
rect -5846 306334 -5226 341778
rect -5846 306098 -5814 306334
rect -5578 306098 -5494 306334
rect -5258 306098 -5226 306334
rect -5846 306014 -5226 306098
rect -5846 305778 -5814 306014
rect -5578 305778 -5494 306014
rect -5258 305778 -5226 306014
rect -5846 270334 -5226 305778
rect -5846 270098 -5814 270334
rect -5578 270098 -5494 270334
rect -5258 270098 -5226 270334
rect -5846 270014 -5226 270098
rect -5846 269778 -5814 270014
rect -5578 269778 -5494 270014
rect -5258 269778 -5226 270014
rect -5846 234334 -5226 269778
rect -5846 234098 -5814 234334
rect -5578 234098 -5494 234334
rect -5258 234098 -5226 234334
rect -5846 234014 -5226 234098
rect -5846 233778 -5814 234014
rect -5578 233778 -5494 234014
rect -5258 233778 -5226 234014
rect -5846 198334 -5226 233778
rect -5846 198098 -5814 198334
rect -5578 198098 -5494 198334
rect -5258 198098 -5226 198334
rect -5846 198014 -5226 198098
rect -5846 197778 -5814 198014
rect -5578 197778 -5494 198014
rect -5258 197778 -5226 198014
rect -5846 162334 -5226 197778
rect -5846 162098 -5814 162334
rect -5578 162098 -5494 162334
rect -5258 162098 -5226 162334
rect -5846 162014 -5226 162098
rect -5846 161778 -5814 162014
rect -5578 161778 -5494 162014
rect -5258 161778 -5226 162014
rect -5846 126334 -5226 161778
rect -5846 126098 -5814 126334
rect -5578 126098 -5494 126334
rect -5258 126098 -5226 126334
rect -5846 126014 -5226 126098
rect -5846 125778 -5814 126014
rect -5578 125778 -5494 126014
rect -5258 125778 -5226 126014
rect -5846 90334 -5226 125778
rect -5846 90098 -5814 90334
rect -5578 90098 -5494 90334
rect -5258 90098 -5226 90334
rect -5846 90014 -5226 90098
rect -5846 89778 -5814 90014
rect -5578 89778 -5494 90014
rect -5258 89778 -5226 90014
rect -5846 54334 -5226 89778
rect -5846 54098 -5814 54334
rect -5578 54098 -5494 54334
rect -5258 54098 -5226 54334
rect -5846 54014 -5226 54098
rect -5846 53778 -5814 54014
rect -5578 53778 -5494 54014
rect -5258 53778 -5226 54014
rect -5846 18334 -5226 53778
rect -5846 18098 -5814 18334
rect -5578 18098 -5494 18334
rect -5258 18098 -5226 18334
rect -5846 18014 -5226 18098
rect -5846 17778 -5814 18014
rect -5578 17778 -5494 18014
rect -5258 17778 -5226 18014
rect -5846 -4186 -5226 17778
rect -4886 707718 -4266 707750
rect -4886 707482 -4854 707718
rect -4618 707482 -4534 707718
rect -4298 707482 -4266 707718
rect -4886 707398 -4266 707482
rect -4886 707162 -4854 707398
rect -4618 707162 -4534 707398
rect -4298 707162 -4266 707398
rect -4886 698614 -4266 707162
rect -4886 698378 -4854 698614
rect -4618 698378 -4534 698614
rect -4298 698378 -4266 698614
rect -4886 698294 -4266 698378
rect -4886 698058 -4854 698294
rect -4618 698058 -4534 698294
rect -4298 698058 -4266 698294
rect -4886 662614 -4266 698058
rect -4886 662378 -4854 662614
rect -4618 662378 -4534 662614
rect -4298 662378 -4266 662614
rect -4886 662294 -4266 662378
rect -4886 662058 -4854 662294
rect -4618 662058 -4534 662294
rect -4298 662058 -4266 662294
rect -4886 626614 -4266 662058
rect -4886 626378 -4854 626614
rect -4618 626378 -4534 626614
rect -4298 626378 -4266 626614
rect -4886 626294 -4266 626378
rect -4886 626058 -4854 626294
rect -4618 626058 -4534 626294
rect -4298 626058 -4266 626294
rect -4886 590614 -4266 626058
rect -4886 590378 -4854 590614
rect -4618 590378 -4534 590614
rect -4298 590378 -4266 590614
rect -4886 590294 -4266 590378
rect -4886 590058 -4854 590294
rect -4618 590058 -4534 590294
rect -4298 590058 -4266 590294
rect -4886 554614 -4266 590058
rect -4886 554378 -4854 554614
rect -4618 554378 -4534 554614
rect -4298 554378 -4266 554614
rect -4886 554294 -4266 554378
rect -4886 554058 -4854 554294
rect -4618 554058 -4534 554294
rect -4298 554058 -4266 554294
rect -4886 518614 -4266 554058
rect -4886 518378 -4854 518614
rect -4618 518378 -4534 518614
rect -4298 518378 -4266 518614
rect -4886 518294 -4266 518378
rect -4886 518058 -4854 518294
rect -4618 518058 -4534 518294
rect -4298 518058 -4266 518294
rect -4886 482614 -4266 518058
rect -4886 482378 -4854 482614
rect -4618 482378 -4534 482614
rect -4298 482378 -4266 482614
rect -4886 482294 -4266 482378
rect -4886 482058 -4854 482294
rect -4618 482058 -4534 482294
rect -4298 482058 -4266 482294
rect -4886 446614 -4266 482058
rect -4886 446378 -4854 446614
rect -4618 446378 -4534 446614
rect -4298 446378 -4266 446614
rect -4886 446294 -4266 446378
rect -4886 446058 -4854 446294
rect -4618 446058 -4534 446294
rect -4298 446058 -4266 446294
rect -4886 410614 -4266 446058
rect -4886 410378 -4854 410614
rect -4618 410378 -4534 410614
rect -4298 410378 -4266 410614
rect -4886 410294 -4266 410378
rect -4886 410058 -4854 410294
rect -4618 410058 -4534 410294
rect -4298 410058 -4266 410294
rect -4886 374614 -4266 410058
rect -4886 374378 -4854 374614
rect -4618 374378 -4534 374614
rect -4298 374378 -4266 374614
rect -4886 374294 -4266 374378
rect -4886 374058 -4854 374294
rect -4618 374058 -4534 374294
rect -4298 374058 -4266 374294
rect -4886 338614 -4266 374058
rect -4886 338378 -4854 338614
rect -4618 338378 -4534 338614
rect -4298 338378 -4266 338614
rect -4886 338294 -4266 338378
rect -4886 338058 -4854 338294
rect -4618 338058 -4534 338294
rect -4298 338058 -4266 338294
rect -4886 302614 -4266 338058
rect -4886 302378 -4854 302614
rect -4618 302378 -4534 302614
rect -4298 302378 -4266 302614
rect -4886 302294 -4266 302378
rect -4886 302058 -4854 302294
rect -4618 302058 -4534 302294
rect -4298 302058 -4266 302294
rect -4886 266614 -4266 302058
rect -4886 266378 -4854 266614
rect -4618 266378 -4534 266614
rect -4298 266378 -4266 266614
rect -4886 266294 -4266 266378
rect -4886 266058 -4854 266294
rect -4618 266058 -4534 266294
rect -4298 266058 -4266 266294
rect -4886 230614 -4266 266058
rect -4886 230378 -4854 230614
rect -4618 230378 -4534 230614
rect -4298 230378 -4266 230614
rect -4886 230294 -4266 230378
rect -4886 230058 -4854 230294
rect -4618 230058 -4534 230294
rect -4298 230058 -4266 230294
rect -4886 194614 -4266 230058
rect -4886 194378 -4854 194614
rect -4618 194378 -4534 194614
rect -4298 194378 -4266 194614
rect -4886 194294 -4266 194378
rect -4886 194058 -4854 194294
rect -4618 194058 -4534 194294
rect -4298 194058 -4266 194294
rect -4886 158614 -4266 194058
rect -4886 158378 -4854 158614
rect -4618 158378 -4534 158614
rect -4298 158378 -4266 158614
rect -4886 158294 -4266 158378
rect -4886 158058 -4854 158294
rect -4618 158058 -4534 158294
rect -4298 158058 -4266 158294
rect -4886 122614 -4266 158058
rect -4886 122378 -4854 122614
rect -4618 122378 -4534 122614
rect -4298 122378 -4266 122614
rect -4886 122294 -4266 122378
rect -4886 122058 -4854 122294
rect -4618 122058 -4534 122294
rect -4298 122058 -4266 122294
rect -4886 86614 -4266 122058
rect -4886 86378 -4854 86614
rect -4618 86378 -4534 86614
rect -4298 86378 -4266 86614
rect -4886 86294 -4266 86378
rect -4886 86058 -4854 86294
rect -4618 86058 -4534 86294
rect -4298 86058 -4266 86294
rect -4886 50614 -4266 86058
rect -4886 50378 -4854 50614
rect -4618 50378 -4534 50614
rect -4298 50378 -4266 50614
rect -4886 50294 -4266 50378
rect -4886 50058 -4854 50294
rect -4618 50058 -4534 50294
rect -4298 50058 -4266 50294
rect -4886 14614 -4266 50058
rect -4886 14378 -4854 14614
rect -4618 14378 -4534 14614
rect -4298 14378 -4266 14614
rect -4886 14294 -4266 14378
rect -4886 14058 -4854 14294
rect -4618 14058 -4534 14294
rect -4298 14058 -4266 14294
rect -4886 -3226 -4266 14058
rect -3926 706758 -3306 706790
rect -3926 706522 -3894 706758
rect -3658 706522 -3574 706758
rect -3338 706522 -3306 706758
rect -3926 706438 -3306 706522
rect -3926 706202 -3894 706438
rect -3658 706202 -3574 706438
rect -3338 706202 -3306 706438
rect -3926 694894 -3306 706202
rect -3926 694658 -3894 694894
rect -3658 694658 -3574 694894
rect -3338 694658 -3306 694894
rect -3926 694574 -3306 694658
rect -3926 694338 -3894 694574
rect -3658 694338 -3574 694574
rect -3338 694338 -3306 694574
rect -3926 658894 -3306 694338
rect -3926 658658 -3894 658894
rect -3658 658658 -3574 658894
rect -3338 658658 -3306 658894
rect -3926 658574 -3306 658658
rect -3926 658338 -3894 658574
rect -3658 658338 -3574 658574
rect -3338 658338 -3306 658574
rect -3926 622894 -3306 658338
rect -3926 622658 -3894 622894
rect -3658 622658 -3574 622894
rect -3338 622658 -3306 622894
rect -3926 622574 -3306 622658
rect -3926 622338 -3894 622574
rect -3658 622338 -3574 622574
rect -3338 622338 -3306 622574
rect -3926 586894 -3306 622338
rect -3926 586658 -3894 586894
rect -3658 586658 -3574 586894
rect -3338 586658 -3306 586894
rect -3926 586574 -3306 586658
rect -3926 586338 -3894 586574
rect -3658 586338 -3574 586574
rect -3338 586338 -3306 586574
rect -3926 550894 -3306 586338
rect -3926 550658 -3894 550894
rect -3658 550658 -3574 550894
rect -3338 550658 -3306 550894
rect -3926 550574 -3306 550658
rect -3926 550338 -3894 550574
rect -3658 550338 -3574 550574
rect -3338 550338 -3306 550574
rect -3926 514894 -3306 550338
rect -3926 514658 -3894 514894
rect -3658 514658 -3574 514894
rect -3338 514658 -3306 514894
rect -3926 514574 -3306 514658
rect -3926 514338 -3894 514574
rect -3658 514338 -3574 514574
rect -3338 514338 -3306 514574
rect -3926 478894 -3306 514338
rect -3926 478658 -3894 478894
rect -3658 478658 -3574 478894
rect -3338 478658 -3306 478894
rect -3926 478574 -3306 478658
rect -3926 478338 -3894 478574
rect -3658 478338 -3574 478574
rect -3338 478338 -3306 478574
rect -3926 442894 -3306 478338
rect -3926 442658 -3894 442894
rect -3658 442658 -3574 442894
rect -3338 442658 -3306 442894
rect -3926 442574 -3306 442658
rect -3926 442338 -3894 442574
rect -3658 442338 -3574 442574
rect -3338 442338 -3306 442574
rect -3926 406894 -3306 442338
rect -3926 406658 -3894 406894
rect -3658 406658 -3574 406894
rect -3338 406658 -3306 406894
rect -3926 406574 -3306 406658
rect -3926 406338 -3894 406574
rect -3658 406338 -3574 406574
rect -3338 406338 -3306 406574
rect -3926 370894 -3306 406338
rect -3926 370658 -3894 370894
rect -3658 370658 -3574 370894
rect -3338 370658 -3306 370894
rect -3926 370574 -3306 370658
rect -3926 370338 -3894 370574
rect -3658 370338 -3574 370574
rect -3338 370338 -3306 370574
rect -3926 334894 -3306 370338
rect -3926 334658 -3894 334894
rect -3658 334658 -3574 334894
rect -3338 334658 -3306 334894
rect -3926 334574 -3306 334658
rect -3926 334338 -3894 334574
rect -3658 334338 -3574 334574
rect -3338 334338 -3306 334574
rect -3926 298894 -3306 334338
rect -3926 298658 -3894 298894
rect -3658 298658 -3574 298894
rect -3338 298658 -3306 298894
rect -3926 298574 -3306 298658
rect -3926 298338 -3894 298574
rect -3658 298338 -3574 298574
rect -3338 298338 -3306 298574
rect -3926 262894 -3306 298338
rect -3926 262658 -3894 262894
rect -3658 262658 -3574 262894
rect -3338 262658 -3306 262894
rect -3926 262574 -3306 262658
rect -3926 262338 -3894 262574
rect -3658 262338 -3574 262574
rect -3338 262338 -3306 262574
rect -3926 226894 -3306 262338
rect -3926 226658 -3894 226894
rect -3658 226658 -3574 226894
rect -3338 226658 -3306 226894
rect -3926 226574 -3306 226658
rect -3926 226338 -3894 226574
rect -3658 226338 -3574 226574
rect -3338 226338 -3306 226574
rect -3926 190894 -3306 226338
rect -3926 190658 -3894 190894
rect -3658 190658 -3574 190894
rect -3338 190658 -3306 190894
rect -3926 190574 -3306 190658
rect -3926 190338 -3894 190574
rect -3658 190338 -3574 190574
rect -3338 190338 -3306 190574
rect -3926 154894 -3306 190338
rect -3926 154658 -3894 154894
rect -3658 154658 -3574 154894
rect -3338 154658 -3306 154894
rect -3926 154574 -3306 154658
rect -3926 154338 -3894 154574
rect -3658 154338 -3574 154574
rect -3338 154338 -3306 154574
rect -3926 118894 -3306 154338
rect -3926 118658 -3894 118894
rect -3658 118658 -3574 118894
rect -3338 118658 -3306 118894
rect -3926 118574 -3306 118658
rect -3926 118338 -3894 118574
rect -3658 118338 -3574 118574
rect -3338 118338 -3306 118574
rect -3926 82894 -3306 118338
rect -3926 82658 -3894 82894
rect -3658 82658 -3574 82894
rect -3338 82658 -3306 82894
rect -3926 82574 -3306 82658
rect -3926 82338 -3894 82574
rect -3658 82338 -3574 82574
rect -3338 82338 -3306 82574
rect -3926 46894 -3306 82338
rect -3926 46658 -3894 46894
rect -3658 46658 -3574 46894
rect -3338 46658 -3306 46894
rect -3926 46574 -3306 46658
rect -3926 46338 -3894 46574
rect -3658 46338 -3574 46574
rect -3338 46338 -3306 46574
rect -3926 10894 -3306 46338
rect -3926 10658 -3894 10894
rect -3658 10658 -3574 10894
rect -3338 10658 -3306 10894
rect -3926 10574 -3306 10658
rect -3926 10338 -3894 10574
rect -3658 10338 -3574 10574
rect -3338 10338 -3306 10574
rect -3926 -2266 -3306 10338
rect -2966 705798 -2346 705830
rect -2966 705562 -2934 705798
rect -2698 705562 -2614 705798
rect -2378 705562 -2346 705798
rect -2966 705478 -2346 705562
rect -2966 705242 -2934 705478
rect -2698 705242 -2614 705478
rect -2378 705242 -2346 705478
rect -2966 691174 -2346 705242
rect -2966 690938 -2934 691174
rect -2698 690938 -2614 691174
rect -2378 690938 -2346 691174
rect -2966 690854 -2346 690938
rect -2966 690618 -2934 690854
rect -2698 690618 -2614 690854
rect -2378 690618 -2346 690854
rect -2966 655174 -2346 690618
rect -2966 654938 -2934 655174
rect -2698 654938 -2614 655174
rect -2378 654938 -2346 655174
rect -2966 654854 -2346 654938
rect -2966 654618 -2934 654854
rect -2698 654618 -2614 654854
rect -2378 654618 -2346 654854
rect -2966 619174 -2346 654618
rect -2966 618938 -2934 619174
rect -2698 618938 -2614 619174
rect -2378 618938 -2346 619174
rect -2966 618854 -2346 618938
rect -2966 618618 -2934 618854
rect -2698 618618 -2614 618854
rect -2378 618618 -2346 618854
rect -2966 583174 -2346 618618
rect -2966 582938 -2934 583174
rect -2698 582938 -2614 583174
rect -2378 582938 -2346 583174
rect -2966 582854 -2346 582938
rect -2966 582618 -2934 582854
rect -2698 582618 -2614 582854
rect -2378 582618 -2346 582854
rect -2966 547174 -2346 582618
rect -2966 546938 -2934 547174
rect -2698 546938 -2614 547174
rect -2378 546938 -2346 547174
rect -2966 546854 -2346 546938
rect -2966 546618 -2934 546854
rect -2698 546618 -2614 546854
rect -2378 546618 -2346 546854
rect -2966 511174 -2346 546618
rect -2966 510938 -2934 511174
rect -2698 510938 -2614 511174
rect -2378 510938 -2346 511174
rect -2966 510854 -2346 510938
rect -2966 510618 -2934 510854
rect -2698 510618 -2614 510854
rect -2378 510618 -2346 510854
rect -2966 475174 -2346 510618
rect -2966 474938 -2934 475174
rect -2698 474938 -2614 475174
rect -2378 474938 -2346 475174
rect -2966 474854 -2346 474938
rect -2966 474618 -2934 474854
rect -2698 474618 -2614 474854
rect -2378 474618 -2346 474854
rect -2966 439174 -2346 474618
rect -2966 438938 -2934 439174
rect -2698 438938 -2614 439174
rect -2378 438938 -2346 439174
rect -2966 438854 -2346 438938
rect -2966 438618 -2934 438854
rect -2698 438618 -2614 438854
rect -2378 438618 -2346 438854
rect -2966 403174 -2346 438618
rect -2966 402938 -2934 403174
rect -2698 402938 -2614 403174
rect -2378 402938 -2346 403174
rect -2966 402854 -2346 402938
rect -2966 402618 -2934 402854
rect -2698 402618 -2614 402854
rect -2378 402618 -2346 402854
rect -2966 367174 -2346 402618
rect -2966 366938 -2934 367174
rect -2698 366938 -2614 367174
rect -2378 366938 -2346 367174
rect -2966 366854 -2346 366938
rect -2966 366618 -2934 366854
rect -2698 366618 -2614 366854
rect -2378 366618 -2346 366854
rect -2966 331174 -2346 366618
rect -2966 330938 -2934 331174
rect -2698 330938 -2614 331174
rect -2378 330938 -2346 331174
rect -2966 330854 -2346 330938
rect -2966 330618 -2934 330854
rect -2698 330618 -2614 330854
rect -2378 330618 -2346 330854
rect -2966 295174 -2346 330618
rect -2966 294938 -2934 295174
rect -2698 294938 -2614 295174
rect -2378 294938 -2346 295174
rect -2966 294854 -2346 294938
rect -2966 294618 -2934 294854
rect -2698 294618 -2614 294854
rect -2378 294618 -2346 294854
rect -2966 259174 -2346 294618
rect -2966 258938 -2934 259174
rect -2698 258938 -2614 259174
rect -2378 258938 -2346 259174
rect -2966 258854 -2346 258938
rect -2966 258618 -2934 258854
rect -2698 258618 -2614 258854
rect -2378 258618 -2346 258854
rect -2966 223174 -2346 258618
rect -2966 222938 -2934 223174
rect -2698 222938 -2614 223174
rect -2378 222938 -2346 223174
rect -2966 222854 -2346 222938
rect -2966 222618 -2934 222854
rect -2698 222618 -2614 222854
rect -2378 222618 -2346 222854
rect -2966 187174 -2346 222618
rect -2966 186938 -2934 187174
rect -2698 186938 -2614 187174
rect -2378 186938 -2346 187174
rect -2966 186854 -2346 186938
rect -2966 186618 -2934 186854
rect -2698 186618 -2614 186854
rect -2378 186618 -2346 186854
rect -2966 151174 -2346 186618
rect -2966 150938 -2934 151174
rect -2698 150938 -2614 151174
rect -2378 150938 -2346 151174
rect -2966 150854 -2346 150938
rect -2966 150618 -2934 150854
rect -2698 150618 -2614 150854
rect -2378 150618 -2346 150854
rect -2966 115174 -2346 150618
rect -2966 114938 -2934 115174
rect -2698 114938 -2614 115174
rect -2378 114938 -2346 115174
rect -2966 114854 -2346 114938
rect -2966 114618 -2934 114854
rect -2698 114618 -2614 114854
rect -2378 114618 -2346 114854
rect -2966 79174 -2346 114618
rect -2966 78938 -2934 79174
rect -2698 78938 -2614 79174
rect -2378 78938 -2346 79174
rect -2966 78854 -2346 78938
rect -2966 78618 -2934 78854
rect -2698 78618 -2614 78854
rect -2378 78618 -2346 78854
rect -2966 43174 -2346 78618
rect -2966 42938 -2934 43174
rect -2698 42938 -2614 43174
rect -2378 42938 -2346 43174
rect -2966 42854 -2346 42938
rect -2966 42618 -2934 42854
rect -2698 42618 -2614 42854
rect -2378 42618 -2346 42854
rect -2966 7174 -2346 42618
rect -2966 6938 -2934 7174
rect -2698 6938 -2614 7174
rect -2378 6938 -2346 7174
rect -2966 6854 -2346 6938
rect -2966 6618 -2934 6854
rect -2698 6618 -2614 6854
rect -2378 6618 -2346 6854
rect -2966 -1306 -2346 6618
rect -2006 704838 -1386 704870
rect -2006 704602 -1974 704838
rect -1738 704602 -1654 704838
rect -1418 704602 -1386 704838
rect -2006 704518 -1386 704602
rect -2006 704282 -1974 704518
rect -1738 704282 -1654 704518
rect -1418 704282 -1386 704518
rect -2006 687454 -1386 704282
rect -2006 687218 -1974 687454
rect -1738 687218 -1654 687454
rect -1418 687218 -1386 687454
rect -2006 687134 -1386 687218
rect -2006 686898 -1974 687134
rect -1738 686898 -1654 687134
rect -1418 686898 -1386 687134
rect -2006 651454 -1386 686898
rect -2006 651218 -1974 651454
rect -1738 651218 -1654 651454
rect -1418 651218 -1386 651454
rect -2006 651134 -1386 651218
rect -2006 650898 -1974 651134
rect -1738 650898 -1654 651134
rect -1418 650898 -1386 651134
rect -2006 615454 -1386 650898
rect -2006 615218 -1974 615454
rect -1738 615218 -1654 615454
rect -1418 615218 -1386 615454
rect -2006 615134 -1386 615218
rect -2006 614898 -1974 615134
rect -1738 614898 -1654 615134
rect -1418 614898 -1386 615134
rect -2006 579454 -1386 614898
rect -2006 579218 -1974 579454
rect -1738 579218 -1654 579454
rect -1418 579218 -1386 579454
rect -2006 579134 -1386 579218
rect -2006 578898 -1974 579134
rect -1738 578898 -1654 579134
rect -1418 578898 -1386 579134
rect -2006 543454 -1386 578898
rect -2006 543218 -1974 543454
rect -1738 543218 -1654 543454
rect -1418 543218 -1386 543454
rect -2006 543134 -1386 543218
rect -2006 542898 -1974 543134
rect -1738 542898 -1654 543134
rect -1418 542898 -1386 543134
rect -2006 507454 -1386 542898
rect -2006 507218 -1974 507454
rect -1738 507218 -1654 507454
rect -1418 507218 -1386 507454
rect -2006 507134 -1386 507218
rect -2006 506898 -1974 507134
rect -1738 506898 -1654 507134
rect -1418 506898 -1386 507134
rect -2006 471454 -1386 506898
rect -2006 471218 -1974 471454
rect -1738 471218 -1654 471454
rect -1418 471218 -1386 471454
rect -2006 471134 -1386 471218
rect -2006 470898 -1974 471134
rect -1738 470898 -1654 471134
rect -1418 470898 -1386 471134
rect -2006 435454 -1386 470898
rect -2006 435218 -1974 435454
rect -1738 435218 -1654 435454
rect -1418 435218 -1386 435454
rect -2006 435134 -1386 435218
rect -2006 434898 -1974 435134
rect -1738 434898 -1654 435134
rect -1418 434898 -1386 435134
rect -2006 399454 -1386 434898
rect -2006 399218 -1974 399454
rect -1738 399218 -1654 399454
rect -1418 399218 -1386 399454
rect -2006 399134 -1386 399218
rect -2006 398898 -1974 399134
rect -1738 398898 -1654 399134
rect -1418 398898 -1386 399134
rect -2006 363454 -1386 398898
rect -2006 363218 -1974 363454
rect -1738 363218 -1654 363454
rect -1418 363218 -1386 363454
rect -2006 363134 -1386 363218
rect -2006 362898 -1974 363134
rect -1738 362898 -1654 363134
rect -1418 362898 -1386 363134
rect -2006 327454 -1386 362898
rect -2006 327218 -1974 327454
rect -1738 327218 -1654 327454
rect -1418 327218 -1386 327454
rect -2006 327134 -1386 327218
rect -2006 326898 -1974 327134
rect -1738 326898 -1654 327134
rect -1418 326898 -1386 327134
rect -2006 291454 -1386 326898
rect -2006 291218 -1974 291454
rect -1738 291218 -1654 291454
rect -1418 291218 -1386 291454
rect -2006 291134 -1386 291218
rect -2006 290898 -1974 291134
rect -1738 290898 -1654 291134
rect -1418 290898 -1386 291134
rect -2006 255454 -1386 290898
rect -2006 255218 -1974 255454
rect -1738 255218 -1654 255454
rect -1418 255218 -1386 255454
rect -2006 255134 -1386 255218
rect -2006 254898 -1974 255134
rect -1738 254898 -1654 255134
rect -1418 254898 -1386 255134
rect -2006 219454 -1386 254898
rect -2006 219218 -1974 219454
rect -1738 219218 -1654 219454
rect -1418 219218 -1386 219454
rect -2006 219134 -1386 219218
rect -2006 218898 -1974 219134
rect -1738 218898 -1654 219134
rect -1418 218898 -1386 219134
rect -2006 183454 -1386 218898
rect -2006 183218 -1974 183454
rect -1738 183218 -1654 183454
rect -1418 183218 -1386 183454
rect -2006 183134 -1386 183218
rect -2006 182898 -1974 183134
rect -1738 182898 -1654 183134
rect -1418 182898 -1386 183134
rect -2006 147454 -1386 182898
rect -2006 147218 -1974 147454
rect -1738 147218 -1654 147454
rect -1418 147218 -1386 147454
rect -2006 147134 -1386 147218
rect -2006 146898 -1974 147134
rect -1738 146898 -1654 147134
rect -1418 146898 -1386 147134
rect -2006 111454 -1386 146898
rect -2006 111218 -1974 111454
rect -1738 111218 -1654 111454
rect -1418 111218 -1386 111454
rect -2006 111134 -1386 111218
rect -2006 110898 -1974 111134
rect -1738 110898 -1654 111134
rect -1418 110898 -1386 111134
rect -2006 75454 -1386 110898
rect -2006 75218 -1974 75454
rect -1738 75218 -1654 75454
rect -1418 75218 -1386 75454
rect -2006 75134 -1386 75218
rect -2006 74898 -1974 75134
rect -1738 74898 -1654 75134
rect -1418 74898 -1386 75134
rect -2006 39454 -1386 74898
rect -2006 39218 -1974 39454
rect -1738 39218 -1654 39454
rect -1418 39218 -1386 39454
rect -2006 39134 -1386 39218
rect -2006 38898 -1974 39134
rect -1738 38898 -1654 39134
rect -1418 38898 -1386 39134
rect -2006 3454 -1386 38898
rect -2006 3218 -1974 3454
rect -1738 3218 -1654 3454
rect -1418 3218 -1386 3454
rect -2006 3134 -1386 3218
rect -2006 2898 -1974 3134
rect -1738 2898 -1654 3134
rect -1418 2898 -1386 3134
rect -2006 -346 -1386 2898
rect -2006 -582 -1974 -346
rect -1738 -582 -1654 -346
rect -1418 -582 -1386 -346
rect -2006 -666 -1386 -582
rect -2006 -902 -1974 -666
rect -1738 -902 -1654 -666
rect -1418 -902 -1386 -666
rect -2006 -934 -1386 -902
rect 1794 704838 2414 711590
rect 1794 704602 1826 704838
rect 2062 704602 2146 704838
rect 2382 704602 2414 704838
rect 1794 704518 2414 704602
rect 1794 704282 1826 704518
rect 2062 704282 2146 704518
rect 2382 704282 2414 704518
rect 1794 687454 2414 704282
rect 1794 687218 1826 687454
rect 2062 687218 2146 687454
rect 2382 687218 2414 687454
rect 1794 687134 2414 687218
rect 1794 686898 1826 687134
rect 2062 686898 2146 687134
rect 2382 686898 2414 687134
rect 1794 651454 2414 686898
rect 1794 651218 1826 651454
rect 2062 651218 2146 651454
rect 2382 651218 2414 651454
rect 1794 651134 2414 651218
rect 1794 650898 1826 651134
rect 2062 650898 2146 651134
rect 2382 650898 2414 651134
rect 1794 615454 2414 650898
rect 1794 615218 1826 615454
rect 2062 615218 2146 615454
rect 2382 615218 2414 615454
rect 1794 615134 2414 615218
rect 1794 614898 1826 615134
rect 2062 614898 2146 615134
rect 2382 614898 2414 615134
rect 1794 579454 2414 614898
rect 1794 579218 1826 579454
rect 2062 579218 2146 579454
rect 2382 579218 2414 579454
rect 1794 579134 2414 579218
rect 1794 578898 1826 579134
rect 2062 578898 2146 579134
rect 2382 578898 2414 579134
rect 1794 543454 2414 578898
rect 1794 543218 1826 543454
rect 2062 543218 2146 543454
rect 2382 543218 2414 543454
rect 1794 543134 2414 543218
rect 1794 542898 1826 543134
rect 2062 542898 2146 543134
rect 2382 542898 2414 543134
rect 1794 507454 2414 542898
rect 1794 507218 1826 507454
rect 2062 507218 2146 507454
rect 2382 507218 2414 507454
rect 1794 507134 2414 507218
rect 1794 506898 1826 507134
rect 2062 506898 2146 507134
rect 2382 506898 2414 507134
rect 1794 471454 2414 506898
rect 1794 471218 1826 471454
rect 2062 471218 2146 471454
rect 2382 471218 2414 471454
rect 1794 471134 2414 471218
rect 1794 470898 1826 471134
rect 2062 470898 2146 471134
rect 2382 470898 2414 471134
rect 1794 435454 2414 470898
rect 1794 435218 1826 435454
rect 2062 435218 2146 435454
rect 2382 435218 2414 435454
rect 1794 435134 2414 435218
rect 1794 434898 1826 435134
rect 2062 434898 2146 435134
rect 2382 434898 2414 435134
rect 1794 399454 2414 434898
rect 1794 399218 1826 399454
rect 2062 399218 2146 399454
rect 2382 399218 2414 399454
rect 1794 399134 2414 399218
rect 1794 398898 1826 399134
rect 2062 398898 2146 399134
rect 2382 398898 2414 399134
rect 1794 363454 2414 398898
rect 1794 363218 1826 363454
rect 2062 363218 2146 363454
rect 2382 363218 2414 363454
rect 1794 363134 2414 363218
rect 1794 362898 1826 363134
rect 2062 362898 2146 363134
rect 2382 362898 2414 363134
rect 1794 327454 2414 362898
rect 1794 327218 1826 327454
rect 2062 327218 2146 327454
rect 2382 327218 2414 327454
rect 1794 327134 2414 327218
rect 1794 326898 1826 327134
rect 2062 326898 2146 327134
rect 2382 326898 2414 327134
rect 1794 291454 2414 326898
rect 1794 291218 1826 291454
rect 2062 291218 2146 291454
rect 2382 291218 2414 291454
rect 1794 291134 2414 291218
rect 1794 290898 1826 291134
rect 2062 290898 2146 291134
rect 2382 290898 2414 291134
rect 1794 255454 2414 290898
rect 1794 255218 1826 255454
rect 2062 255218 2146 255454
rect 2382 255218 2414 255454
rect 1794 255134 2414 255218
rect 1794 254898 1826 255134
rect 2062 254898 2146 255134
rect 2382 254898 2414 255134
rect 1794 219454 2414 254898
rect 1794 219218 1826 219454
rect 2062 219218 2146 219454
rect 2382 219218 2414 219454
rect 1794 219134 2414 219218
rect 1794 218898 1826 219134
rect 2062 218898 2146 219134
rect 2382 218898 2414 219134
rect 1794 183454 2414 218898
rect 1794 183218 1826 183454
rect 2062 183218 2146 183454
rect 2382 183218 2414 183454
rect 1794 183134 2414 183218
rect 1794 182898 1826 183134
rect 2062 182898 2146 183134
rect 2382 182898 2414 183134
rect 1794 147454 2414 182898
rect 1794 147218 1826 147454
rect 2062 147218 2146 147454
rect 2382 147218 2414 147454
rect 1794 147134 2414 147218
rect 1794 146898 1826 147134
rect 2062 146898 2146 147134
rect 2382 146898 2414 147134
rect 1794 111454 2414 146898
rect 1794 111218 1826 111454
rect 2062 111218 2146 111454
rect 2382 111218 2414 111454
rect 1794 111134 2414 111218
rect 1794 110898 1826 111134
rect 2062 110898 2146 111134
rect 2382 110898 2414 111134
rect 1794 75454 2414 110898
rect 1794 75218 1826 75454
rect 2062 75218 2146 75454
rect 2382 75218 2414 75454
rect 1794 75134 2414 75218
rect 1794 74898 1826 75134
rect 2062 74898 2146 75134
rect 2382 74898 2414 75134
rect 1794 39454 2414 74898
rect 1794 39218 1826 39454
rect 2062 39218 2146 39454
rect 2382 39218 2414 39454
rect 1794 39134 2414 39218
rect 1794 38898 1826 39134
rect 2062 38898 2146 39134
rect 2382 38898 2414 39134
rect 1794 3454 2414 38898
rect 1794 3218 1826 3454
rect 2062 3218 2146 3454
rect 2382 3218 2414 3454
rect 1794 3134 2414 3218
rect 1794 2898 1826 3134
rect 2062 2898 2146 3134
rect 2382 2898 2414 3134
rect 1794 -346 2414 2898
rect 1794 -582 1826 -346
rect 2062 -582 2146 -346
rect 2382 -582 2414 -346
rect 1794 -666 2414 -582
rect 1794 -902 1826 -666
rect 2062 -902 2146 -666
rect 2382 -902 2414 -666
rect -2966 -1542 -2934 -1306
rect -2698 -1542 -2614 -1306
rect -2378 -1542 -2346 -1306
rect -2966 -1626 -2346 -1542
rect -2966 -1862 -2934 -1626
rect -2698 -1862 -2614 -1626
rect -2378 -1862 -2346 -1626
rect -2966 -1894 -2346 -1862
rect -3926 -2502 -3894 -2266
rect -3658 -2502 -3574 -2266
rect -3338 -2502 -3306 -2266
rect -3926 -2586 -3306 -2502
rect -3926 -2822 -3894 -2586
rect -3658 -2822 -3574 -2586
rect -3338 -2822 -3306 -2586
rect -3926 -2854 -3306 -2822
rect -4886 -3462 -4854 -3226
rect -4618 -3462 -4534 -3226
rect -4298 -3462 -4266 -3226
rect -4886 -3546 -4266 -3462
rect -4886 -3782 -4854 -3546
rect -4618 -3782 -4534 -3546
rect -4298 -3782 -4266 -3546
rect -4886 -3814 -4266 -3782
rect -5846 -4422 -5814 -4186
rect -5578 -4422 -5494 -4186
rect -5258 -4422 -5226 -4186
rect -5846 -4506 -5226 -4422
rect -5846 -4742 -5814 -4506
rect -5578 -4742 -5494 -4506
rect -5258 -4742 -5226 -4506
rect -5846 -4774 -5226 -4742
rect -6806 -5382 -6774 -5146
rect -6538 -5382 -6454 -5146
rect -6218 -5382 -6186 -5146
rect -6806 -5466 -6186 -5382
rect -6806 -5702 -6774 -5466
rect -6538 -5702 -6454 -5466
rect -6218 -5702 -6186 -5466
rect -6806 -5734 -6186 -5702
rect -7766 -6342 -7734 -6106
rect -7498 -6342 -7414 -6106
rect -7178 -6342 -7146 -6106
rect -7766 -6426 -7146 -6342
rect -7766 -6662 -7734 -6426
rect -7498 -6662 -7414 -6426
rect -7178 -6662 -7146 -6426
rect -7766 -6694 -7146 -6662
rect -8726 -7302 -8694 -7066
rect -8458 -7302 -8374 -7066
rect -8138 -7302 -8106 -7066
rect -8726 -7386 -8106 -7302
rect -8726 -7622 -8694 -7386
rect -8458 -7622 -8374 -7386
rect -8138 -7622 -8106 -7386
rect -8726 -7654 -8106 -7622
rect 1794 -7654 2414 -902
rect 5514 705798 6134 711590
rect 5514 705562 5546 705798
rect 5782 705562 5866 705798
rect 6102 705562 6134 705798
rect 5514 705478 6134 705562
rect 5514 705242 5546 705478
rect 5782 705242 5866 705478
rect 6102 705242 6134 705478
rect 5514 691174 6134 705242
rect 5514 690938 5546 691174
rect 5782 690938 5866 691174
rect 6102 690938 6134 691174
rect 5514 690854 6134 690938
rect 5514 690618 5546 690854
rect 5782 690618 5866 690854
rect 6102 690618 6134 690854
rect 5514 655174 6134 690618
rect 5514 654938 5546 655174
rect 5782 654938 5866 655174
rect 6102 654938 6134 655174
rect 5514 654854 6134 654938
rect 5514 654618 5546 654854
rect 5782 654618 5866 654854
rect 6102 654618 6134 654854
rect 5514 619174 6134 654618
rect 5514 618938 5546 619174
rect 5782 618938 5866 619174
rect 6102 618938 6134 619174
rect 5514 618854 6134 618938
rect 5514 618618 5546 618854
rect 5782 618618 5866 618854
rect 6102 618618 6134 618854
rect 5514 583174 6134 618618
rect 5514 582938 5546 583174
rect 5782 582938 5866 583174
rect 6102 582938 6134 583174
rect 5514 582854 6134 582938
rect 5514 582618 5546 582854
rect 5782 582618 5866 582854
rect 6102 582618 6134 582854
rect 5514 547174 6134 582618
rect 5514 546938 5546 547174
rect 5782 546938 5866 547174
rect 6102 546938 6134 547174
rect 5514 546854 6134 546938
rect 5514 546618 5546 546854
rect 5782 546618 5866 546854
rect 6102 546618 6134 546854
rect 5514 511174 6134 546618
rect 5514 510938 5546 511174
rect 5782 510938 5866 511174
rect 6102 510938 6134 511174
rect 5514 510854 6134 510938
rect 5514 510618 5546 510854
rect 5782 510618 5866 510854
rect 6102 510618 6134 510854
rect 5514 475174 6134 510618
rect 5514 474938 5546 475174
rect 5782 474938 5866 475174
rect 6102 474938 6134 475174
rect 5514 474854 6134 474938
rect 5514 474618 5546 474854
rect 5782 474618 5866 474854
rect 6102 474618 6134 474854
rect 5514 439174 6134 474618
rect 5514 438938 5546 439174
rect 5782 438938 5866 439174
rect 6102 438938 6134 439174
rect 5514 438854 6134 438938
rect 5514 438618 5546 438854
rect 5782 438618 5866 438854
rect 6102 438618 6134 438854
rect 5514 403174 6134 438618
rect 5514 402938 5546 403174
rect 5782 402938 5866 403174
rect 6102 402938 6134 403174
rect 5514 402854 6134 402938
rect 5514 402618 5546 402854
rect 5782 402618 5866 402854
rect 6102 402618 6134 402854
rect 5514 367174 6134 402618
rect 5514 366938 5546 367174
rect 5782 366938 5866 367174
rect 6102 366938 6134 367174
rect 5514 366854 6134 366938
rect 5514 366618 5546 366854
rect 5782 366618 5866 366854
rect 6102 366618 6134 366854
rect 5514 331174 6134 366618
rect 5514 330938 5546 331174
rect 5782 330938 5866 331174
rect 6102 330938 6134 331174
rect 5514 330854 6134 330938
rect 5514 330618 5546 330854
rect 5782 330618 5866 330854
rect 6102 330618 6134 330854
rect 5514 295174 6134 330618
rect 5514 294938 5546 295174
rect 5782 294938 5866 295174
rect 6102 294938 6134 295174
rect 5514 294854 6134 294938
rect 5514 294618 5546 294854
rect 5782 294618 5866 294854
rect 6102 294618 6134 294854
rect 5514 259174 6134 294618
rect 5514 258938 5546 259174
rect 5782 258938 5866 259174
rect 6102 258938 6134 259174
rect 5514 258854 6134 258938
rect 5514 258618 5546 258854
rect 5782 258618 5866 258854
rect 6102 258618 6134 258854
rect 5514 223174 6134 258618
rect 5514 222938 5546 223174
rect 5782 222938 5866 223174
rect 6102 222938 6134 223174
rect 5514 222854 6134 222938
rect 5514 222618 5546 222854
rect 5782 222618 5866 222854
rect 6102 222618 6134 222854
rect 5514 187174 6134 222618
rect 5514 186938 5546 187174
rect 5782 186938 5866 187174
rect 6102 186938 6134 187174
rect 5514 186854 6134 186938
rect 5514 186618 5546 186854
rect 5782 186618 5866 186854
rect 6102 186618 6134 186854
rect 5514 151174 6134 186618
rect 5514 150938 5546 151174
rect 5782 150938 5866 151174
rect 6102 150938 6134 151174
rect 5514 150854 6134 150938
rect 5514 150618 5546 150854
rect 5782 150618 5866 150854
rect 6102 150618 6134 150854
rect 5514 115174 6134 150618
rect 5514 114938 5546 115174
rect 5782 114938 5866 115174
rect 6102 114938 6134 115174
rect 5514 114854 6134 114938
rect 5514 114618 5546 114854
rect 5782 114618 5866 114854
rect 6102 114618 6134 114854
rect 5514 79174 6134 114618
rect 5514 78938 5546 79174
rect 5782 78938 5866 79174
rect 6102 78938 6134 79174
rect 5514 78854 6134 78938
rect 5514 78618 5546 78854
rect 5782 78618 5866 78854
rect 6102 78618 6134 78854
rect 5514 43174 6134 78618
rect 5514 42938 5546 43174
rect 5782 42938 5866 43174
rect 6102 42938 6134 43174
rect 5514 42854 6134 42938
rect 5514 42618 5546 42854
rect 5782 42618 5866 42854
rect 6102 42618 6134 42854
rect 5514 7174 6134 42618
rect 5514 6938 5546 7174
rect 5782 6938 5866 7174
rect 6102 6938 6134 7174
rect 5514 6854 6134 6938
rect 5514 6618 5546 6854
rect 5782 6618 5866 6854
rect 6102 6618 6134 6854
rect 5514 -1306 6134 6618
rect 5514 -1542 5546 -1306
rect 5782 -1542 5866 -1306
rect 6102 -1542 6134 -1306
rect 5514 -1626 6134 -1542
rect 5514 -1862 5546 -1626
rect 5782 -1862 5866 -1626
rect 6102 -1862 6134 -1626
rect 5514 -7654 6134 -1862
rect 9234 706758 9854 711590
rect 9234 706522 9266 706758
rect 9502 706522 9586 706758
rect 9822 706522 9854 706758
rect 9234 706438 9854 706522
rect 9234 706202 9266 706438
rect 9502 706202 9586 706438
rect 9822 706202 9854 706438
rect 9234 694894 9854 706202
rect 9234 694658 9266 694894
rect 9502 694658 9586 694894
rect 9822 694658 9854 694894
rect 9234 694574 9854 694658
rect 9234 694338 9266 694574
rect 9502 694338 9586 694574
rect 9822 694338 9854 694574
rect 9234 658894 9854 694338
rect 9234 658658 9266 658894
rect 9502 658658 9586 658894
rect 9822 658658 9854 658894
rect 9234 658574 9854 658658
rect 9234 658338 9266 658574
rect 9502 658338 9586 658574
rect 9822 658338 9854 658574
rect 9234 622894 9854 658338
rect 9234 622658 9266 622894
rect 9502 622658 9586 622894
rect 9822 622658 9854 622894
rect 9234 622574 9854 622658
rect 9234 622338 9266 622574
rect 9502 622338 9586 622574
rect 9822 622338 9854 622574
rect 9234 586894 9854 622338
rect 9234 586658 9266 586894
rect 9502 586658 9586 586894
rect 9822 586658 9854 586894
rect 9234 586574 9854 586658
rect 9234 586338 9266 586574
rect 9502 586338 9586 586574
rect 9822 586338 9854 586574
rect 9234 550894 9854 586338
rect 9234 550658 9266 550894
rect 9502 550658 9586 550894
rect 9822 550658 9854 550894
rect 9234 550574 9854 550658
rect 9234 550338 9266 550574
rect 9502 550338 9586 550574
rect 9822 550338 9854 550574
rect 9234 514894 9854 550338
rect 9234 514658 9266 514894
rect 9502 514658 9586 514894
rect 9822 514658 9854 514894
rect 9234 514574 9854 514658
rect 9234 514338 9266 514574
rect 9502 514338 9586 514574
rect 9822 514338 9854 514574
rect 9234 478894 9854 514338
rect 9234 478658 9266 478894
rect 9502 478658 9586 478894
rect 9822 478658 9854 478894
rect 9234 478574 9854 478658
rect 9234 478338 9266 478574
rect 9502 478338 9586 478574
rect 9822 478338 9854 478574
rect 9234 442894 9854 478338
rect 9234 442658 9266 442894
rect 9502 442658 9586 442894
rect 9822 442658 9854 442894
rect 9234 442574 9854 442658
rect 9234 442338 9266 442574
rect 9502 442338 9586 442574
rect 9822 442338 9854 442574
rect 9234 406894 9854 442338
rect 9234 406658 9266 406894
rect 9502 406658 9586 406894
rect 9822 406658 9854 406894
rect 9234 406574 9854 406658
rect 9234 406338 9266 406574
rect 9502 406338 9586 406574
rect 9822 406338 9854 406574
rect 9234 370894 9854 406338
rect 9234 370658 9266 370894
rect 9502 370658 9586 370894
rect 9822 370658 9854 370894
rect 9234 370574 9854 370658
rect 9234 370338 9266 370574
rect 9502 370338 9586 370574
rect 9822 370338 9854 370574
rect 9234 334894 9854 370338
rect 9234 334658 9266 334894
rect 9502 334658 9586 334894
rect 9822 334658 9854 334894
rect 9234 334574 9854 334658
rect 9234 334338 9266 334574
rect 9502 334338 9586 334574
rect 9822 334338 9854 334574
rect 9234 298894 9854 334338
rect 9234 298658 9266 298894
rect 9502 298658 9586 298894
rect 9822 298658 9854 298894
rect 9234 298574 9854 298658
rect 9234 298338 9266 298574
rect 9502 298338 9586 298574
rect 9822 298338 9854 298574
rect 9234 262894 9854 298338
rect 9234 262658 9266 262894
rect 9502 262658 9586 262894
rect 9822 262658 9854 262894
rect 9234 262574 9854 262658
rect 9234 262338 9266 262574
rect 9502 262338 9586 262574
rect 9822 262338 9854 262574
rect 9234 226894 9854 262338
rect 9234 226658 9266 226894
rect 9502 226658 9586 226894
rect 9822 226658 9854 226894
rect 9234 226574 9854 226658
rect 9234 226338 9266 226574
rect 9502 226338 9586 226574
rect 9822 226338 9854 226574
rect 9234 190894 9854 226338
rect 9234 190658 9266 190894
rect 9502 190658 9586 190894
rect 9822 190658 9854 190894
rect 9234 190574 9854 190658
rect 9234 190338 9266 190574
rect 9502 190338 9586 190574
rect 9822 190338 9854 190574
rect 9234 154894 9854 190338
rect 9234 154658 9266 154894
rect 9502 154658 9586 154894
rect 9822 154658 9854 154894
rect 9234 154574 9854 154658
rect 9234 154338 9266 154574
rect 9502 154338 9586 154574
rect 9822 154338 9854 154574
rect 9234 118894 9854 154338
rect 9234 118658 9266 118894
rect 9502 118658 9586 118894
rect 9822 118658 9854 118894
rect 9234 118574 9854 118658
rect 9234 118338 9266 118574
rect 9502 118338 9586 118574
rect 9822 118338 9854 118574
rect 9234 82894 9854 118338
rect 9234 82658 9266 82894
rect 9502 82658 9586 82894
rect 9822 82658 9854 82894
rect 9234 82574 9854 82658
rect 9234 82338 9266 82574
rect 9502 82338 9586 82574
rect 9822 82338 9854 82574
rect 9234 46894 9854 82338
rect 9234 46658 9266 46894
rect 9502 46658 9586 46894
rect 9822 46658 9854 46894
rect 9234 46574 9854 46658
rect 9234 46338 9266 46574
rect 9502 46338 9586 46574
rect 9822 46338 9854 46574
rect 9234 10894 9854 46338
rect 9234 10658 9266 10894
rect 9502 10658 9586 10894
rect 9822 10658 9854 10894
rect 9234 10574 9854 10658
rect 9234 10338 9266 10574
rect 9502 10338 9586 10574
rect 9822 10338 9854 10574
rect 9234 -2266 9854 10338
rect 9234 -2502 9266 -2266
rect 9502 -2502 9586 -2266
rect 9822 -2502 9854 -2266
rect 9234 -2586 9854 -2502
rect 9234 -2822 9266 -2586
rect 9502 -2822 9586 -2586
rect 9822 -2822 9854 -2586
rect 9234 -7654 9854 -2822
rect 12954 707718 13574 711590
rect 12954 707482 12986 707718
rect 13222 707482 13306 707718
rect 13542 707482 13574 707718
rect 12954 707398 13574 707482
rect 12954 707162 12986 707398
rect 13222 707162 13306 707398
rect 13542 707162 13574 707398
rect 12954 698614 13574 707162
rect 12954 698378 12986 698614
rect 13222 698378 13306 698614
rect 13542 698378 13574 698614
rect 12954 698294 13574 698378
rect 12954 698058 12986 698294
rect 13222 698058 13306 698294
rect 13542 698058 13574 698294
rect 12954 662614 13574 698058
rect 12954 662378 12986 662614
rect 13222 662378 13306 662614
rect 13542 662378 13574 662614
rect 12954 662294 13574 662378
rect 12954 662058 12986 662294
rect 13222 662058 13306 662294
rect 13542 662058 13574 662294
rect 12954 626614 13574 662058
rect 12954 626378 12986 626614
rect 13222 626378 13306 626614
rect 13542 626378 13574 626614
rect 12954 626294 13574 626378
rect 12954 626058 12986 626294
rect 13222 626058 13306 626294
rect 13542 626058 13574 626294
rect 12954 590614 13574 626058
rect 12954 590378 12986 590614
rect 13222 590378 13306 590614
rect 13542 590378 13574 590614
rect 12954 590294 13574 590378
rect 12954 590058 12986 590294
rect 13222 590058 13306 590294
rect 13542 590058 13574 590294
rect 12954 554614 13574 590058
rect 12954 554378 12986 554614
rect 13222 554378 13306 554614
rect 13542 554378 13574 554614
rect 12954 554294 13574 554378
rect 12954 554058 12986 554294
rect 13222 554058 13306 554294
rect 13542 554058 13574 554294
rect 12954 518614 13574 554058
rect 12954 518378 12986 518614
rect 13222 518378 13306 518614
rect 13542 518378 13574 518614
rect 12954 518294 13574 518378
rect 12954 518058 12986 518294
rect 13222 518058 13306 518294
rect 13542 518058 13574 518294
rect 12954 482614 13574 518058
rect 12954 482378 12986 482614
rect 13222 482378 13306 482614
rect 13542 482378 13574 482614
rect 12954 482294 13574 482378
rect 12954 482058 12986 482294
rect 13222 482058 13306 482294
rect 13542 482058 13574 482294
rect 12954 446614 13574 482058
rect 12954 446378 12986 446614
rect 13222 446378 13306 446614
rect 13542 446378 13574 446614
rect 12954 446294 13574 446378
rect 12954 446058 12986 446294
rect 13222 446058 13306 446294
rect 13542 446058 13574 446294
rect 12954 410614 13574 446058
rect 12954 410378 12986 410614
rect 13222 410378 13306 410614
rect 13542 410378 13574 410614
rect 12954 410294 13574 410378
rect 12954 410058 12986 410294
rect 13222 410058 13306 410294
rect 13542 410058 13574 410294
rect 12954 374614 13574 410058
rect 12954 374378 12986 374614
rect 13222 374378 13306 374614
rect 13542 374378 13574 374614
rect 12954 374294 13574 374378
rect 12954 374058 12986 374294
rect 13222 374058 13306 374294
rect 13542 374058 13574 374294
rect 12954 338614 13574 374058
rect 12954 338378 12986 338614
rect 13222 338378 13306 338614
rect 13542 338378 13574 338614
rect 12954 338294 13574 338378
rect 12954 338058 12986 338294
rect 13222 338058 13306 338294
rect 13542 338058 13574 338294
rect 12954 302614 13574 338058
rect 12954 302378 12986 302614
rect 13222 302378 13306 302614
rect 13542 302378 13574 302614
rect 12954 302294 13574 302378
rect 12954 302058 12986 302294
rect 13222 302058 13306 302294
rect 13542 302058 13574 302294
rect 12954 266614 13574 302058
rect 12954 266378 12986 266614
rect 13222 266378 13306 266614
rect 13542 266378 13574 266614
rect 12954 266294 13574 266378
rect 12954 266058 12986 266294
rect 13222 266058 13306 266294
rect 13542 266058 13574 266294
rect 12954 230614 13574 266058
rect 12954 230378 12986 230614
rect 13222 230378 13306 230614
rect 13542 230378 13574 230614
rect 12954 230294 13574 230378
rect 12954 230058 12986 230294
rect 13222 230058 13306 230294
rect 13542 230058 13574 230294
rect 12954 194614 13574 230058
rect 12954 194378 12986 194614
rect 13222 194378 13306 194614
rect 13542 194378 13574 194614
rect 12954 194294 13574 194378
rect 12954 194058 12986 194294
rect 13222 194058 13306 194294
rect 13542 194058 13574 194294
rect 12954 158614 13574 194058
rect 12954 158378 12986 158614
rect 13222 158378 13306 158614
rect 13542 158378 13574 158614
rect 12954 158294 13574 158378
rect 12954 158058 12986 158294
rect 13222 158058 13306 158294
rect 13542 158058 13574 158294
rect 12954 122614 13574 158058
rect 12954 122378 12986 122614
rect 13222 122378 13306 122614
rect 13542 122378 13574 122614
rect 12954 122294 13574 122378
rect 12954 122058 12986 122294
rect 13222 122058 13306 122294
rect 13542 122058 13574 122294
rect 12954 86614 13574 122058
rect 12954 86378 12986 86614
rect 13222 86378 13306 86614
rect 13542 86378 13574 86614
rect 12954 86294 13574 86378
rect 12954 86058 12986 86294
rect 13222 86058 13306 86294
rect 13542 86058 13574 86294
rect 12954 50614 13574 86058
rect 12954 50378 12986 50614
rect 13222 50378 13306 50614
rect 13542 50378 13574 50614
rect 12954 50294 13574 50378
rect 12954 50058 12986 50294
rect 13222 50058 13306 50294
rect 13542 50058 13574 50294
rect 12954 14614 13574 50058
rect 12954 14378 12986 14614
rect 13222 14378 13306 14614
rect 13542 14378 13574 14614
rect 12954 14294 13574 14378
rect 12954 14058 12986 14294
rect 13222 14058 13306 14294
rect 13542 14058 13574 14294
rect 12954 -3226 13574 14058
rect 12954 -3462 12986 -3226
rect 13222 -3462 13306 -3226
rect 13542 -3462 13574 -3226
rect 12954 -3546 13574 -3462
rect 12954 -3782 12986 -3546
rect 13222 -3782 13306 -3546
rect 13542 -3782 13574 -3546
rect 12954 -7654 13574 -3782
rect 16674 708678 17294 711590
rect 16674 708442 16706 708678
rect 16942 708442 17026 708678
rect 17262 708442 17294 708678
rect 16674 708358 17294 708442
rect 16674 708122 16706 708358
rect 16942 708122 17026 708358
rect 17262 708122 17294 708358
rect 16674 666334 17294 708122
rect 16674 666098 16706 666334
rect 16942 666098 17026 666334
rect 17262 666098 17294 666334
rect 16674 666014 17294 666098
rect 16674 665778 16706 666014
rect 16942 665778 17026 666014
rect 17262 665778 17294 666014
rect 16674 630334 17294 665778
rect 16674 630098 16706 630334
rect 16942 630098 17026 630334
rect 17262 630098 17294 630334
rect 16674 630014 17294 630098
rect 16674 629778 16706 630014
rect 16942 629778 17026 630014
rect 17262 629778 17294 630014
rect 16674 594334 17294 629778
rect 16674 594098 16706 594334
rect 16942 594098 17026 594334
rect 17262 594098 17294 594334
rect 16674 594014 17294 594098
rect 16674 593778 16706 594014
rect 16942 593778 17026 594014
rect 17262 593778 17294 594014
rect 16674 558334 17294 593778
rect 16674 558098 16706 558334
rect 16942 558098 17026 558334
rect 17262 558098 17294 558334
rect 16674 558014 17294 558098
rect 16674 557778 16706 558014
rect 16942 557778 17026 558014
rect 17262 557778 17294 558014
rect 16674 522334 17294 557778
rect 16674 522098 16706 522334
rect 16942 522098 17026 522334
rect 17262 522098 17294 522334
rect 16674 522014 17294 522098
rect 16674 521778 16706 522014
rect 16942 521778 17026 522014
rect 17262 521778 17294 522014
rect 16674 486334 17294 521778
rect 16674 486098 16706 486334
rect 16942 486098 17026 486334
rect 17262 486098 17294 486334
rect 16674 486014 17294 486098
rect 16674 485778 16706 486014
rect 16942 485778 17026 486014
rect 17262 485778 17294 486014
rect 16674 450334 17294 485778
rect 16674 450098 16706 450334
rect 16942 450098 17026 450334
rect 17262 450098 17294 450334
rect 16674 450014 17294 450098
rect 16674 449778 16706 450014
rect 16942 449778 17026 450014
rect 17262 449778 17294 450014
rect 16674 414334 17294 449778
rect 16674 414098 16706 414334
rect 16942 414098 17026 414334
rect 17262 414098 17294 414334
rect 16674 414014 17294 414098
rect 16674 413778 16706 414014
rect 16942 413778 17026 414014
rect 17262 413778 17294 414014
rect 16674 378334 17294 413778
rect 16674 378098 16706 378334
rect 16942 378098 17026 378334
rect 17262 378098 17294 378334
rect 16674 378014 17294 378098
rect 16674 377778 16706 378014
rect 16942 377778 17026 378014
rect 17262 377778 17294 378014
rect 16674 342334 17294 377778
rect 16674 342098 16706 342334
rect 16942 342098 17026 342334
rect 17262 342098 17294 342334
rect 16674 342014 17294 342098
rect 16674 341778 16706 342014
rect 16942 341778 17026 342014
rect 17262 341778 17294 342014
rect 16674 306334 17294 341778
rect 16674 306098 16706 306334
rect 16942 306098 17026 306334
rect 17262 306098 17294 306334
rect 16674 306014 17294 306098
rect 16674 305778 16706 306014
rect 16942 305778 17026 306014
rect 17262 305778 17294 306014
rect 16674 270334 17294 305778
rect 16674 270098 16706 270334
rect 16942 270098 17026 270334
rect 17262 270098 17294 270334
rect 16674 270014 17294 270098
rect 16674 269778 16706 270014
rect 16942 269778 17026 270014
rect 17262 269778 17294 270014
rect 16674 234334 17294 269778
rect 16674 234098 16706 234334
rect 16942 234098 17026 234334
rect 17262 234098 17294 234334
rect 16674 234014 17294 234098
rect 16674 233778 16706 234014
rect 16942 233778 17026 234014
rect 17262 233778 17294 234014
rect 16674 198334 17294 233778
rect 16674 198098 16706 198334
rect 16942 198098 17026 198334
rect 17262 198098 17294 198334
rect 16674 198014 17294 198098
rect 16674 197778 16706 198014
rect 16942 197778 17026 198014
rect 17262 197778 17294 198014
rect 16674 162334 17294 197778
rect 16674 162098 16706 162334
rect 16942 162098 17026 162334
rect 17262 162098 17294 162334
rect 16674 162014 17294 162098
rect 16674 161778 16706 162014
rect 16942 161778 17026 162014
rect 17262 161778 17294 162014
rect 16674 126334 17294 161778
rect 16674 126098 16706 126334
rect 16942 126098 17026 126334
rect 17262 126098 17294 126334
rect 16674 126014 17294 126098
rect 16674 125778 16706 126014
rect 16942 125778 17026 126014
rect 17262 125778 17294 126014
rect 16674 90334 17294 125778
rect 16674 90098 16706 90334
rect 16942 90098 17026 90334
rect 17262 90098 17294 90334
rect 16674 90014 17294 90098
rect 16674 89778 16706 90014
rect 16942 89778 17026 90014
rect 17262 89778 17294 90014
rect 16674 54334 17294 89778
rect 16674 54098 16706 54334
rect 16942 54098 17026 54334
rect 17262 54098 17294 54334
rect 16674 54014 17294 54098
rect 16674 53778 16706 54014
rect 16942 53778 17026 54014
rect 17262 53778 17294 54014
rect 16674 18334 17294 53778
rect 16674 18098 16706 18334
rect 16942 18098 17026 18334
rect 17262 18098 17294 18334
rect 16674 18014 17294 18098
rect 16674 17778 16706 18014
rect 16942 17778 17026 18014
rect 17262 17778 17294 18014
rect 16674 -4186 17294 17778
rect 16674 -4422 16706 -4186
rect 16942 -4422 17026 -4186
rect 17262 -4422 17294 -4186
rect 16674 -4506 17294 -4422
rect 16674 -4742 16706 -4506
rect 16942 -4742 17026 -4506
rect 17262 -4742 17294 -4506
rect 16674 -7654 17294 -4742
rect 20394 709638 21014 711590
rect 20394 709402 20426 709638
rect 20662 709402 20746 709638
rect 20982 709402 21014 709638
rect 20394 709318 21014 709402
rect 20394 709082 20426 709318
rect 20662 709082 20746 709318
rect 20982 709082 21014 709318
rect 20394 670054 21014 709082
rect 20394 669818 20426 670054
rect 20662 669818 20746 670054
rect 20982 669818 21014 670054
rect 20394 669734 21014 669818
rect 20394 669498 20426 669734
rect 20662 669498 20746 669734
rect 20982 669498 21014 669734
rect 20394 634054 21014 669498
rect 20394 633818 20426 634054
rect 20662 633818 20746 634054
rect 20982 633818 21014 634054
rect 20394 633734 21014 633818
rect 20394 633498 20426 633734
rect 20662 633498 20746 633734
rect 20982 633498 21014 633734
rect 20394 598054 21014 633498
rect 20394 597818 20426 598054
rect 20662 597818 20746 598054
rect 20982 597818 21014 598054
rect 20394 597734 21014 597818
rect 20394 597498 20426 597734
rect 20662 597498 20746 597734
rect 20982 597498 21014 597734
rect 20394 562054 21014 597498
rect 20394 561818 20426 562054
rect 20662 561818 20746 562054
rect 20982 561818 21014 562054
rect 20394 561734 21014 561818
rect 20394 561498 20426 561734
rect 20662 561498 20746 561734
rect 20982 561498 21014 561734
rect 20394 526054 21014 561498
rect 20394 525818 20426 526054
rect 20662 525818 20746 526054
rect 20982 525818 21014 526054
rect 20394 525734 21014 525818
rect 20394 525498 20426 525734
rect 20662 525498 20746 525734
rect 20982 525498 21014 525734
rect 20394 490054 21014 525498
rect 20394 489818 20426 490054
rect 20662 489818 20746 490054
rect 20982 489818 21014 490054
rect 20394 489734 21014 489818
rect 20394 489498 20426 489734
rect 20662 489498 20746 489734
rect 20982 489498 21014 489734
rect 20394 454054 21014 489498
rect 20394 453818 20426 454054
rect 20662 453818 20746 454054
rect 20982 453818 21014 454054
rect 20394 453734 21014 453818
rect 20394 453498 20426 453734
rect 20662 453498 20746 453734
rect 20982 453498 21014 453734
rect 20394 418054 21014 453498
rect 20394 417818 20426 418054
rect 20662 417818 20746 418054
rect 20982 417818 21014 418054
rect 20394 417734 21014 417818
rect 20394 417498 20426 417734
rect 20662 417498 20746 417734
rect 20982 417498 21014 417734
rect 20394 382054 21014 417498
rect 20394 381818 20426 382054
rect 20662 381818 20746 382054
rect 20982 381818 21014 382054
rect 20394 381734 21014 381818
rect 20394 381498 20426 381734
rect 20662 381498 20746 381734
rect 20982 381498 21014 381734
rect 20394 346054 21014 381498
rect 20394 345818 20426 346054
rect 20662 345818 20746 346054
rect 20982 345818 21014 346054
rect 20394 345734 21014 345818
rect 20394 345498 20426 345734
rect 20662 345498 20746 345734
rect 20982 345498 21014 345734
rect 20394 310054 21014 345498
rect 20394 309818 20426 310054
rect 20662 309818 20746 310054
rect 20982 309818 21014 310054
rect 20394 309734 21014 309818
rect 20394 309498 20426 309734
rect 20662 309498 20746 309734
rect 20982 309498 21014 309734
rect 20394 274054 21014 309498
rect 20394 273818 20426 274054
rect 20662 273818 20746 274054
rect 20982 273818 21014 274054
rect 20394 273734 21014 273818
rect 20394 273498 20426 273734
rect 20662 273498 20746 273734
rect 20982 273498 21014 273734
rect 20394 238054 21014 273498
rect 20394 237818 20426 238054
rect 20662 237818 20746 238054
rect 20982 237818 21014 238054
rect 20394 237734 21014 237818
rect 20394 237498 20426 237734
rect 20662 237498 20746 237734
rect 20982 237498 21014 237734
rect 20394 202054 21014 237498
rect 20394 201818 20426 202054
rect 20662 201818 20746 202054
rect 20982 201818 21014 202054
rect 20394 201734 21014 201818
rect 20394 201498 20426 201734
rect 20662 201498 20746 201734
rect 20982 201498 21014 201734
rect 20394 166054 21014 201498
rect 20394 165818 20426 166054
rect 20662 165818 20746 166054
rect 20982 165818 21014 166054
rect 20394 165734 21014 165818
rect 20394 165498 20426 165734
rect 20662 165498 20746 165734
rect 20982 165498 21014 165734
rect 20394 130054 21014 165498
rect 20394 129818 20426 130054
rect 20662 129818 20746 130054
rect 20982 129818 21014 130054
rect 20394 129734 21014 129818
rect 20394 129498 20426 129734
rect 20662 129498 20746 129734
rect 20982 129498 21014 129734
rect 20394 94054 21014 129498
rect 20394 93818 20426 94054
rect 20662 93818 20746 94054
rect 20982 93818 21014 94054
rect 20394 93734 21014 93818
rect 20394 93498 20426 93734
rect 20662 93498 20746 93734
rect 20982 93498 21014 93734
rect 20394 58054 21014 93498
rect 20394 57818 20426 58054
rect 20662 57818 20746 58054
rect 20982 57818 21014 58054
rect 20394 57734 21014 57818
rect 20394 57498 20426 57734
rect 20662 57498 20746 57734
rect 20982 57498 21014 57734
rect 20394 22054 21014 57498
rect 20394 21818 20426 22054
rect 20662 21818 20746 22054
rect 20982 21818 21014 22054
rect 20394 21734 21014 21818
rect 20394 21498 20426 21734
rect 20662 21498 20746 21734
rect 20982 21498 21014 21734
rect 20394 -5146 21014 21498
rect 20394 -5382 20426 -5146
rect 20662 -5382 20746 -5146
rect 20982 -5382 21014 -5146
rect 20394 -5466 21014 -5382
rect 20394 -5702 20426 -5466
rect 20662 -5702 20746 -5466
rect 20982 -5702 21014 -5466
rect 20394 -7654 21014 -5702
rect 24114 710598 24734 711590
rect 24114 710362 24146 710598
rect 24382 710362 24466 710598
rect 24702 710362 24734 710598
rect 24114 710278 24734 710362
rect 24114 710042 24146 710278
rect 24382 710042 24466 710278
rect 24702 710042 24734 710278
rect 24114 673774 24734 710042
rect 24114 673538 24146 673774
rect 24382 673538 24466 673774
rect 24702 673538 24734 673774
rect 24114 673454 24734 673538
rect 24114 673218 24146 673454
rect 24382 673218 24466 673454
rect 24702 673218 24734 673454
rect 24114 637774 24734 673218
rect 24114 637538 24146 637774
rect 24382 637538 24466 637774
rect 24702 637538 24734 637774
rect 24114 637454 24734 637538
rect 24114 637218 24146 637454
rect 24382 637218 24466 637454
rect 24702 637218 24734 637454
rect 24114 601774 24734 637218
rect 24114 601538 24146 601774
rect 24382 601538 24466 601774
rect 24702 601538 24734 601774
rect 24114 601454 24734 601538
rect 24114 601218 24146 601454
rect 24382 601218 24466 601454
rect 24702 601218 24734 601454
rect 24114 565774 24734 601218
rect 24114 565538 24146 565774
rect 24382 565538 24466 565774
rect 24702 565538 24734 565774
rect 24114 565454 24734 565538
rect 24114 565218 24146 565454
rect 24382 565218 24466 565454
rect 24702 565218 24734 565454
rect 24114 529774 24734 565218
rect 24114 529538 24146 529774
rect 24382 529538 24466 529774
rect 24702 529538 24734 529774
rect 24114 529454 24734 529538
rect 24114 529218 24146 529454
rect 24382 529218 24466 529454
rect 24702 529218 24734 529454
rect 24114 493774 24734 529218
rect 24114 493538 24146 493774
rect 24382 493538 24466 493774
rect 24702 493538 24734 493774
rect 24114 493454 24734 493538
rect 24114 493218 24146 493454
rect 24382 493218 24466 493454
rect 24702 493218 24734 493454
rect 24114 457774 24734 493218
rect 24114 457538 24146 457774
rect 24382 457538 24466 457774
rect 24702 457538 24734 457774
rect 24114 457454 24734 457538
rect 24114 457218 24146 457454
rect 24382 457218 24466 457454
rect 24702 457218 24734 457454
rect 24114 421774 24734 457218
rect 24114 421538 24146 421774
rect 24382 421538 24466 421774
rect 24702 421538 24734 421774
rect 24114 421454 24734 421538
rect 24114 421218 24146 421454
rect 24382 421218 24466 421454
rect 24702 421218 24734 421454
rect 24114 385774 24734 421218
rect 24114 385538 24146 385774
rect 24382 385538 24466 385774
rect 24702 385538 24734 385774
rect 24114 385454 24734 385538
rect 24114 385218 24146 385454
rect 24382 385218 24466 385454
rect 24702 385218 24734 385454
rect 24114 349774 24734 385218
rect 24114 349538 24146 349774
rect 24382 349538 24466 349774
rect 24702 349538 24734 349774
rect 24114 349454 24734 349538
rect 24114 349218 24146 349454
rect 24382 349218 24466 349454
rect 24702 349218 24734 349454
rect 24114 313774 24734 349218
rect 24114 313538 24146 313774
rect 24382 313538 24466 313774
rect 24702 313538 24734 313774
rect 24114 313454 24734 313538
rect 24114 313218 24146 313454
rect 24382 313218 24466 313454
rect 24702 313218 24734 313454
rect 24114 277774 24734 313218
rect 24114 277538 24146 277774
rect 24382 277538 24466 277774
rect 24702 277538 24734 277774
rect 24114 277454 24734 277538
rect 24114 277218 24146 277454
rect 24382 277218 24466 277454
rect 24702 277218 24734 277454
rect 24114 241774 24734 277218
rect 24114 241538 24146 241774
rect 24382 241538 24466 241774
rect 24702 241538 24734 241774
rect 24114 241454 24734 241538
rect 24114 241218 24146 241454
rect 24382 241218 24466 241454
rect 24702 241218 24734 241454
rect 24114 205774 24734 241218
rect 24114 205538 24146 205774
rect 24382 205538 24466 205774
rect 24702 205538 24734 205774
rect 24114 205454 24734 205538
rect 24114 205218 24146 205454
rect 24382 205218 24466 205454
rect 24702 205218 24734 205454
rect 24114 169774 24734 205218
rect 24114 169538 24146 169774
rect 24382 169538 24466 169774
rect 24702 169538 24734 169774
rect 24114 169454 24734 169538
rect 24114 169218 24146 169454
rect 24382 169218 24466 169454
rect 24702 169218 24734 169454
rect 24114 133774 24734 169218
rect 27834 711558 28454 711590
rect 27834 711322 27866 711558
rect 28102 711322 28186 711558
rect 28422 711322 28454 711558
rect 27834 711238 28454 711322
rect 27834 711002 27866 711238
rect 28102 711002 28186 711238
rect 28422 711002 28454 711238
rect 27834 677494 28454 711002
rect 27834 677258 27866 677494
rect 28102 677258 28186 677494
rect 28422 677258 28454 677494
rect 27834 677174 28454 677258
rect 27834 676938 27866 677174
rect 28102 676938 28186 677174
rect 28422 676938 28454 677174
rect 27834 641494 28454 676938
rect 27834 641258 27866 641494
rect 28102 641258 28186 641494
rect 28422 641258 28454 641494
rect 27834 641174 28454 641258
rect 27834 640938 27866 641174
rect 28102 640938 28186 641174
rect 28422 640938 28454 641174
rect 27834 605494 28454 640938
rect 27834 605258 27866 605494
rect 28102 605258 28186 605494
rect 28422 605258 28454 605494
rect 27834 605174 28454 605258
rect 27834 604938 27866 605174
rect 28102 604938 28186 605174
rect 28422 604938 28454 605174
rect 27834 569494 28454 604938
rect 37794 704838 38414 711590
rect 37794 704602 37826 704838
rect 38062 704602 38146 704838
rect 38382 704602 38414 704838
rect 37794 704518 38414 704602
rect 37794 704282 37826 704518
rect 38062 704282 38146 704518
rect 38382 704282 38414 704518
rect 37794 687454 38414 704282
rect 37794 687218 37826 687454
rect 38062 687218 38146 687454
rect 38382 687218 38414 687454
rect 37794 687134 38414 687218
rect 37794 686898 37826 687134
rect 38062 686898 38146 687134
rect 38382 686898 38414 687134
rect 37794 651454 38414 686898
rect 37794 651218 37826 651454
rect 38062 651218 38146 651454
rect 38382 651218 38414 651454
rect 37794 651134 38414 651218
rect 37794 650898 37826 651134
rect 38062 650898 38146 651134
rect 38382 650898 38414 651134
rect 37794 615454 38414 650898
rect 37794 615218 37826 615454
rect 38062 615218 38146 615454
rect 38382 615218 38414 615454
rect 37794 615134 38414 615218
rect 37794 614898 37826 615134
rect 38062 614898 38146 615134
rect 38382 614898 38414 615134
rect 34208 579454 34528 579486
rect 34208 579218 34250 579454
rect 34486 579218 34528 579454
rect 34208 579134 34528 579218
rect 34208 578898 34250 579134
rect 34486 578898 34528 579134
rect 34208 578866 34528 578898
rect 37794 579454 38414 614898
rect 37794 579218 37826 579454
rect 38062 579218 38146 579454
rect 38382 579218 38414 579454
rect 37794 579134 38414 579218
rect 37794 578898 37826 579134
rect 38062 578898 38146 579134
rect 38382 578898 38414 579134
rect 27834 569258 27866 569494
rect 28102 569258 28186 569494
rect 28422 569258 28454 569494
rect 27834 569174 28454 569258
rect 27834 568938 27866 569174
rect 28102 568938 28186 569174
rect 28422 568938 28454 569174
rect 27834 533494 28454 568938
rect 34208 543454 34528 543486
rect 34208 543218 34250 543454
rect 34486 543218 34528 543454
rect 34208 543134 34528 543218
rect 34208 542898 34250 543134
rect 34486 542898 34528 543134
rect 34208 542866 34528 542898
rect 37794 543454 38414 578898
rect 37794 543218 37826 543454
rect 38062 543218 38146 543454
rect 38382 543218 38414 543454
rect 37794 543134 38414 543218
rect 37794 542898 37826 543134
rect 38062 542898 38146 543134
rect 38382 542898 38414 543134
rect 27834 533258 27866 533494
rect 28102 533258 28186 533494
rect 28422 533258 28454 533494
rect 27834 533174 28454 533258
rect 27834 532938 27866 533174
rect 28102 532938 28186 533174
rect 28422 532938 28454 533174
rect 27834 497494 28454 532938
rect 34208 507454 34528 507486
rect 34208 507218 34250 507454
rect 34486 507218 34528 507454
rect 34208 507134 34528 507218
rect 34208 506898 34250 507134
rect 34486 506898 34528 507134
rect 34208 506866 34528 506898
rect 37794 507454 38414 542898
rect 37794 507218 37826 507454
rect 38062 507218 38146 507454
rect 38382 507218 38414 507454
rect 37794 507134 38414 507218
rect 37794 506898 37826 507134
rect 38062 506898 38146 507134
rect 38382 506898 38414 507134
rect 27834 497258 27866 497494
rect 28102 497258 28186 497494
rect 28422 497258 28454 497494
rect 27834 497174 28454 497258
rect 27834 496938 27866 497174
rect 28102 496938 28186 497174
rect 28422 496938 28454 497174
rect 27834 461494 28454 496938
rect 34208 471454 34528 471486
rect 34208 471218 34250 471454
rect 34486 471218 34528 471454
rect 34208 471134 34528 471218
rect 34208 470898 34250 471134
rect 34486 470898 34528 471134
rect 34208 470866 34528 470898
rect 37794 471454 38414 506898
rect 37794 471218 37826 471454
rect 38062 471218 38146 471454
rect 38382 471218 38414 471454
rect 37794 471134 38414 471218
rect 37794 470898 37826 471134
rect 38062 470898 38146 471134
rect 38382 470898 38414 471134
rect 27834 461258 27866 461494
rect 28102 461258 28186 461494
rect 28422 461258 28454 461494
rect 27834 461174 28454 461258
rect 27834 460938 27866 461174
rect 28102 460938 28186 461174
rect 28422 460938 28454 461174
rect 27834 425494 28454 460938
rect 27834 425258 27866 425494
rect 28102 425258 28186 425494
rect 28422 425258 28454 425494
rect 27834 425174 28454 425258
rect 27834 424938 27866 425174
rect 28102 424938 28186 425174
rect 28422 424938 28454 425174
rect 27834 389494 28454 424938
rect 27834 389258 27866 389494
rect 28102 389258 28186 389494
rect 28422 389258 28454 389494
rect 27834 389174 28454 389258
rect 27834 388938 27866 389174
rect 28102 388938 28186 389174
rect 28422 388938 28454 389174
rect 27834 353494 28454 388938
rect 27834 353258 27866 353494
rect 28102 353258 28186 353494
rect 28422 353258 28454 353494
rect 27834 353174 28454 353258
rect 27834 352938 27866 353174
rect 28102 352938 28186 353174
rect 28422 352938 28454 353174
rect 27834 317494 28454 352938
rect 27834 317258 27866 317494
rect 28102 317258 28186 317494
rect 28422 317258 28454 317494
rect 27834 317174 28454 317258
rect 27834 316938 27866 317174
rect 28102 316938 28186 317174
rect 28422 316938 28454 317174
rect 27834 281494 28454 316938
rect 37794 435454 38414 470898
rect 37794 435218 37826 435454
rect 38062 435218 38146 435454
rect 38382 435218 38414 435454
rect 37794 435134 38414 435218
rect 37794 434898 37826 435134
rect 38062 434898 38146 435134
rect 38382 434898 38414 435134
rect 37794 399454 38414 434898
rect 37794 399218 37826 399454
rect 38062 399218 38146 399454
rect 38382 399218 38414 399454
rect 37794 399134 38414 399218
rect 37794 398898 37826 399134
rect 38062 398898 38146 399134
rect 38382 398898 38414 399134
rect 37794 363454 38414 398898
rect 37794 363218 37826 363454
rect 38062 363218 38146 363454
rect 38382 363218 38414 363454
rect 37794 363134 38414 363218
rect 37794 362898 37826 363134
rect 38062 362898 38146 363134
rect 38382 362898 38414 363134
rect 37794 327454 38414 362898
rect 37794 327218 37826 327454
rect 38062 327218 38146 327454
rect 38382 327218 38414 327454
rect 37794 327134 38414 327218
rect 37794 326898 37826 327134
rect 38062 326898 38146 327134
rect 38382 326898 38414 327134
rect 34208 291454 34528 291486
rect 34208 291218 34250 291454
rect 34486 291218 34528 291454
rect 34208 291134 34528 291218
rect 34208 290898 34250 291134
rect 34486 290898 34528 291134
rect 34208 290866 34528 290898
rect 37794 291454 38414 326898
rect 37794 291218 37826 291454
rect 38062 291218 38146 291454
rect 38382 291218 38414 291454
rect 37794 291134 38414 291218
rect 37794 290898 37826 291134
rect 38062 290898 38146 291134
rect 38382 290898 38414 291134
rect 27834 281258 27866 281494
rect 28102 281258 28186 281494
rect 28422 281258 28454 281494
rect 27834 281174 28454 281258
rect 27834 280938 27866 281174
rect 28102 280938 28186 281174
rect 28422 280938 28454 281174
rect 27834 245494 28454 280938
rect 34208 255454 34528 255486
rect 34208 255218 34250 255454
rect 34486 255218 34528 255454
rect 34208 255134 34528 255218
rect 34208 254898 34250 255134
rect 34486 254898 34528 255134
rect 34208 254866 34528 254898
rect 37794 255454 38414 290898
rect 37794 255218 37826 255454
rect 38062 255218 38146 255454
rect 38382 255218 38414 255454
rect 37794 255134 38414 255218
rect 37794 254898 37826 255134
rect 38062 254898 38146 255134
rect 38382 254898 38414 255134
rect 27834 245258 27866 245494
rect 28102 245258 28186 245494
rect 28422 245258 28454 245494
rect 27834 245174 28454 245258
rect 27834 244938 27866 245174
rect 28102 244938 28186 245174
rect 28422 244938 28454 245174
rect 27834 209494 28454 244938
rect 34208 219454 34528 219486
rect 34208 219218 34250 219454
rect 34486 219218 34528 219454
rect 34208 219134 34528 219218
rect 34208 218898 34250 219134
rect 34486 218898 34528 219134
rect 34208 218866 34528 218898
rect 37794 219454 38414 254898
rect 37794 219218 37826 219454
rect 38062 219218 38146 219454
rect 38382 219218 38414 219454
rect 37794 219134 38414 219218
rect 37794 218898 37826 219134
rect 38062 218898 38146 219134
rect 38382 218898 38414 219134
rect 27834 209258 27866 209494
rect 28102 209258 28186 209494
rect 28422 209258 28454 209494
rect 27834 209174 28454 209258
rect 27834 208938 27866 209174
rect 28102 208938 28186 209174
rect 28422 208938 28454 209174
rect 27834 173494 28454 208938
rect 34208 183454 34528 183486
rect 34208 183218 34250 183454
rect 34486 183218 34528 183454
rect 34208 183134 34528 183218
rect 34208 182898 34250 183134
rect 34486 182898 34528 183134
rect 34208 182866 34528 182898
rect 37794 183454 38414 218898
rect 37794 183218 37826 183454
rect 38062 183218 38146 183454
rect 38382 183218 38414 183454
rect 37794 183134 38414 183218
rect 37794 182898 37826 183134
rect 38062 182898 38146 183134
rect 38382 182898 38414 183134
rect 27834 173258 27866 173494
rect 28102 173258 28186 173494
rect 28422 173258 28454 173494
rect 27834 173174 28454 173258
rect 27834 172938 27866 173174
rect 28102 172938 28186 173174
rect 28422 172938 28454 173174
rect 27834 137494 28454 172938
rect 27834 137258 27866 137494
rect 28102 137258 28186 137494
rect 28422 137258 28454 137494
rect 27834 137174 28454 137258
rect 27834 136938 27866 137174
rect 28102 136938 28186 137174
rect 28422 136938 28454 137174
rect 27834 133820 28454 136938
rect 37794 147454 38414 182898
rect 37794 147218 37826 147454
rect 38062 147218 38146 147454
rect 38382 147218 38414 147454
rect 37794 147134 38414 147218
rect 37794 146898 37826 147134
rect 38062 146898 38146 147134
rect 38382 146898 38414 147134
rect 24114 133538 24146 133774
rect 24382 133538 24466 133774
rect 24702 133538 24734 133774
rect 24114 133454 24734 133538
rect 24114 133218 24146 133454
rect 24382 133218 24466 133454
rect 24702 133218 24734 133454
rect 24114 97774 24734 133218
rect 37794 133057 38414 146898
rect 41514 705798 42134 711590
rect 41514 705562 41546 705798
rect 41782 705562 41866 705798
rect 42102 705562 42134 705798
rect 41514 705478 42134 705562
rect 41514 705242 41546 705478
rect 41782 705242 41866 705478
rect 42102 705242 42134 705478
rect 41514 691174 42134 705242
rect 41514 690938 41546 691174
rect 41782 690938 41866 691174
rect 42102 690938 42134 691174
rect 41514 690854 42134 690938
rect 41514 690618 41546 690854
rect 41782 690618 41866 690854
rect 42102 690618 42134 690854
rect 41514 655174 42134 690618
rect 41514 654938 41546 655174
rect 41782 654938 41866 655174
rect 42102 654938 42134 655174
rect 41514 654854 42134 654938
rect 41514 654618 41546 654854
rect 41782 654618 41866 654854
rect 42102 654618 42134 654854
rect 41514 619174 42134 654618
rect 41514 618938 41546 619174
rect 41782 618938 41866 619174
rect 42102 618938 42134 619174
rect 41514 618854 42134 618938
rect 41514 618618 41546 618854
rect 41782 618618 41866 618854
rect 42102 618618 42134 618854
rect 41514 583174 42134 618618
rect 41514 582938 41546 583174
rect 41782 582938 41866 583174
rect 42102 582938 42134 583174
rect 41514 582854 42134 582938
rect 41514 582618 41546 582854
rect 41782 582618 41866 582854
rect 42102 582618 42134 582854
rect 41514 547174 42134 582618
rect 41514 546938 41546 547174
rect 41782 546938 41866 547174
rect 42102 546938 42134 547174
rect 41514 546854 42134 546938
rect 41514 546618 41546 546854
rect 41782 546618 41866 546854
rect 42102 546618 42134 546854
rect 41514 511174 42134 546618
rect 41514 510938 41546 511174
rect 41782 510938 41866 511174
rect 42102 510938 42134 511174
rect 41514 510854 42134 510938
rect 41514 510618 41546 510854
rect 41782 510618 41866 510854
rect 42102 510618 42134 510854
rect 41514 475174 42134 510618
rect 41514 474938 41546 475174
rect 41782 474938 41866 475174
rect 42102 474938 42134 475174
rect 41514 474854 42134 474938
rect 41514 474618 41546 474854
rect 41782 474618 41866 474854
rect 42102 474618 42134 474854
rect 41514 439174 42134 474618
rect 41514 438938 41546 439174
rect 41782 438938 41866 439174
rect 42102 438938 42134 439174
rect 41514 438854 42134 438938
rect 41514 438618 41546 438854
rect 41782 438618 41866 438854
rect 42102 438618 42134 438854
rect 41514 403174 42134 438618
rect 41514 402938 41546 403174
rect 41782 402938 41866 403174
rect 42102 402938 42134 403174
rect 41514 402854 42134 402938
rect 41514 402618 41546 402854
rect 41782 402618 41866 402854
rect 42102 402618 42134 402854
rect 41514 367174 42134 402618
rect 41514 366938 41546 367174
rect 41782 366938 41866 367174
rect 42102 366938 42134 367174
rect 41514 366854 42134 366938
rect 41514 366618 41546 366854
rect 41782 366618 41866 366854
rect 42102 366618 42134 366854
rect 41514 331174 42134 366618
rect 41514 330938 41546 331174
rect 41782 330938 41866 331174
rect 42102 330938 42134 331174
rect 41514 330854 42134 330938
rect 41514 330618 41546 330854
rect 41782 330618 41866 330854
rect 42102 330618 42134 330854
rect 41514 295174 42134 330618
rect 41514 294938 41546 295174
rect 41782 294938 41866 295174
rect 42102 294938 42134 295174
rect 41514 294854 42134 294938
rect 41514 294618 41546 294854
rect 41782 294618 41866 294854
rect 42102 294618 42134 294854
rect 41514 259174 42134 294618
rect 41514 258938 41546 259174
rect 41782 258938 41866 259174
rect 42102 258938 42134 259174
rect 41514 258854 42134 258938
rect 41514 258618 41546 258854
rect 41782 258618 41866 258854
rect 42102 258618 42134 258854
rect 41514 223174 42134 258618
rect 41514 222938 41546 223174
rect 41782 222938 41866 223174
rect 42102 222938 42134 223174
rect 41514 222854 42134 222938
rect 41514 222618 41546 222854
rect 41782 222618 41866 222854
rect 42102 222618 42134 222854
rect 41514 187174 42134 222618
rect 41514 186938 41546 187174
rect 41782 186938 41866 187174
rect 42102 186938 42134 187174
rect 41514 186854 42134 186938
rect 41514 186618 41546 186854
rect 41782 186618 41866 186854
rect 42102 186618 42134 186854
rect 41514 151174 42134 186618
rect 41514 150938 41546 151174
rect 41782 150938 41866 151174
rect 42102 150938 42134 151174
rect 41514 150854 42134 150938
rect 41514 150618 41546 150854
rect 41782 150618 41866 150854
rect 42102 150618 42134 150854
rect 41514 133057 42134 150618
rect 45234 706758 45854 711590
rect 45234 706522 45266 706758
rect 45502 706522 45586 706758
rect 45822 706522 45854 706758
rect 45234 706438 45854 706522
rect 45234 706202 45266 706438
rect 45502 706202 45586 706438
rect 45822 706202 45854 706438
rect 45234 694894 45854 706202
rect 45234 694658 45266 694894
rect 45502 694658 45586 694894
rect 45822 694658 45854 694894
rect 45234 694574 45854 694658
rect 45234 694338 45266 694574
rect 45502 694338 45586 694574
rect 45822 694338 45854 694574
rect 45234 658894 45854 694338
rect 45234 658658 45266 658894
rect 45502 658658 45586 658894
rect 45822 658658 45854 658894
rect 45234 658574 45854 658658
rect 45234 658338 45266 658574
rect 45502 658338 45586 658574
rect 45822 658338 45854 658574
rect 45234 622894 45854 658338
rect 45234 622658 45266 622894
rect 45502 622658 45586 622894
rect 45822 622658 45854 622894
rect 45234 622574 45854 622658
rect 45234 622338 45266 622574
rect 45502 622338 45586 622574
rect 45822 622338 45854 622574
rect 45234 586894 45854 622338
rect 48954 707718 49574 711590
rect 48954 707482 48986 707718
rect 49222 707482 49306 707718
rect 49542 707482 49574 707718
rect 48954 707398 49574 707482
rect 48954 707162 48986 707398
rect 49222 707162 49306 707398
rect 49542 707162 49574 707398
rect 48954 698614 49574 707162
rect 48954 698378 48986 698614
rect 49222 698378 49306 698614
rect 49542 698378 49574 698614
rect 48954 698294 49574 698378
rect 48954 698058 48986 698294
rect 49222 698058 49306 698294
rect 49542 698058 49574 698294
rect 48954 662614 49574 698058
rect 48954 662378 48986 662614
rect 49222 662378 49306 662614
rect 49542 662378 49574 662614
rect 48954 662294 49574 662378
rect 48954 662058 48986 662294
rect 49222 662058 49306 662294
rect 49542 662058 49574 662294
rect 48954 626614 49574 662058
rect 48954 626378 48986 626614
rect 49222 626378 49306 626614
rect 49542 626378 49574 626614
rect 48954 626294 49574 626378
rect 48954 626058 48986 626294
rect 49222 626058 49306 626294
rect 49542 626058 49574 626294
rect 48954 599868 49574 626058
rect 52674 708678 53294 711590
rect 52674 708442 52706 708678
rect 52942 708442 53026 708678
rect 53262 708442 53294 708678
rect 52674 708358 53294 708442
rect 52674 708122 52706 708358
rect 52942 708122 53026 708358
rect 53262 708122 53294 708358
rect 52674 666334 53294 708122
rect 52674 666098 52706 666334
rect 52942 666098 53026 666334
rect 53262 666098 53294 666334
rect 52674 666014 53294 666098
rect 52674 665778 52706 666014
rect 52942 665778 53026 666014
rect 53262 665778 53294 666014
rect 52674 630334 53294 665778
rect 52674 630098 52706 630334
rect 52942 630098 53026 630334
rect 53262 630098 53294 630334
rect 52674 630014 53294 630098
rect 52674 629778 52706 630014
rect 52942 629778 53026 630014
rect 53262 629778 53294 630014
rect 45234 586658 45266 586894
rect 45502 586658 45586 586894
rect 45822 586658 45854 586894
rect 45234 586574 45854 586658
rect 45234 586338 45266 586574
rect 45502 586338 45586 586574
rect 45822 586338 45854 586574
rect 45234 550894 45854 586338
rect 52674 594334 53294 629778
rect 52674 594098 52706 594334
rect 52942 594098 53026 594334
rect 53262 594098 53294 594334
rect 52674 594014 53294 594098
rect 52674 593778 52706 594014
rect 52942 593778 53026 594014
rect 53262 593778 53294 594014
rect 49568 583174 49888 583206
rect 49568 582938 49610 583174
rect 49846 582938 49888 583174
rect 49568 582854 49888 582938
rect 49568 582618 49610 582854
rect 49846 582618 49888 582854
rect 49568 582586 49888 582618
rect 45234 550658 45266 550894
rect 45502 550658 45586 550894
rect 45822 550658 45854 550894
rect 45234 550574 45854 550658
rect 45234 550338 45266 550574
rect 45502 550338 45586 550574
rect 45822 550338 45854 550574
rect 45234 514894 45854 550338
rect 52674 558334 53294 593778
rect 52674 558098 52706 558334
rect 52942 558098 53026 558334
rect 53262 558098 53294 558334
rect 52674 558014 53294 558098
rect 52674 557778 52706 558014
rect 52942 557778 53026 558014
rect 53262 557778 53294 558014
rect 49568 547174 49888 547206
rect 49568 546938 49610 547174
rect 49846 546938 49888 547174
rect 49568 546854 49888 546938
rect 49568 546618 49610 546854
rect 49846 546618 49888 546854
rect 49568 546586 49888 546618
rect 45234 514658 45266 514894
rect 45502 514658 45586 514894
rect 45822 514658 45854 514894
rect 45234 514574 45854 514658
rect 45234 514338 45266 514574
rect 45502 514338 45586 514574
rect 45822 514338 45854 514574
rect 45234 478894 45854 514338
rect 52674 522334 53294 557778
rect 52674 522098 52706 522334
rect 52942 522098 53026 522334
rect 53262 522098 53294 522334
rect 52674 522014 53294 522098
rect 52674 521778 52706 522014
rect 52942 521778 53026 522014
rect 53262 521778 53294 522014
rect 49568 511174 49888 511206
rect 49568 510938 49610 511174
rect 49846 510938 49888 511174
rect 49568 510854 49888 510938
rect 49568 510618 49610 510854
rect 49846 510618 49888 510854
rect 49568 510586 49888 510618
rect 45234 478658 45266 478894
rect 45502 478658 45586 478894
rect 45822 478658 45854 478894
rect 45234 478574 45854 478658
rect 45234 478338 45266 478574
rect 45502 478338 45586 478574
rect 45822 478338 45854 478574
rect 45234 442894 45854 478338
rect 52674 486334 53294 521778
rect 52674 486098 52706 486334
rect 52942 486098 53026 486334
rect 53262 486098 53294 486334
rect 52674 486014 53294 486098
rect 52674 485778 52706 486014
rect 52942 485778 53026 486014
rect 53262 485778 53294 486014
rect 49568 475174 49888 475206
rect 49568 474938 49610 475174
rect 49846 474938 49888 475174
rect 49568 474854 49888 474938
rect 49568 474618 49610 474854
rect 49846 474618 49888 474854
rect 49568 474586 49888 474618
rect 45234 442658 45266 442894
rect 45502 442658 45586 442894
rect 45822 442658 45854 442894
rect 45234 442574 45854 442658
rect 45234 442338 45266 442574
rect 45502 442338 45586 442574
rect 45822 442338 45854 442574
rect 45234 406894 45854 442338
rect 52674 450334 53294 485778
rect 52674 450098 52706 450334
rect 52942 450098 53026 450334
rect 53262 450098 53294 450334
rect 52674 450014 53294 450098
rect 52674 449778 52706 450014
rect 52942 449778 53026 450014
rect 53262 449778 53294 450014
rect 45234 406658 45266 406894
rect 45502 406658 45586 406894
rect 45822 406658 45854 406894
rect 45234 406574 45854 406658
rect 45234 406338 45266 406574
rect 45502 406338 45586 406574
rect 45822 406338 45854 406574
rect 45234 370894 45854 406338
rect 45234 370658 45266 370894
rect 45502 370658 45586 370894
rect 45822 370658 45854 370894
rect 45234 370574 45854 370658
rect 45234 370338 45266 370574
rect 45502 370338 45586 370574
rect 45822 370338 45854 370574
rect 45234 334894 45854 370338
rect 45234 334658 45266 334894
rect 45502 334658 45586 334894
rect 45822 334658 45854 334894
rect 45234 334574 45854 334658
rect 45234 334338 45266 334574
rect 45502 334338 45586 334574
rect 45822 334338 45854 334574
rect 45234 298894 45854 334338
rect 48954 410614 49574 440068
rect 48954 410378 48986 410614
rect 49222 410378 49306 410614
rect 49542 410378 49574 410614
rect 48954 410294 49574 410378
rect 48954 410058 48986 410294
rect 49222 410058 49306 410294
rect 49542 410058 49574 410294
rect 48954 374614 49574 410058
rect 48954 374378 48986 374614
rect 49222 374378 49306 374614
rect 49542 374378 49574 374614
rect 48954 374294 49574 374378
rect 48954 374058 48986 374294
rect 49222 374058 49306 374294
rect 49542 374058 49574 374294
rect 48954 338614 49574 374058
rect 48954 338378 48986 338614
rect 49222 338378 49306 338614
rect 49542 338378 49574 338614
rect 48954 338294 49574 338378
rect 48954 338058 48986 338294
rect 49222 338058 49306 338294
rect 49542 338058 49574 338294
rect 48954 323676 49574 338058
rect 52674 414334 53294 449778
rect 52674 414098 52706 414334
rect 52942 414098 53026 414334
rect 53262 414098 53294 414334
rect 52674 414014 53294 414098
rect 52674 413778 52706 414014
rect 52942 413778 53026 414014
rect 53262 413778 53294 414014
rect 52674 378334 53294 413778
rect 52674 378098 52706 378334
rect 52942 378098 53026 378334
rect 53262 378098 53294 378334
rect 52674 378014 53294 378098
rect 52674 377778 52706 378014
rect 52942 377778 53026 378014
rect 53262 377778 53294 378014
rect 52674 342334 53294 377778
rect 52674 342098 52706 342334
rect 52942 342098 53026 342334
rect 53262 342098 53294 342334
rect 52674 342014 53294 342098
rect 52674 341778 52706 342014
rect 52942 341778 53026 342014
rect 53262 341778 53294 342014
rect 45234 298658 45266 298894
rect 45502 298658 45586 298894
rect 45822 298658 45854 298894
rect 45234 298574 45854 298658
rect 45234 298338 45266 298574
rect 45502 298338 45586 298574
rect 45822 298338 45854 298574
rect 45234 262894 45854 298338
rect 52674 306334 53294 341778
rect 52674 306098 52706 306334
rect 52942 306098 53026 306334
rect 53262 306098 53294 306334
rect 52674 306014 53294 306098
rect 52674 305778 52706 306014
rect 52942 305778 53026 306014
rect 53262 305778 53294 306014
rect 49568 295174 49888 295206
rect 49568 294938 49610 295174
rect 49846 294938 49888 295174
rect 49568 294854 49888 294938
rect 49568 294618 49610 294854
rect 49846 294618 49888 294854
rect 49568 294586 49888 294618
rect 45234 262658 45266 262894
rect 45502 262658 45586 262894
rect 45822 262658 45854 262894
rect 45234 262574 45854 262658
rect 45234 262338 45266 262574
rect 45502 262338 45586 262574
rect 45822 262338 45854 262574
rect 45234 226894 45854 262338
rect 52674 270334 53294 305778
rect 52674 270098 52706 270334
rect 52942 270098 53026 270334
rect 53262 270098 53294 270334
rect 52674 270014 53294 270098
rect 52674 269778 52706 270014
rect 52942 269778 53026 270014
rect 53262 269778 53294 270014
rect 49568 259174 49888 259206
rect 49568 258938 49610 259174
rect 49846 258938 49888 259174
rect 49568 258854 49888 258938
rect 49568 258618 49610 258854
rect 49846 258618 49888 258854
rect 49568 258586 49888 258618
rect 45234 226658 45266 226894
rect 45502 226658 45586 226894
rect 45822 226658 45854 226894
rect 45234 226574 45854 226658
rect 45234 226338 45266 226574
rect 45502 226338 45586 226574
rect 45822 226338 45854 226574
rect 45234 190894 45854 226338
rect 52674 234334 53294 269778
rect 52674 234098 52706 234334
rect 52942 234098 53026 234334
rect 53262 234098 53294 234334
rect 52674 234014 53294 234098
rect 52674 233778 52706 234014
rect 52942 233778 53026 234014
rect 53262 233778 53294 234014
rect 49568 223174 49888 223206
rect 49568 222938 49610 223174
rect 49846 222938 49888 223174
rect 49568 222854 49888 222938
rect 49568 222618 49610 222854
rect 49846 222618 49888 222854
rect 49568 222586 49888 222618
rect 45234 190658 45266 190894
rect 45502 190658 45586 190894
rect 45822 190658 45854 190894
rect 45234 190574 45854 190658
rect 45234 190338 45266 190574
rect 45502 190338 45586 190574
rect 45822 190338 45854 190574
rect 45234 154894 45854 190338
rect 52674 198334 53294 233778
rect 52674 198098 52706 198334
rect 52942 198098 53026 198334
rect 53262 198098 53294 198334
rect 52674 198014 53294 198098
rect 52674 197778 52706 198014
rect 52942 197778 53026 198014
rect 53262 197778 53294 198014
rect 49568 187174 49888 187206
rect 49568 186938 49610 187174
rect 49846 186938 49888 187174
rect 49568 186854 49888 186938
rect 49568 186618 49610 186854
rect 49846 186618 49888 186854
rect 49568 186586 49888 186618
rect 45234 154658 45266 154894
rect 45502 154658 45586 154894
rect 45822 154658 45854 154894
rect 45234 154574 45854 154658
rect 45234 154338 45266 154574
rect 45502 154338 45586 154574
rect 45822 154338 45854 154574
rect 45234 133057 45854 154338
rect 52674 162334 53294 197778
rect 52674 162098 52706 162334
rect 52942 162098 53026 162334
rect 53262 162098 53294 162334
rect 52674 162014 53294 162098
rect 52674 161778 52706 162014
rect 52942 161778 53026 162014
rect 53262 161778 53294 162014
rect 52674 133057 53294 161778
rect 56394 709638 57014 711590
rect 56394 709402 56426 709638
rect 56662 709402 56746 709638
rect 56982 709402 57014 709638
rect 56394 709318 57014 709402
rect 56394 709082 56426 709318
rect 56662 709082 56746 709318
rect 56982 709082 57014 709318
rect 56394 670054 57014 709082
rect 56394 669818 56426 670054
rect 56662 669818 56746 670054
rect 56982 669818 57014 670054
rect 56394 669734 57014 669818
rect 56394 669498 56426 669734
rect 56662 669498 56746 669734
rect 56982 669498 57014 669734
rect 56394 634054 57014 669498
rect 56394 633818 56426 634054
rect 56662 633818 56746 634054
rect 56982 633818 57014 634054
rect 56394 633734 57014 633818
rect 56394 633498 56426 633734
rect 56662 633498 56746 633734
rect 56982 633498 57014 633734
rect 56394 598054 57014 633498
rect 56394 597818 56426 598054
rect 56662 597818 56746 598054
rect 56982 597818 57014 598054
rect 56394 597734 57014 597818
rect 56394 597498 56426 597734
rect 56662 597498 56746 597734
rect 56982 597498 57014 597734
rect 56394 562054 57014 597498
rect 56394 561818 56426 562054
rect 56662 561818 56746 562054
rect 56982 561818 57014 562054
rect 56394 561734 57014 561818
rect 56394 561498 56426 561734
rect 56662 561498 56746 561734
rect 56982 561498 57014 561734
rect 56394 526054 57014 561498
rect 56394 525818 56426 526054
rect 56662 525818 56746 526054
rect 56982 525818 57014 526054
rect 56394 525734 57014 525818
rect 56394 525498 56426 525734
rect 56662 525498 56746 525734
rect 56982 525498 57014 525734
rect 56394 490054 57014 525498
rect 56394 489818 56426 490054
rect 56662 489818 56746 490054
rect 56982 489818 57014 490054
rect 56394 489734 57014 489818
rect 56394 489498 56426 489734
rect 56662 489498 56746 489734
rect 56982 489498 57014 489734
rect 56394 454054 57014 489498
rect 56394 453818 56426 454054
rect 56662 453818 56746 454054
rect 56982 453818 57014 454054
rect 56394 453734 57014 453818
rect 56394 453498 56426 453734
rect 56662 453498 56746 453734
rect 56982 453498 57014 453734
rect 56394 418054 57014 453498
rect 56394 417818 56426 418054
rect 56662 417818 56746 418054
rect 56982 417818 57014 418054
rect 56394 417734 57014 417818
rect 56394 417498 56426 417734
rect 56662 417498 56746 417734
rect 56982 417498 57014 417734
rect 56394 382054 57014 417498
rect 56394 381818 56426 382054
rect 56662 381818 56746 382054
rect 56982 381818 57014 382054
rect 56394 381734 57014 381818
rect 56394 381498 56426 381734
rect 56662 381498 56746 381734
rect 56982 381498 57014 381734
rect 56394 346054 57014 381498
rect 56394 345818 56426 346054
rect 56662 345818 56746 346054
rect 56982 345818 57014 346054
rect 56394 345734 57014 345818
rect 56394 345498 56426 345734
rect 56662 345498 56746 345734
rect 56982 345498 57014 345734
rect 56394 310054 57014 345498
rect 56394 309818 56426 310054
rect 56662 309818 56746 310054
rect 56982 309818 57014 310054
rect 56394 309734 57014 309818
rect 56394 309498 56426 309734
rect 56662 309498 56746 309734
rect 56982 309498 57014 309734
rect 56394 274054 57014 309498
rect 56394 273818 56426 274054
rect 56662 273818 56746 274054
rect 56982 273818 57014 274054
rect 56394 273734 57014 273818
rect 56394 273498 56426 273734
rect 56662 273498 56746 273734
rect 56982 273498 57014 273734
rect 56394 238054 57014 273498
rect 56394 237818 56426 238054
rect 56662 237818 56746 238054
rect 56982 237818 57014 238054
rect 56394 237734 57014 237818
rect 56394 237498 56426 237734
rect 56662 237498 56746 237734
rect 56982 237498 57014 237734
rect 56394 202054 57014 237498
rect 56394 201818 56426 202054
rect 56662 201818 56746 202054
rect 56982 201818 57014 202054
rect 56394 201734 57014 201818
rect 56394 201498 56426 201734
rect 56662 201498 56746 201734
rect 56982 201498 57014 201734
rect 56394 166054 57014 201498
rect 56394 165818 56426 166054
rect 56662 165818 56746 166054
rect 56982 165818 57014 166054
rect 56394 165734 57014 165818
rect 56394 165498 56426 165734
rect 56662 165498 56746 165734
rect 56982 165498 57014 165734
rect 56394 133057 57014 165498
rect 60114 710598 60734 711590
rect 60114 710362 60146 710598
rect 60382 710362 60466 710598
rect 60702 710362 60734 710598
rect 60114 710278 60734 710362
rect 60114 710042 60146 710278
rect 60382 710042 60466 710278
rect 60702 710042 60734 710278
rect 60114 673774 60734 710042
rect 60114 673538 60146 673774
rect 60382 673538 60466 673774
rect 60702 673538 60734 673774
rect 60114 673454 60734 673538
rect 60114 673218 60146 673454
rect 60382 673218 60466 673454
rect 60702 673218 60734 673454
rect 60114 637774 60734 673218
rect 60114 637538 60146 637774
rect 60382 637538 60466 637774
rect 60702 637538 60734 637774
rect 60114 637454 60734 637538
rect 60114 637218 60146 637454
rect 60382 637218 60466 637454
rect 60702 637218 60734 637454
rect 60114 601774 60734 637218
rect 60114 601538 60146 601774
rect 60382 601538 60466 601774
rect 60702 601538 60734 601774
rect 60114 601454 60734 601538
rect 60114 601218 60146 601454
rect 60382 601218 60466 601454
rect 60702 601218 60734 601454
rect 60114 565774 60734 601218
rect 63834 711558 64454 711590
rect 63834 711322 63866 711558
rect 64102 711322 64186 711558
rect 64422 711322 64454 711558
rect 63834 711238 64454 711322
rect 63834 711002 63866 711238
rect 64102 711002 64186 711238
rect 64422 711002 64454 711238
rect 63834 677494 64454 711002
rect 63834 677258 63866 677494
rect 64102 677258 64186 677494
rect 64422 677258 64454 677494
rect 63834 677174 64454 677258
rect 63834 676938 63866 677174
rect 64102 676938 64186 677174
rect 64422 676938 64454 677174
rect 63834 641494 64454 676938
rect 63834 641258 63866 641494
rect 64102 641258 64186 641494
rect 64422 641258 64454 641494
rect 63834 641174 64454 641258
rect 63834 640938 63866 641174
rect 64102 640938 64186 641174
rect 64422 640938 64454 641174
rect 63834 605494 64454 640938
rect 63834 605258 63866 605494
rect 64102 605258 64186 605494
rect 64422 605258 64454 605494
rect 63834 605174 64454 605258
rect 63834 604938 63866 605174
rect 64102 604938 64186 605174
rect 64422 604938 64454 605174
rect 63834 595705 64454 604938
rect 73794 704838 74414 711590
rect 73794 704602 73826 704838
rect 74062 704602 74146 704838
rect 74382 704602 74414 704838
rect 73794 704518 74414 704602
rect 73794 704282 73826 704518
rect 74062 704282 74146 704518
rect 74382 704282 74414 704518
rect 73794 687454 74414 704282
rect 73794 687218 73826 687454
rect 74062 687218 74146 687454
rect 74382 687218 74414 687454
rect 73794 687134 74414 687218
rect 73794 686898 73826 687134
rect 74062 686898 74146 687134
rect 74382 686898 74414 687134
rect 73794 651454 74414 686898
rect 73794 651218 73826 651454
rect 74062 651218 74146 651454
rect 74382 651218 74414 651454
rect 73794 651134 74414 651218
rect 73794 650898 73826 651134
rect 74062 650898 74146 651134
rect 74382 650898 74414 651134
rect 73794 615454 74414 650898
rect 73794 615218 73826 615454
rect 74062 615218 74146 615454
rect 74382 615218 74414 615454
rect 73794 615134 74414 615218
rect 73794 614898 73826 615134
rect 74062 614898 74146 615134
rect 74382 614898 74414 615134
rect 73794 595705 74414 614898
rect 77514 705798 78134 711590
rect 77514 705562 77546 705798
rect 77782 705562 77866 705798
rect 78102 705562 78134 705798
rect 77514 705478 78134 705562
rect 77514 705242 77546 705478
rect 77782 705242 77866 705478
rect 78102 705242 78134 705478
rect 77514 691174 78134 705242
rect 77514 690938 77546 691174
rect 77782 690938 77866 691174
rect 78102 690938 78134 691174
rect 77514 690854 78134 690938
rect 77514 690618 77546 690854
rect 77782 690618 77866 690854
rect 78102 690618 78134 690854
rect 77514 655174 78134 690618
rect 77514 654938 77546 655174
rect 77782 654938 77866 655174
rect 78102 654938 78134 655174
rect 77514 654854 78134 654938
rect 77514 654618 77546 654854
rect 77782 654618 77866 654854
rect 78102 654618 78134 654854
rect 77514 619174 78134 654618
rect 77514 618938 77546 619174
rect 77782 618938 77866 619174
rect 78102 618938 78134 619174
rect 77514 618854 78134 618938
rect 77514 618618 77546 618854
rect 77782 618618 77866 618854
rect 78102 618618 78134 618854
rect 77514 595705 78134 618618
rect 81234 706758 81854 711590
rect 81234 706522 81266 706758
rect 81502 706522 81586 706758
rect 81822 706522 81854 706758
rect 81234 706438 81854 706522
rect 81234 706202 81266 706438
rect 81502 706202 81586 706438
rect 81822 706202 81854 706438
rect 81234 694894 81854 706202
rect 81234 694658 81266 694894
rect 81502 694658 81586 694894
rect 81822 694658 81854 694894
rect 81234 694574 81854 694658
rect 81234 694338 81266 694574
rect 81502 694338 81586 694574
rect 81822 694338 81854 694574
rect 81234 658894 81854 694338
rect 81234 658658 81266 658894
rect 81502 658658 81586 658894
rect 81822 658658 81854 658894
rect 81234 658574 81854 658658
rect 81234 658338 81266 658574
rect 81502 658338 81586 658574
rect 81822 658338 81854 658574
rect 81234 622894 81854 658338
rect 81234 622658 81266 622894
rect 81502 622658 81586 622894
rect 81822 622658 81854 622894
rect 81234 622574 81854 622658
rect 81234 622338 81266 622574
rect 81502 622338 81586 622574
rect 81822 622338 81854 622574
rect 81234 595705 81854 622338
rect 84954 707718 85574 711590
rect 84954 707482 84986 707718
rect 85222 707482 85306 707718
rect 85542 707482 85574 707718
rect 84954 707398 85574 707482
rect 84954 707162 84986 707398
rect 85222 707162 85306 707398
rect 85542 707162 85574 707398
rect 84954 698614 85574 707162
rect 84954 698378 84986 698614
rect 85222 698378 85306 698614
rect 85542 698378 85574 698614
rect 84954 698294 85574 698378
rect 84954 698058 84986 698294
rect 85222 698058 85306 698294
rect 85542 698058 85574 698294
rect 84954 662614 85574 698058
rect 84954 662378 84986 662614
rect 85222 662378 85306 662614
rect 85542 662378 85574 662614
rect 84954 662294 85574 662378
rect 84954 662058 84986 662294
rect 85222 662058 85306 662294
rect 85542 662058 85574 662294
rect 84954 626614 85574 662058
rect 84954 626378 84986 626614
rect 85222 626378 85306 626614
rect 85542 626378 85574 626614
rect 84954 626294 85574 626378
rect 84954 626058 84986 626294
rect 85222 626058 85306 626294
rect 85542 626058 85574 626294
rect 84954 595705 85574 626058
rect 88674 708678 89294 711590
rect 88674 708442 88706 708678
rect 88942 708442 89026 708678
rect 89262 708442 89294 708678
rect 88674 708358 89294 708442
rect 88674 708122 88706 708358
rect 88942 708122 89026 708358
rect 89262 708122 89294 708358
rect 88674 666334 89294 708122
rect 88674 666098 88706 666334
rect 88942 666098 89026 666334
rect 89262 666098 89294 666334
rect 88674 666014 89294 666098
rect 88674 665778 88706 666014
rect 88942 665778 89026 666014
rect 89262 665778 89294 666014
rect 88674 630334 89294 665778
rect 88674 630098 88706 630334
rect 88942 630098 89026 630334
rect 89262 630098 89294 630334
rect 88674 630014 89294 630098
rect 88674 629778 88706 630014
rect 88942 629778 89026 630014
rect 89262 629778 89294 630014
rect 88674 595705 89294 629778
rect 92394 709638 93014 711590
rect 92394 709402 92426 709638
rect 92662 709402 92746 709638
rect 92982 709402 93014 709638
rect 92394 709318 93014 709402
rect 92394 709082 92426 709318
rect 92662 709082 92746 709318
rect 92982 709082 93014 709318
rect 92394 670054 93014 709082
rect 92394 669818 92426 670054
rect 92662 669818 92746 670054
rect 92982 669818 93014 670054
rect 92394 669734 93014 669818
rect 92394 669498 92426 669734
rect 92662 669498 92746 669734
rect 92982 669498 93014 669734
rect 92394 634054 93014 669498
rect 92394 633818 92426 634054
rect 92662 633818 92746 634054
rect 92982 633818 93014 634054
rect 92394 633734 93014 633818
rect 92394 633498 92426 633734
rect 92662 633498 92746 633734
rect 92982 633498 93014 633734
rect 92394 598054 93014 633498
rect 92394 597818 92426 598054
rect 92662 597818 92746 598054
rect 92982 597818 93014 598054
rect 92394 597734 93014 597818
rect 92394 597498 92426 597734
rect 92662 597498 92746 597734
rect 92982 597498 93014 597734
rect 92394 595705 93014 597498
rect 96114 710598 96734 711590
rect 96114 710362 96146 710598
rect 96382 710362 96466 710598
rect 96702 710362 96734 710598
rect 96114 710278 96734 710362
rect 96114 710042 96146 710278
rect 96382 710042 96466 710278
rect 96702 710042 96734 710278
rect 96114 673774 96734 710042
rect 96114 673538 96146 673774
rect 96382 673538 96466 673774
rect 96702 673538 96734 673774
rect 96114 673454 96734 673538
rect 96114 673218 96146 673454
rect 96382 673218 96466 673454
rect 96702 673218 96734 673454
rect 96114 637774 96734 673218
rect 96114 637538 96146 637774
rect 96382 637538 96466 637774
rect 96702 637538 96734 637774
rect 96114 637454 96734 637538
rect 96114 637218 96146 637454
rect 96382 637218 96466 637454
rect 96702 637218 96734 637454
rect 96114 601774 96734 637218
rect 96114 601538 96146 601774
rect 96382 601538 96466 601774
rect 96702 601538 96734 601774
rect 96114 601454 96734 601538
rect 96114 601218 96146 601454
rect 96382 601218 96466 601454
rect 96702 601218 96734 601454
rect 96114 595705 96734 601218
rect 99834 711558 100454 711590
rect 99834 711322 99866 711558
rect 100102 711322 100186 711558
rect 100422 711322 100454 711558
rect 99834 711238 100454 711322
rect 99834 711002 99866 711238
rect 100102 711002 100186 711238
rect 100422 711002 100454 711238
rect 99834 677494 100454 711002
rect 99834 677258 99866 677494
rect 100102 677258 100186 677494
rect 100422 677258 100454 677494
rect 99834 677174 100454 677258
rect 99834 676938 99866 677174
rect 100102 676938 100186 677174
rect 100422 676938 100454 677174
rect 99834 641494 100454 676938
rect 99834 641258 99866 641494
rect 100102 641258 100186 641494
rect 100422 641258 100454 641494
rect 99834 641174 100454 641258
rect 99834 640938 99866 641174
rect 100102 640938 100186 641174
rect 100422 640938 100454 641174
rect 99834 605494 100454 640938
rect 99834 605258 99866 605494
rect 100102 605258 100186 605494
rect 100422 605258 100454 605494
rect 99834 605174 100454 605258
rect 99834 604938 99866 605174
rect 100102 604938 100186 605174
rect 100422 604938 100454 605174
rect 99834 595705 100454 604938
rect 109794 704838 110414 711590
rect 109794 704602 109826 704838
rect 110062 704602 110146 704838
rect 110382 704602 110414 704838
rect 109794 704518 110414 704602
rect 109794 704282 109826 704518
rect 110062 704282 110146 704518
rect 110382 704282 110414 704518
rect 109794 687454 110414 704282
rect 109794 687218 109826 687454
rect 110062 687218 110146 687454
rect 110382 687218 110414 687454
rect 109794 687134 110414 687218
rect 109794 686898 109826 687134
rect 110062 686898 110146 687134
rect 110382 686898 110414 687134
rect 109794 651454 110414 686898
rect 109794 651218 109826 651454
rect 110062 651218 110146 651454
rect 110382 651218 110414 651454
rect 109794 651134 110414 651218
rect 109794 650898 109826 651134
rect 110062 650898 110146 651134
rect 110382 650898 110414 651134
rect 109794 615454 110414 650898
rect 109794 615218 109826 615454
rect 110062 615218 110146 615454
rect 110382 615218 110414 615454
rect 109794 615134 110414 615218
rect 109794 614898 109826 615134
rect 110062 614898 110146 615134
rect 110382 614898 110414 615134
rect 80288 583174 80608 583206
rect 80288 582938 80330 583174
rect 80566 582938 80608 583174
rect 80288 582854 80608 582938
rect 80288 582618 80330 582854
rect 80566 582618 80608 582854
rect 80288 582586 80608 582618
rect 64928 579454 65248 579486
rect 64928 579218 64970 579454
rect 65206 579218 65248 579454
rect 64928 579134 65248 579218
rect 64928 578898 64970 579134
rect 65206 578898 65248 579134
rect 64928 578866 65248 578898
rect 95648 579454 95968 579486
rect 95648 579218 95690 579454
rect 95926 579218 95968 579454
rect 95648 579134 95968 579218
rect 95648 578898 95690 579134
rect 95926 578898 95968 579134
rect 95648 578866 95968 578898
rect 109794 579454 110414 614898
rect 109794 579218 109826 579454
rect 110062 579218 110146 579454
rect 110382 579218 110414 579454
rect 109794 579134 110414 579218
rect 109794 578898 109826 579134
rect 110062 578898 110146 579134
rect 110382 578898 110414 579134
rect 60114 565538 60146 565774
rect 60382 565538 60466 565774
rect 60702 565538 60734 565774
rect 60114 565454 60734 565538
rect 60114 565218 60146 565454
rect 60382 565218 60466 565454
rect 60702 565218 60734 565454
rect 60114 529774 60734 565218
rect 80288 547174 80608 547206
rect 80288 546938 80330 547174
rect 80566 546938 80608 547174
rect 80288 546854 80608 546938
rect 80288 546618 80330 546854
rect 80566 546618 80608 546854
rect 80288 546586 80608 546618
rect 64928 543454 65248 543486
rect 64928 543218 64970 543454
rect 65206 543218 65248 543454
rect 64928 543134 65248 543218
rect 64928 542898 64970 543134
rect 65206 542898 65248 543134
rect 64928 542866 65248 542898
rect 95648 543454 95968 543486
rect 95648 543218 95690 543454
rect 95926 543218 95968 543454
rect 95648 543134 95968 543218
rect 95648 542898 95690 543134
rect 95926 542898 95968 543134
rect 95648 542866 95968 542898
rect 109794 543454 110414 578898
rect 109794 543218 109826 543454
rect 110062 543218 110146 543454
rect 110382 543218 110414 543454
rect 109794 543134 110414 543218
rect 109794 542898 109826 543134
rect 110062 542898 110146 543134
rect 110382 542898 110414 543134
rect 60114 529538 60146 529774
rect 60382 529538 60466 529774
rect 60702 529538 60734 529774
rect 60114 529454 60734 529538
rect 60114 529218 60146 529454
rect 60382 529218 60466 529454
rect 60702 529218 60734 529454
rect 60114 493774 60734 529218
rect 80288 511174 80608 511206
rect 80288 510938 80330 511174
rect 80566 510938 80608 511174
rect 80288 510854 80608 510938
rect 80288 510618 80330 510854
rect 80566 510618 80608 510854
rect 80288 510586 80608 510618
rect 64928 507454 65248 507486
rect 64928 507218 64970 507454
rect 65206 507218 65248 507454
rect 64928 507134 65248 507218
rect 64928 506898 64970 507134
rect 65206 506898 65248 507134
rect 64928 506866 65248 506898
rect 95648 507454 95968 507486
rect 95648 507218 95690 507454
rect 95926 507218 95968 507454
rect 95648 507134 95968 507218
rect 95648 506898 95690 507134
rect 95926 506898 95968 507134
rect 95648 506866 95968 506898
rect 109794 507454 110414 542898
rect 109794 507218 109826 507454
rect 110062 507218 110146 507454
rect 110382 507218 110414 507454
rect 109794 507134 110414 507218
rect 109794 506898 109826 507134
rect 110062 506898 110146 507134
rect 110382 506898 110414 507134
rect 60114 493538 60146 493774
rect 60382 493538 60466 493774
rect 60702 493538 60734 493774
rect 60114 493454 60734 493538
rect 60114 493218 60146 493454
rect 60382 493218 60466 493454
rect 60702 493218 60734 493454
rect 60114 457774 60734 493218
rect 80288 475174 80608 475206
rect 80288 474938 80330 475174
rect 80566 474938 80608 475174
rect 80288 474854 80608 474938
rect 80288 474618 80330 474854
rect 80566 474618 80608 474854
rect 80288 474586 80608 474618
rect 64928 471454 65248 471486
rect 64928 471218 64970 471454
rect 65206 471218 65248 471454
rect 64928 471134 65248 471218
rect 64928 470898 64970 471134
rect 65206 470898 65248 471134
rect 64928 470866 65248 470898
rect 95648 471454 95968 471486
rect 95648 471218 95690 471454
rect 95926 471218 95968 471454
rect 95648 471134 95968 471218
rect 95648 470898 95690 471134
rect 95926 470898 95968 471134
rect 95648 470866 95968 470898
rect 109794 471454 110414 506898
rect 109794 471218 109826 471454
rect 110062 471218 110146 471454
rect 110382 471218 110414 471454
rect 109794 471134 110414 471218
rect 109794 470898 109826 471134
rect 110062 470898 110146 471134
rect 110382 470898 110414 471134
rect 60114 457538 60146 457774
rect 60382 457538 60466 457774
rect 60702 457538 60734 457774
rect 60114 457454 60734 457538
rect 60114 457218 60146 457454
rect 60382 457218 60466 457454
rect 60702 457218 60734 457454
rect 60114 421774 60734 457218
rect 60114 421538 60146 421774
rect 60382 421538 60466 421774
rect 60702 421538 60734 421774
rect 60114 421454 60734 421538
rect 60114 421218 60146 421454
rect 60382 421218 60466 421454
rect 60702 421218 60734 421454
rect 60114 385774 60734 421218
rect 60114 385538 60146 385774
rect 60382 385538 60466 385774
rect 60702 385538 60734 385774
rect 60114 385454 60734 385538
rect 60114 385218 60146 385454
rect 60382 385218 60466 385454
rect 60702 385218 60734 385454
rect 60114 349774 60734 385218
rect 60114 349538 60146 349774
rect 60382 349538 60466 349774
rect 60702 349538 60734 349774
rect 60114 349454 60734 349538
rect 60114 349218 60146 349454
rect 60382 349218 60466 349454
rect 60702 349218 60734 349454
rect 60114 313774 60734 349218
rect 63834 425494 64454 447495
rect 63834 425258 63866 425494
rect 64102 425258 64186 425494
rect 64422 425258 64454 425494
rect 63834 425174 64454 425258
rect 63834 424938 63866 425174
rect 64102 424938 64186 425174
rect 64422 424938 64454 425174
rect 63834 389494 64454 424938
rect 63834 389258 63866 389494
rect 64102 389258 64186 389494
rect 64422 389258 64454 389494
rect 63834 389174 64454 389258
rect 63834 388938 63866 389174
rect 64102 388938 64186 389174
rect 64422 388938 64454 389174
rect 63834 353494 64454 388938
rect 63834 353258 63866 353494
rect 64102 353258 64186 353494
rect 64422 353258 64454 353494
rect 63834 353174 64454 353258
rect 63834 352938 63866 353174
rect 64102 352938 64186 353174
rect 64422 352938 64454 353174
rect 63834 320601 64454 352938
rect 73794 435454 74414 447495
rect 73794 435218 73826 435454
rect 74062 435218 74146 435454
rect 74382 435218 74414 435454
rect 73794 435134 74414 435218
rect 73794 434898 73826 435134
rect 74062 434898 74146 435134
rect 74382 434898 74414 435134
rect 73794 399454 74414 434898
rect 73794 399218 73826 399454
rect 74062 399218 74146 399454
rect 74382 399218 74414 399454
rect 73794 399134 74414 399218
rect 73794 398898 73826 399134
rect 74062 398898 74146 399134
rect 74382 398898 74414 399134
rect 73794 363454 74414 398898
rect 73794 363218 73826 363454
rect 74062 363218 74146 363454
rect 74382 363218 74414 363454
rect 73794 363134 74414 363218
rect 73794 362898 73826 363134
rect 74062 362898 74146 363134
rect 74382 362898 74414 363134
rect 73794 327454 74414 362898
rect 73794 327218 73826 327454
rect 74062 327218 74146 327454
rect 74382 327218 74414 327454
rect 73794 327134 74414 327218
rect 73794 326898 73826 327134
rect 74062 326898 74146 327134
rect 74382 326898 74414 327134
rect 73794 320601 74414 326898
rect 77514 439174 78134 447495
rect 77514 438938 77546 439174
rect 77782 438938 77866 439174
rect 78102 438938 78134 439174
rect 77514 438854 78134 438938
rect 77514 438618 77546 438854
rect 77782 438618 77866 438854
rect 78102 438618 78134 438854
rect 77514 403174 78134 438618
rect 77514 402938 77546 403174
rect 77782 402938 77866 403174
rect 78102 402938 78134 403174
rect 77514 402854 78134 402938
rect 77514 402618 77546 402854
rect 77782 402618 77866 402854
rect 78102 402618 78134 402854
rect 77514 367174 78134 402618
rect 77514 366938 77546 367174
rect 77782 366938 77866 367174
rect 78102 366938 78134 367174
rect 77514 366854 78134 366938
rect 77514 366618 77546 366854
rect 77782 366618 77866 366854
rect 78102 366618 78134 366854
rect 77514 331174 78134 366618
rect 77514 330938 77546 331174
rect 77782 330938 77866 331174
rect 78102 330938 78134 331174
rect 77514 330854 78134 330938
rect 77514 330618 77546 330854
rect 77782 330618 77866 330854
rect 78102 330618 78134 330854
rect 77514 320601 78134 330618
rect 81234 442894 81854 447495
rect 81234 442658 81266 442894
rect 81502 442658 81586 442894
rect 81822 442658 81854 442894
rect 81234 442574 81854 442658
rect 81234 442338 81266 442574
rect 81502 442338 81586 442574
rect 81822 442338 81854 442574
rect 81234 406894 81854 442338
rect 81234 406658 81266 406894
rect 81502 406658 81586 406894
rect 81822 406658 81854 406894
rect 81234 406574 81854 406658
rect 81234 406338 81266 406574
rect 81502 406338 81586 406574
rect 81822 406338 81854 406574
rect 81234 370894 81854 406338
rect 81234 370658 81266 370894
rect 81502 370658 81586 370894
rect 81822 370658 81854 370894
rect 81234 370574 81854 370658
rect 81234 370338 81266 370574
rect 81502 370338 81586 370574
rect 81822 370338 81854 370574
rect 81234 334894 81854 370338
rect 81234 334658 81266 334894
rect 81502 334658 81586 334894
rect 81822 334658 81854 334894
rect 81234 334574 81854 334658
rect 81234 334338 81266 334574
rect 81502 334338 81586 334574
rect 81822 334338 81854 334574
rect 81234 320601 81854 334338
rect 84954 446614 85574 447495
rect 84954 446378 84986 446614
rect 85222 446378 85306 446614
rect 85542 446378 85574 446614
rect 84954 446294 85574 446378
rect 84954 446058 84986 446294
rect 85222 446058 85306 446294
rect 85542 446058 85574 446294
rect 84954 410614 85574 446058
rect 84954 410378 84986 410614
rect 85222 410378 85306 410614
rect 85542 410378 85574 410614
rect 84954 410294 85574 410378
rect 84954 410058 84986 410294
rect 85222 410058 85306 410294
rect 85542 410058 85574 410294
rect 84954 374614 85574 410058
rect 84954 374378 84986 374614
rect 85222 374378 85306 374614
rect 85542 374378 85574 374614
rect 84954 374294 85574 374378
rect 84954 374058 84986 374294
rect 85222 374058 85306 374294
rect 85542 374058 85574 374294
rect 84954 338614 85574 374058
rect 84954 338378 84986 338614
rect 85222 338378 85306 338614
rect 85542 338378 85574 338614
rect 84954 338294 85574 338378
rect 84954 338058 84986 338294
rect 85222 338058 85306 338294
rect 85542 338058 85574 338294
rect 84954 320601 85574 338058
rect 88674 414334 89294 447495
rect 88674 414098 88706 414334
rect 88942 414098 89026 414334
rect 89262 414098 89294 414334
rect 88674 414014 89294 414098
rect 88674 413778 88706 414014
rect 88942 413778 89026 414014
rect 89262 413778 89294 414014
rect 88674 378334 89294 413778
rect 88674 378098 88706 378334
rect 88942 378098 89026 378334
rect 89262 378098 89294 378334
rect 88674 378014 89294 378098
rect 88674 377778 88706 378014
rect 88942 377778 89026 378014
rect 89262 377778 89294 378014
rect 88674 342334 89294 377778
rect 88674 342098 88706 342334
rect 88942 342098 89026 342334
rect 89262 342098 89294 342334
rect 88674 342014 89294 342098
rect 88674 341778 88706 342014
rect 88942 341778 89026 342014
rect 89262 341778 89294 342014
rect 88674 320601 89294 341778
rect 92394 418054 93014 447495
rect 92394 417818 92426 418054
rect 92662 417818 92746 418054
rect 92982 417818 93014 418054
rect 92394 417734 93014 417818
rect 92394 417498 92426 417734
rect 92662 417498 92746 417734
rect 92982 417498 93014 417734
rect 92394 382054 93014 417498
rect 92394 381818 92426 382054
rect 92662 381818 92746 382054
rect 92982 381818 93014 382054
rect 92394 381734 93014 381818
rect 92394 381498 92426 381734
rect 92662 381498 92746 381734
rect 92982 381498 93014 381734
rect 92394 346054 93014 381498
rect 92394 345818 92426 346054
rect 92662 345818 92746 346054
rect 92982 345818 93014 346054
rect 92394 345734 93014 345818
rect 92394 345498 92426 345734
rect 92662 345498 92746 345734
rect 92982 345498 93014 345734
rect 92394 320601 93014 345498
rect 96114 421774 96734 447495
rect 96114 421538 96146 421774
rect 96382 421538 96466 421774
rect 96702 421538 96734 421774
rect 96114 421454 96734 421538
rect 96114 421218 96146 421454
rect 96382 421218 96466 421454
rect 96702 421218 96734 421454
rect 96114 385774 96734 421218
rect 96114 385538 96146 385774
rect 96382 385538 96466 385774
rect 96702 385538 96734 385774
rect 96114 385454 96734 385538
rect 96114 385218 96146 385454
rect 96382 385218 96466 385454
rect 96702 385218 96734 385454
rect 96114 349774 96734 385218
rect 96114 349538 96146 349774
rect 96382 349538 96466 349774
rect 96702 349538 96734 349774
rect 96114 349454 96734 349538
rect 96114 349218 96146 349454
rect 96382 349218 96466 349454
rect 96702 349218 96734 349454
rect 96114 320601 96734 349218
rect 99834 425494 100454 447495
rect 99834 425258 99866 425494
rect 100102 425258 100186 425494
rect 100422 425258 100454 425494
rect 99834 425174 100454 425258
rect 99834 424938 99866 425174
rect 100102 424938 100186 425174
rect 100422 424938 100454 425174
rect 99834 389494 100454 424938
rect 99834 389258 99866 389494
rect 100102 389258 100186 389494
rect 100422 389258 100454 389494
rect 99834 389174 100454 389258
rect 99834 388938 99866 389174
rect 100102 388938 100186 389174
rect 100422 388938 100454 389174
rect 99834 353494 100454 388938
rect 99834 353258 99866 353494
rect 100102 353258 100186 353494
rect 100422 353258 100454 353494
rect 99834 353174 100454 353258
rect 99834 352938 99866 353174
rect 100102 352938 100186 353174
rect 100422 352938 100454 353174
rect 99834 320601 100454 352938
rect 109794 435454 110414 470898
rect 109794 435218 109826 435454
rect 110062 435218 110146 435454
rect 110382 435218 110414 435454
rect 109794 435134 110414 435218
rect 109794 434898 109826 435134
rect 110062 434898 110146 435134
rect 110382 434898 110414 435134
rect 109794 399454 110414 434898
rect 109794 399218 109826 399454
rect 110062 399218 110146 399454
rect 110382 399218 110414 399454
rect 109794 399134 110414 399218
rect 109794 398898 109826 399134
rect 110062 398898 110146 399134
rect 110382 398898 110414 399134
rect 109794 363454 110414 398898
rect 109794 363218 109826 363454
rect 110062 363218 110146 363454
rect 110382 363218 110414 363454
rect 109794 363134 110414 363218
rect 109794 362898 109826 363134
rect 110062 362898 110146 363134
rect 110382 362898 110414 363134
rect 109794 327454 110414 362898
rect 109794 327218 109826 327454
rect 110062 327218 110146 327454
rect 110382 327218 110414 327454
rect 109794 327134 110414 327218
rect 109794 326898 109826 327134
rect 110062 326898 110146 327134
rect 110382 326898 110414 327134
rect 60114 313538 60146 313774
rect 60382 313538 60466 313774
rect 60702 313538 60734 313774
rect 60114 313454 60734 313538
rect 60114 313218 60146 313454
rect 60382 313218 60466 313454
rect 60702 313218 60734 313454
rect 60114 277774 60734 313218
rect 80288 295174 80608 295206
rect 80288 294938 80330 295174
rect 80566 294938 80608 295174
rect 80288 294854 80608 294938
rect 80288 294618 80330 294854
rect 80566 294618 80608 294854
rect 80288 294586 80608 294618
rect 64928 291454 65248 291486
rect 64928 291218 64970 291454
rect 65206 291218 65248 291454
rect 64928 291134 65248 291218
rect 64928 290898 64970 291134
rect 65206 290898 65248 291134
rect 64928 290866 65248 290898
rect 95648 291454 95968 291486
rect 95648 291218 95690 291454
rect 95926 291218 95968 291454
rect 95648 291134 95968 291218
rect 95648 290898 95690 291134
rect 95926 290898 95968 291134
rect 95648 290866 95968 290898
rect 109794 291454 110414 326898
rect 109794 291218 109826 291454
rect 110062 291218 110146 291454
rect 110382 291218 110414 291454
rect 109794 291134 110414 291218
rect 109794 290898 109826 291134
rect 110062 290898 110146 291134
rect 110382 290898 110414 291134
rect 60114 277538 60146 277774
rect 60382 277538 60466 277774
rect 60702 277538 60734 277774
rect 60114 277454 60734 277538
rect 60114 277218 60146 277454
rect 60382 277218 60466 277454
rect 60702 277218 60734 277454
rect 60114 241774 60734 277218
rect 80288 259174 80608 259206
rect 80288 258938 80330 259174
rect 80566 258938 80608 259174
rect 80288 258854 80608 258938
rect 80288 258618 80330 258854
rect 80566 258618 80608 258854
rect 80288 258586 80608 258618
rect 64928 255454 65248 255486
rect 64928 255218 64970 255454
rect 65206 255218 65248 255454
rect 64928 255134 65248 255218
rect 64928 254898 64970 255134
rect 65206 254898 65248 255134
rect 64928 254866 65248 254898
rect 95648 255454 95968 255486
rect 95648 255218 95690 255454
rect 95926 255218 95968 255454
rect 95648 255134 95968 255218
rect 95648 254898 95690 255134
rect 95926 254898 95968 255134
rect 95648 254866 95968 254898
rect 109794 255454 110414 290898
rect 109794 255218 109826 255454
rect 110062 255218 110146 255454
rect 110382 255218 110414 255454
rect 109794 255134 110414 255218
rect 109794 254898 109826 255134
rect 110062 254898 110146 255134
rect 110382 254898 110414 255134
rect 60114 241538 60146 241774
rect 60382 241538 60466 241774
rect 60702 241538 60734 241774
rect 60114 241454 60734 241538
rect 60114 241218 60146 241454
rect 60382 241218 60466 241454
rect 60702 241218 60734 241454
rect 60114 205774 60734 241218
rect 80288 223174 80608 223206
rect 80288 222938 80330 223174
rect 80566 222938 80608 223174
rect 80288 222854 80608 222938
rect 80288 222618 80330 222854
rect 80566 222618 80608 222854
rect 80288 222586 80608 222618
rect 64928 219454 65248 219486
rect 64928 219218 64970 219454
rect 65206 219218 65248 219454
rect 64928 219134 65248 219218
rect 64928 218898 64970 219134
rect 65206 218898 65248 219134
rect 64928 218866 65248 218898
rect 95648 219454 95968 219486
rect 95648 219218 95690 219454
rect 95926 219218 95968 219454
rect 95648 219134 95968 219218
rect 95648 218898 95690 219134
rect 95926 218898 95968 219134
rect 95648 218866 95968 218898
rect 109794 219454 110414 254898
rect 109794 219218 109826 219454
rect 110062 219218 110146 219454
rect 110382 219218 110414 219454
rect 109794 219134 110414 219218
rect 109794 218898 109826 219134
rect 110062 218898 110146 219134
rect 110382 218898 110414 219134
rect 60114 205538 60146 205774
rect 60382 205538 60466 205774
rect 60702 205538 60734 205774
rect 60114 205454 60734 205538
rect 60114 205218 60146 205454
rect 60382 205218 60466 205454
rect 60702 205218 60734 205454
rect 60114 169774 60734 205218
rect 80288 187174 80608 187206
rect 80288 186938 80330 187174
rect 80566 186938 80608 187174
rect 80288 186854 80608 186938
rect 80288 186618 80330 186854
rect 80566 186618 80608 186854
rect 80288 186586 80608 186618
rect 64928 183454 65248 183486
rect 64928 183218 64970 183454
rect 65206 183218 65248 183454
rect 64928 183134 65248 183218
rect 64928 182898 64970 183134
rect 65206 182898 65248 183134
rect 64928 182866 65248 182898
rect 95648 183454 95968 183486
rect 95648 183218 95690 183454
rect 95926 183218 95968 183454
rect 95648 183134 95968 183218
rect 95648 182898 95690 183134
rect 95926 182898 95968 183134
rect 95648 182866 95968 182898
rect 109794 183454 110414 218898
rect 109794 183218 109826 183454
rect 110062 183218 110146 183454
rect 110382 183218 110414 183454
rect 109794 183134 110414 183218
rect 109794 182898 109826 183134
rect 110062 182898 110146 183134
rect 110382 182898 110414 183134
rect 60114 169538 60146 169774
rect 60382 169538 60466 169774
rect 60702 169538 60734 169774
rect 60114 169454 60734 169538
rect 60114 169218 60146 169454
rect 60382 169218 60466 169454
rect 60702 169218 60734 169454
rect 60114 133774 60734 169218
rect 60114 133538 60146 133774
rect 60382 133538 60466 133774
rect 60702 133538 60734 133774
rect 60114 133454 60734 133538
rect 60114 133218 60146 133454
rect 60382 133218 60466 133454
rect 60702 133218 60734 133454
rect 60114 133057 60734 133218
rect 88674 162334 89294 167495
rect 88674 162098 88706 162334
rect 88942 162098 89026 162334
rect 89262 162098 89294 162334
rect 88674 162014 89294 162098
rect 88674 161778 88706 162014
rect 88942 161778 89026 162014
rect 89262 161778 89294 162014
rect 88674 133057 89294 161778
rect 92394 166054 93014 167495
rect 92394 165818 92426 166054
rect 92662 165818 92746 166054
rect 92982 165818 93014 166054
rect 92394 165734 93014 165818
rect 92394 165498 92426 165734
rect 92662 165498 92746 165734
rect 92982 165498 93014 165734
rect 92394 133057 93014 165498
rect 96114 133774 96734 167495
rect 96114 133538 96146 133774
rect 96382 133538 96466 133774
rect 96702 133538 96734 133774
rect 96114 133454 96734 133538
rect 96114 133218 96146 133454
rect 96382 133218 96466 133454
rect 96702 133218 96734 133454
rect 96114 133057 96734 133218
rect 109794 147454 110414 182898
rect 109794 147218 109826 147454
rect 110062 147218 110146 147454
rect 110382 147218 110414 147454
rect 109794 147134 110414 147218
rect 109794 146898 109826 147134
rect 110062 146898 110146 147134
rect 110382 146898 110414 147134
rect 109794 133057 110414 146898
rect 113514 705798 114134 711590
rect 113514 705562 113546 705798
rect 113782 705562 113866 705798
rect 114102 705562 114134 705798
rect 113514 705478 114134 705562
rect 113514 705242 113546 705478
rect 113782 705242 113866 705478
rect 114102 705242 114134 705478
rect 113514 691174 114134 705242
rect 113514 690938 113546 691174
rect 113782 690938 113866 691174
rect 114102 690938 114134 691174
rect 113514 690854 114134 690938
rect 113514 690618 113546 690854
rect 113782 690618 113866 690854
rect 114102 690618 114134 690854
rect 113514 655174 114134 690618
rect 113514 654938 113546 655174
rect 113782 654938 113866 655174
rect 114102 654938 114134 655174
rect 113514 654854 114134 654938
rect 113514 654618 113546 654854
rect 113782 654618 113866 654854
rect 114102 654618 114134 654854
rect 113514 619174 114134 654618
rect 113514 618938 113546 619174
rect 113782 618938 113866 619174
rect 114102 618938 114134 619174
rect 113514 618854 114134 618938
rect 113514 618618 113546 618854
rect 113782 618618 113866 618854
rect 114102 618618 114134 618854
rect 113514 583174 114134 618618
rect 113514 582938 113546 583174
rect 113782 582938 113866 583174
rect 114102 582938 114134 583174
rect 113514 582854 114134 582938
rect 113514 582618 113546 582854
rect 113782 582618 113866 582854
rect 114102 582618 114134 582854
rect 113514 547174 114134 582618
rect 113514 546938 113546 547174
rect 113782 546938 113866 547174
rect 114102 546938 114134 547174
rect 113514 546854 114134 546938
rect 113514 546618 113546 546854
rect 113782 546618 113866 546854
rect 114102 546618 114134 546854
rect 113514 511174 114134 546618
rect 113514 510938 113546 511174
rect 113782 510938 113866 511174
rect 114102 510938 114134 511174
rect 113514 510854 114134 510938
rect 113514 510618 113546 510854
rect 113782 510618 113866 510854
rect 114102 510618 114134 510854
rect 113514 475174 114134 510618
rect 113514 474938 113546 475174
rect 113782 474938 113866 475174
rect 114102 474938 114134 475174
rect 113514 474854 114134 474938
rect 113514 474618 113546 474854
rect 113782 474618 113866 474854
rect 114102 474618 114134 474854
rect 113514 439174 114134 474618
rect 113514 438938 113546 439174
rect 113782 438938 113866 439174
rect 114102 438938 114134 439174
rect 113514 438854 114134 438938
rect 113514 438618 113546 438854
rect 113782 438618 113866 438854
rect 114102 438618 114134 438854
rect 113514 403174 114134 438618
rect 113514 402938 113546 403174
rect 113782 402938 113866 403174
rect 114102 402938 114134 403174
rect 113514 402854 114134 402938
rect 113514 402618 113546 402854
rect 113782 402618 113866 402854
rect 114102 402618 114134 402854
rect 113514 367174 114134 402618
rect 113514 366938 113546 367174
rect 113782 366938 113866 367174
rect 114102 366938 114134 367174
rect 113514 366854 114134 366938
rect 113514 366618 113546 366854
rect 113782 366618 113866 366854
rect 114102 366618 114134 366854
rect 113514 331174 114134 366618
rect 113514 330938 113546 331174
rect 113782 330938 113866 331174
rect 114102 330938 114134 331174
rect 113514 330854 114134 330938
rect 113514 330618 113546 330854
rect 113782 330618 113866 330854
rect 114102 330618 114134 330854
rect 113514 295174 114134 330618
rect 113514 294938 113546 295174
rect 113782 294938 113866 295174
rect 114102 294938 114134 295174
rect 113514 294854 114134 294938
rect 113514 294618 113546 294854
rect 113782 294618 113866 294854
rect 114102 294618 114134 294854
rect 113514 259174 114134 294618
rect 113514 258938 113546 259174
rect 113782 258938 113866 259174
rect 114102 258938 114134 259174
rect 113514 258854 114134 258938
rect 113514 258618 113546 258854
rect 113782 258618 113866 258854
rect 114102 258618 114134 258854
rect 113514 223174 114134 258618
rect 113514 222938 113546 223174
rect 113782 222938 113866 223174
rect 114102 222938 114134 223174
rect 113514 222854 114134 222938
rect 113514 222618 113546 222854
rect 113782 222618 113866 222854
rect 114102 222618 114134 222854
rect 113514 187174 114134 222618
rect 113514 186938 113546 187174
rect 113782 186938 113866 187174
rect 114102 186938 114134 187174
rect 113514 186854 114134 186938
rect 113514 186618 113546 186854
rect 113782 186618 113866 186854
rect 114102 186618 114134 186854
rect 113514 151174 114134 186618
rect 113514 150938 113546 151174
rect 113782 150938 113866 151174
rect 114102 150938 114134 151174
rect 113514 150854 114134 150938
rect 113514 150618 113546 150854
rect 113782 150618 113866 150854
rect 114102 150618 114134 150854
rect 113514 133057 114134 150618
rect 117234 706758 117854 711590
rect 117234 706522 117266 706758
rect 117502 706522 117586 706758
rect 117822 706522 117854 706758
rect 117234 706438 117854 706522
rect 117234 706202 117266 706438
rect 117502 706202 117586 706438
rect 117822 706202 117854 706438
rect 117234 694894 117854 706202
rect 117234 694658 117266 694894
rect 117502 694658 117586 694894
rect 117822 694658 117854 694894
rect 117234 694574 117854 694658
rect 117234 694338 117266 694574
rect 117502 694338 117586 694574
rect 117822 694338 117854 694574
rect 117234 658894 117854 694338
rect 117234 658658 117266 658894
rect 117502 658658 117586 658894
rect 117822 658658 117854 658894
rect 117234 658574 117854 658658
rect 117234 658338 117266 658574
rect 117502 658338 117586 658574
rect 117822 658338 117854 658574
rect 117234 622894 117854 658338
rect 117234 622658 117266 622894
rect 117502 622658 117586 622894
rect 117822 622658 117854 622894
rect 117234 622574 117854 622658
rect 117234 622338 117266 622574
rect 117502 622338 117586 622574
rect 117822 622338 117854 622574
rect 117234 586894 117854 622338
rect 117234 586658 117266 586894
rect 117502 586658 117586 586894
rect 117822 586658 117854 586894
rect 117234 586574 117854 586658
rect 117234 586338 117266 586574
rect 117502 586338 117586 586574
rect 117822 586338 117854 586574
rect 117234 550894 117854 586338
rect 117234 550658 117266 550894
rect 117502 550658 117586 550894
rect 117822 550658 117854 550894
rect 117234 550574 117854 550658
rect 117234 550338 117266 550574
rect 117502 550338 117586 550574
rect 117822 550338 117854 550574
rect 117234 514894 117854 550338
rect 117234 514658 117266 514894
rect 117502 514658 117586 514894
rect 117822 514658 117854 514894
rect 117234 514574 117854 514658
rect 117234 514338 117266 514574
rect 117502 514338 117586 514574
rect 117822 514338 117854 514574
rect 117234 478894 117854 514338
rect 117234 478658 117266 478894
rect 117502 478658 117586 478894
rect 117822 478658 117854 478894
rect 117234 478574 117854 478658
rect 117234 478338 117266 478574
rect 117502 478338 117586 478574
rect 117822 478338 117854 478574
rect 117234 442894 117854 478338
rect 117234 442658 117266 442894
rect 117502 442658 117586 442894
rect 117822 442658 117854 442894
rect 117234 442574 117854 442658
rect 117234 442338 117266 442574
rect 117502 442338 117586 442574
rect 117822 442338 117854 442574
rect 117234 406894 117854 442338
rect 117234 406658 117266 406894
rect 117502 406658 117586 406894
rect 117822 406658 117854 406894
rect 117234 406574 117854 406658
rect 117234 406338 117266 406574
rect 117502 406338 117586 406574
rect 117822 406338 117854 406574
rect 117234 370894 117854 406338
rect 117234 370658 117266 370894
rect 117502 370658 117586 370894
rect 117822 370658 117854 370894
rect 117234 370574 117854 370658
rect 117234 370338 117266 370574
rect 117502 370338 117586 370574
rect 117822 370338 117854 370574
rect 117234 334894 117854 370338
rect 117234 334658 117266 334894
rect 117502 334658 117586 334894
rect 117822 334658 117854 334894
rect 117234 334574 117854 334658
rect 117234 334338 117266 334574
rect 117502 334338 117586 334574
rect 117822 334338 117854 334574
rect 117234 298894 117854 334338
rect 117234 298658 117266 298894
rect 117502 298658 117586 298894
rect 117822 298658 117854 298894
rect 117234 298574 117854 298658
rect 117234 298338 117266 298574
rect 117502 298338 117586 298574
rect 117822 298338 117854 298574
rect 117234 262894 117854 298338
rect 117234 262658 117266 262894
rect 117502 262658 117586 262894
rect 117822 262658 117854 262894
rect 117234 262574 117854 262658
rect 117234 262338 117266 262574
rect 117502 262338 117586 262574
rect 117822 262338 117854 262574
rect 117234 226894 117854 262338
rect 117234 226658 117266 226894
rect 117502 226658 117586 226894
rect 117822 226658 117854 226894
rect 117234 226574 117854 226658
rect 117234 226338 117266 226574
rect 117502 226338 117586 226574
rect 117822 226338 117854 226574
rect 117234 190894 117854 226338
rect 117234 190658 117266 190894
rect 117502 190658 117586 190894
rect 117822 190658 117854 190894
rect 117234 190574 117854 190658
rect 117234 190338 117266 190574
rect 117502 190338 117586 190574
rect 117822 190338 117854 190574
rect 117234 154894 117854 190338
rect 117234 154658 117266 154894
rect 117502 154658 117586 154894
rect 117822 154658 117854 154894
rect 117234 154574 117854 154658
rect 117234 154338 117266 154574
rect 117502 154338 117586 154574
rect 117822 154338 117854 154574
rect 117234 133057 117854 154338
rect 120954 707718 121574 711590
rect 120954 707482 120986 707718
rect 121222 707482 121306 707718
rect 121542 707482 121574 707718
rect 120954 707398 121574 707482
rect 120954 707162 120986 707398
rect 121222 707162 121306 707398
rect 121542 707162 121574 707398
rect 120954 698614 121574 707162
rect 120954 698378 120986 698614
rect 121222 698378 121306 698614
rect 121542 698378 121574 698614
rect 120954 698294 121574 698378
rect 120954 698058 120986 698294
rect 121222 698058 121306 698294
rect 121542 698058 121574 698294
rect 120954 662614 121574 698058
rect 120954 662378 120986 662614
rect 121222 662378 121306 662614
rect 121542 662378 121574 662614
rect 120954 662294 121574 662378
rect 120954 662058 120986 662294
rect 121222 662058 121306 662294
rect 121542 662058 121574 662294
rect 120954 626614 121574 662058
rect 120954 626378 120986 626614
rect 121222 626378 121306 626614
rect 121542 626378 121574 626614
rect 120954 626294 121574 626378
rect 120954 626058 120986 626294
rect 121222 626058 121306 626294
rect 121542 626058 121574 626294
rect 120954 590614 121574 626058
rect 120954 590378 120986 590614
rect 121222 590378 121306 590614
rect 121542 590378 121574 590614
rect 120954 590294 121574 590378
rect 120954 590058 120986 590294
rect 121222 590058 121306 590294
rect 121542 590058 121574 590294
rect 120954 554614 121574 590058
rect 120954 554378 120986 554614
rect 121222 554378 121306 554614
rect 121542 554378 121574 554614
rect 120954 554294 121574 554378
rect 120954 554058 120986 554294
rect 121222 554058 121306 554294
rect 121542 554058 121574 554294
rect 120954 518614 121574 554058
rect 120954 518378 120986 518614
rect 121222 518378 121306 518614
rect 121542 518378 121574 518614
rect 120954 518294 121574 518378
rect 120954 518058 120986 518294
rect 121222 518058 121306 518294
rect 121542 518058 121574 518294
rect 120954 482614 121574 518058
rect 120954 482378 120986 482614
rect 121222 482378 121306 482614
rect 121542 482378 121574 482614
rect 120954 482294 121574 482378
rect 120954 482058 120986 482294
rect 121222 482058 121306 482294
rect 121542 482058 121574 482294
rect 120954 446614 121574 482058
rect 120954 446378 120986 446614
rect 121222 446378 121306 446614
rect 121542 446378 121574 446614
rect 120954 446294 121574 446378
rect 120954 446058 120986 446294
rect 121222 446058 121306 446294
rect 121542 446058 121574 446294
rect 120954 410614 121574 446058
rect 120954 410378 120986 410614
rect 121222 410378 121306 410614
rect 121542 410378 121574 410614
rect 120954 410294 121574 410378
rect 120954 410058 120986 410294
rect 121222 410058 121306 410294
rect 121542 410058 121574 410294
rect 120954 374614 121574 410058
rect 120954 374378 120986 374614
rect 121222 374378 121306 374614
rect 121542 374378 121574 374614
rect 120954 374294 121574 374378
rect 120954 374058 120986 374294
rect 121222 374058 121306 374294
rect 121542 374058 121574 374294
rect 120954 338614 121574 374058
rect 120954 338378 120986 338614
rect 121222 338378 121306 338614
rect 121542 338378 121574 338614
rect 120954 338294 121574 338378
rect 120954 338058 120986 338294
rect 121222 338058 121306 338294
rect 121542 338058 121574 338294
rect 120954 302614 121574 338058
rect 120954 302378 120986 302614
rect 121222 302378 121306 302614
rect 121542 302378 121574 302614
rect 120954 302294 121574 302378
rect 120954 302058 120986 302294
rect 121222 302058 121306 302294
rect 121542 302058 121574 302294
rect 120954 266614 121574 302058
rect 120954 266378 120986 266614
rect 121222 266378 121306 266614
rect 121542 266378 121574 266614
rect 120954 266294 121574 266378
rect 120954 266058 120986 266294
rect 121222 266058 121306 266294
rect 121542 266058 121574 266294
rect 120954 230614 121574 266058
rect 120954 230378 120986 230614
rect 121222 230378 121306 230614
rect 121542 230378 121574 230614
rect 120954 230294 121574 230378
rect 120954 230058 120986 230294
rect 121222 230058 121306 230294
rect 121542 230058 121574 230294
rect 120954 194614 121574 230058
rect 120954 194378 120986 194614
rect 121222 194378 121306 194614
rect 121542 194378 121574 194614
rect 120954 194294 121574 194378
rect 120954 194058 120986 194294
rect 121222 194058 121306 194294
rect 121542 194058 121574 194294
rect 120954 158614 121574 194058
rect 120954 158378 120986 158614
rect 121222 158378 121306 158614
rect 121542 158378 121574 158614
rect 120954 158294 121574 158378
rect 120954 158058 120986 158294
rect 121222 158058 121306 158294
rect 121542 158058 121574 158294
rect 120954 133057 121574 158058
rect 124674 708678 125294 711590
rect 124674 708442 124706 708678
rect 124942 708442 125026 708678
rect 125262 708442 125294 708678
rect 124674 708358 125294 708442
rect 124674 708122 124706 708358
rect 124942 708122 125026 708358
rect 125262 708122 125294 708358
rect 124674 666334 125294 708122
rect 124674 666098 124706 666334
rect 124942 666098 125026 666334
rect 125262 666098 125294 666334
rect 124674 666014 125294 666098
rect 124674 665778 124706 666014
rect 124942 665778 125026 666014
rect 125262 665778 125294 666014
rect 124674 630334 125294 665778
rect 124674 630098 124706 630334
rect 124942 630098 125026 630334
rect 125262 630098 125294 630334
rect 124674 630014 125294 630098
rect 124674 629778 124706 630014
rect 124942 629778 125026 630014
rect 125262 629778 125294 630014
rect 124674 594334 125294 629778
rect 124674 594098 124706 594334
rect 124942 594098 125026 594334
rect 125262 594098 125294 594334
rect 124674 594014 125294 594098
rect 124674 593778 124706 594014
rect 124942 593778 125026 594014
rect 125262 593778 125294 594014
rect 124674 558334 125294 593778
rect 124674 558098 124706 558334
rect 124942 558098 125026 558334
rect 125262 558098 125294 558334
rect 124674 558014 125294 558098
rect 124674 557778 124706 558014
rect 124942 557778 125026 558014
rect 125262 557778 125294 558014
rect 124674 522334 125294 557778
rect 124674 522098 124706 522334
rect 124942 522098 125026 522334
rect 125262 522098 125294 522334
rect 124674 522014 125294 522098
rect 124674 521778 124706 522014
rect 124942 521778 125026 522014
rect 125262 521778 125294 522014
rect 124674 486334 125294 521778
rect 124674 486098 124706 486334
rect 124942 486098 125026 486334
rect 125262 486098 125294 486334
rect 124674 486014 125294 486098
rect 124674 485778 124706 486014
rect 124942 485778 125026 486014
rect 125262 485778 125294 486014
rect 124674 450334 125294 485778
rect 124674 450098 124706 450334
rect 124942 450098 125026 450334
rect 125262 450098 125294 450334
rect 124674 450014 125294 450098
rect 124674 449778 124706 450014
rect 124942 449778 125026 450014
rect 125262 449778 125294 450014
rect 124674 414334 125294 449778
rect 124674 414098 124706 414334
rect 124942 414098 125026 414334
rect 125262 414098 125294 414334
rect 124674 414014 125294 414098
rect 124674 413778 124706 414014
rect 124942 413778 125026 414014
rect 125262 413778 125294 414014
rect 124674 378334 125294 413778
rect 124674 378098 124706 378334
rect 124942 378098 125026 378334
rect 125262 378098 125294 378334
rect 124674 378014 125294 378098
rect 124674 377778 124706 378014
rect 124942 377778 125026 378014
rect 125262 377778 125294 378014
rect 124674 342334 125294 377778
rect 124674 342098 124706 342334
rect 124942 342098 125026 342334
rect 125262 342098 125294 342334
rect 124674 342014 125294 342098
rect 124674 341778 124706 342014
rect 124942 341778 125026 342014
rect 125262 341778 125294 342014
rect 124674 306334 125294 341778
rect 124674 306098 124706 306334
rect 124942 306098 125026 306334
rect 125262 306098 125294 306334
rect 124674 306014 125294 306098
rect 124674 305778 124706 306014
rect 124942 305778 125026 306014
rect 125262 305778 125294 306014
rect 124674 270334 125294 305778
rect 124674 270098 124706 270334
rect 124942 270098 125026 270334
rect 125262 270098 125294 270334
rect 124674 270014 125294 270098
rect 124674 269778 124706 270014
rect 124942 269778 125026 270014
rect 125262 269778 125294 270014
rect 124674 234334 125294 269778
rect 124674 234098 124706 234334
rect 124942 234098 125026 234334
rect 125262 234098 125294 234334
rect 124674 234014 125294 234098
rect 124674 233778 124706 234014
rect 124942 233778 125026 234014
rect 125262 233778 125294 234014
rect 124674 198334 125294 233778
rect 124674 198098 124706 198334
rect 124942 198098 125026 198334
rect 125262 198098 125294 198334
rect 124674 198014 125294 198098
rect 124674 197778 124706 198014
rect 124942 197778 125026 198014
rect 125262 197778 125294 198014
rect 124674 162334 125294 197778
rect 124674 162098 124706 162334
rect 124942 162098 125026 162334
rect 125262 162098 125294 162334
rect 124674 162014 125294 162098
rect 124674 161778 124706 162014
rect 124942 161778 125026 162014
rect 125262 161778 125294 162014
rect 124674 133057 125294 161778
rect 128394 709638 129014 711590
rect 128394 709402 128426 709638
rect 128662 709402 128746 709638
rect 128982 709402 129014 709638
rect 128394 709318 129014 709402
rect 128394 709082 128426 709318
rect 128662 709082 128746 709318
rect 128982 709082 129014 709318
rect 128394 670054 129014 709082
rect 128394 669818 128426 670054
rect 128662 669818 128746 670054
rect 128982 669818 129014 670054
rect 128394 669734 129014 669818
rect 128394 669498 128426 669734
rect 128662 669498 128746 669734
rect 128982 669498 129014 669734
rect 128394 634054 129014 669498
rect 128394 633818 128426 634054
rect 128662 633818 128746 634054
rect 128982 633818 129014 634054
rect 128394 633734 129014 633818
rect 128394 633498 128426 633734
rect 128662 633498 128746 633734
rect 128982 633498 129014 633734
rect 128394 598054 129014 633498
rect 128394 597818 128426 598054
rect 128662 597818 128746 598054
rect 128982 597818 129014 598054
rect 128394 597734 129014 597818
rect 128394 597498 128426 597734
rect 128662 597498 128746 597734
rect 128982 597498 129014 597734
rect 128394 562054 129014 597498
rect 128394 561818 128426 562054
rect 128662 561818 128746 562054
rect 128982 561818 129014 562054
rect 128394 561734 129014 561818
rect 128394 561498 128426 561734
rect 128662 561498 128746 561734
rect 128982 561498 129014 561734
rect 128394 526054 129014 561498
rect 128394 525818 128426 526054
rect 128662 525818 128746 526054
rect 128982 525818 129014 526054
rect 128394 525734 129014 525818
rect 128394 525498 128426 525734
rect 128662 525498 128746 525734
rect 128982 525498 129014 525734
rect 128394 490054 129014 525498
rect 128394 489818 128426 490054
rect 128662 489818 128746 490054
rect 128982 489818 129014 490054
rect 128394 489734 129014 489818
rect 128394 489498 128426 489734
rect 128662 489498 128746 489734
rect 128982 489498 129014 489734
rect 128394 454054 129014 489498
rect 128394 453818 128426 454054
rect 128662 453818 128746 454054
rect 128982 453818 129014 454054
rect 128394 453734 129014 453818
rect 128394 453498 128426 453734
rect 128662 453498 128746 453734
rect 128982 453498 129014 453734
rect 128394 418054 129014 453498
rect 128394 417818 128426 418054
rect 128662 417818 128746 418054
rect 128982 417818 129014 418054
rect 128394 417734 129014 417818
rect 128394 417498 128426 417734
rect 128662 417498 128746 417734
rect 128982 417498 129014 417734
rect 128394 382054 129014 417498
rect 128394 381818 128426 382054
rect 128662 381818 128746 382054
rect 128982 381818 129014 382054
rect 128394 381734 129014 381818
rect 128394 381498 128426 381734
rect 128662 381498 128746 381734
rect 128982 381498 129014 381734
rect 128394 346054 129014 381498
rect 128394 345818 128426 346054
rect 128662 345818 128746 346054
rect 128982 345818 129014 346054
rect 128394 345734 129014 345818
rect 128394 345498 128426 345734
rect 128662 345498 128746 345734
rect 128982 345498 129014 345734
rect 128394 310054 129014 345498
rect 128394 309818 128426 310054
rect 128662 309818 128746 310054
rect 128982 309818 129014 310054
rect 128394 309734 129014 309818
rect 128394 309498 128426 309734
rect 128662 309498 128746 309734
rect 128982 309498 129014 309734
rect 128394 274054 129014 309498
rect 128394 273818 128426 274054
rect 128662 273818 128746 274054
rect 128982 273818 129014 274054
rect 128394 273734 129014 273818
rect 128394 273498 128426 273734
rect 128662 273498 128746 273734
rect 128982 273498 129014 273734
rect 128394 238054 129014 273498
rect 128394 237818 128426 238054
rect 128662 237818 128746 238054
rect 128982 237818 129014 238054
rect 128394 237734 129014 237818
rect 128394 237498 128426 237734
rect 128662 237498 128746 237734
rect 128982 237498 129014 237734
rect 128394 202054 129014 237498
rect 128394 201818 128426 202054
rect 128662 201818 128746 202054
rect 128982 201818 129014 202054
rect 128394 201734 129014 201818
rect 128394 201498 128426 201734
rect 128662 201498 128746 201734
rect 128982 201498 129014 201734
rect 128394 166054 129014 201498
rect 128394 165818 128426 166054
rect 128662 165818 128746 166054
rect 128982 165818 129014 166054
rect 128394 165734 129014 165818
rect 128394 165498 128426 165734
rect 128662 165498 128746 165734
rect 128982 165498 129014 165734
rect 128394 133057 129014 165498
rect 132114 710598 132734 711590
rect 132114 710362 132146 710598
rect 132382 710362 132466 710598
rect 132702 710362 132734 710598
rect 132114 710278 132734 710362
rect 132114 710042 132146 710278
rect 132382 710042 132466 710278
rect 132702 710042 132734 710278
rect 132114 673774 132734 710042
rect 132114 673538 132146 673774
rect 132382 673538 132466 673774
rect 132702 673538 132734 673774
rect 132114 673454 132734 673538
rect 132114 673218 132146 673454
rect 132382 673218 132466 673454
rect 132702 673218 132734 673454
rect 132114 637774 132734 673218
rect 132114 637538 132146 637774
rect 132382 637538 132466 637774
rect 132702 637538 132734 637774
rect 132114 637454 132734 637538
rect 132114 637218 132146 637454
rect 132382 637218 132466 637454
rect 132702 637218 132734 637454
rect 132114 601774 132734 637218
rect 132114 601538 132146 601774
rect 132382 601538 132466 601774
rect 132702 601538 132734 601774
rect 132114 601454 132734 601538
rect 132114 601218 132146 601454
rect 132382 601218 132466 601454
rect 132702 601218 132734 601454
rect 132114 565774 132734 601218
rect 132114 565538 132146 565774
rect 132382 565538 132466 565774
rect 132702 565538 132734 565774
rect 132114 565454 132734 565538
rect 132114 565218 132146 565454
rect 132382 565218 132466 565454
rect 132702 565218 132734 565454
rect 132114 529774 132734 565218
rect 132114 529538 132146 529774
rect 132382 529538 132466 529774
rect 132702 529538 132734 529774
rect 132114 529454 132734 529538
rect 132114 529218 132146 529454
rect 132382 529218 132466 529454
rect 132702 529218 132734 529454
rect 132114 493774 132734 529218
rect 132114 493538 132146 493774
rect 132382 493538 132466 493774
rect 132702 493538 132734 493774
rect 132114 493454 132734 493538
rect 132114 493218 132146 493454
rect 132382 493218 132466 493454
rect 132702 493218 132734 493454
rect 132114 457774 132734 493218
rect 132114 457538 132146 457774
rect 132382 457538 132466 457774
rect 132702 457538 132734 457774
rect 132114 457454 132734 457538
rect 132114 457218 132146 457454
rect 132382 457218 132466 457454
rect 132702 457218 132734 457454
rect 132114 421774 132734 457218
rect 132114 421538 132146 421774
rect 132382 421538 132466 421774
rect 132702 421538 132734 421774
rect 132114 421454 132734 421538
rect 132114 421218 132146 421454
rect 132382 421218 132466 421454
rect 132702 421218 132734 421454
rect 132114 385774 132734 421218
rect 132114 385538 132146 385774
rect 132382 385538 132466 385774
rect 132702 385538 132734 385774
rect 132114 385454 132734 385538
rect 132114 385218 132146 385454
rect 132382 385218 132466 385454
rect 132702 385218 132734 385454
rect 132114 349774 132734 385218
rect 132114 349538 132146 349774
rect 132382 349538 132466 349774
rect 132702 349538 132734 349774
rect 132114 349454 132734 349538
rect 132114 349218 132146 349454
rect 132382 349218 132466 349454
rect 132702 349218 132734 349454
rect 132114 313774 132734 349218
rect 132114 313538 132146 313774
rect 132382 313538 132466 313774
rect 132702 313538 132734 313774
rect 132114 313454 132734 313538
rect 132114 313218 132146 313454
rect 132382 313218 132466 313454
rect 132702 313218 132734 313454
rect 132114 277774 132734 313218
rect 132114 277538 132146 277774
rect 132382 277538 132466 277774
rect 132702 277538 132734 277774
rect 132114 277454 132734 277538
rect 132114 277218 132146 277454
rect 132382 277218 132466 277454
rect 132702 277218 132734 277454
rect 132114 241774 132734 277218
rect 132114 241538 132146 241774
rect 132382 241538 132466 241774
rect 132702 241538 132734 241774
rect 132114 241454 132734 241538
rect 132114 241218 132146 241454
rect 132382 241218 132466 241454
rect 132702 241218 132734 241454
rect 132114 205774 132734 241218
rect 132114 205538 132146 205774
rect 132382 205538 132466 205774
rect 132702 205538 132734 205774
rect 132114 205454 132734 205538
rect 132114 205218 132146 205454
rect 132382 205218 132466 205454
rect 132702 205218 132734 205454
rect 132114 169774 132734 205218
rect 132114 169538 132146 169774
rect 132382 169538 132466 169774
rect 132702 169538 132734 169774
rect 132114 169454 132734 169538
rect 132114 169218 132146 169454
rect 132382 169218 132466 169454
rect 132702 169218 132734 169454
rect 132114 133774 132734 169218
rect 132114 133538 132146 133774
rect 132382 133538 132466 133774
rect 132702 133538 132734 133774
rect 132114 133454 132734 133538
rect 132114 133218 132146 133454
rect 132382 133218 132466 133454
rect 132702 133218 132734 133454
rect 132114 133057 132734 133218
rect 135834 711558 136454 711590
rect 135834 711322 135866 711558
rect 136102 711322 136186 711558
rect 136422 711322 136454 711558
rect 135834 711238 136454 711322
rect 135834 711002 135866 711238
rect 136102 711002 136186 711238
rect 136422 711002 136454 711238
rect 135834 677494 136454 711002
rect 135834 677258 135866 677494
rect 136102 677258 136186 677494
rect 136422 677258 136454 677494
rect 135834 677174 136454 677258
rect 135834 676938 135866 677174
rect 136102 676938 136186 677174
rect 136422 676938 136454 677174
rect 135834 641494 136454 676938
rect 135834 641258 135866 641494
rect 136102 641258 136186 641494
rect 136422 641258 136454 641494
rect 135834 641174 136454 641258
rect 135834 640938 135866 641174
rect 136102 640938 136186 641174
rect 136422 640938 136454 641174
rect 135834 605494 136454 640938
rect 135834 605258 135866 605494
rect 136102 605258 136186 605494
rect 136422 605258 136454 605494
rect 135834 605174 136454 605258
rect 135834 604938 135866 605174
rect 136102 604938 136186 605174
rect 136422 604938 136454 605174
rect 135834 569494 136454 604938
rect 135834 569258 135866 569494
rect 136102 569258 136186 569494
rect 136422 569258 136454 569494
rect 135834 569174 136454 569258
rect 135834 568938 135866 569174
rect 136102 568938 136186 569174
rect 136422 568938 136454 569174
rect 135834 533494 136454 568938
rect 135834 533258 135866 533494
rect 136102 533258 136186 533494
rect 136422 533258 136454 533494
rect 135834 533174 136454 533258
rect 135834 532938 135866 533174
rect 136102 532938 136186 533174
rect 136422 532938 136454 533174
rect 135834 497494 136454 532938
rect 135834 497258 135866 497494
rect 136102 497258 136186 497494
rect 136422 497258 136454 497494
rect 135834 497174 136454 497258
rect 135834 496938 135866 497174
rect 136102 496938 136186 497174
rect 136422 496938 136454 497174
rect 135834 461494 136454 496938
rect 135834 461258 135866 461494
rect 136102 461258 136186 461494
rect 136422 461258 136454 461494
rect 135834 461174 136454 461258
rect 135834 460938 135866 461174
rect 136102 460938 136186 461174
rect 136422 460938 136454 461174
rect 135834 425494 136454 460938
rect 135834 425258 135866 425494
rect 136102 425258 136186 425494
rect 136422 425258 136454 425494
rect 135834 425174 136454 425258
rect 135834 424938 135866 425174
rect 136102 424938 136186 425174
rect 136422 424938 136454 425174
rect 135834 389494 136454 424938
rect 135834 389258 135866 389494
rect 136102 389258 136186 389494
rect 136422 389258 136454 389494
rect 135834 389174 136454 389258
rect 135834 388938 135866 389174
rect 136102 388938 136186 389174
rect 136422 388938 136454 389174
rect 135834 353494 136454 388938
rect 135834 353258 135866 353494
rect 136102 353258 136186 353494
rect 136422 353258 136454 353494
rect 135834 353174 136454 353258
rect 135834 352938 135866 353174
rect 136102 352938 136186 353174
rect 136422 352938 136454 353174
rect 135834 317494 136454 352938
rect 135834 317258 135866 317494
rect 136102 317258 136186 317494
rect 136422 317258 136454 317494
rect 135834 317174 136454 317258
rect 135834 316938 135866 317174
rect 136102 316938 136186 317174
rect 136422 316938 136454 317174
rect 135834 281494 136454 316938
rect 135834 281258 135866 281494
rect 136102 281258 136186 281494
rect 136422 281258 136454 281494
rect 135834 281174 136454 281258
rect 135834 280938 135866 281174
rect 136102 280938 136186 281174
rect 136422 280938 136454 281174
rect 135834 245494 136454 280938
rect 135834 245258 135866 245494
rect 136102 245258 136186 245494
rect 136422 245258 136454 245494
rect 135834 245174 136454 245258
rect 135834 244938 135866 245174
rect 136102 244938 136186 245174
rect 136422 244938 136454 245174
rect 135834 209494 136454 244938
rect 135834 209258 135866 209494
rect 136102 209258 136186 209494
rect 136422 209258 136454 209494
rect 135834 209174 136454 209258
rect 135834 208938 135866 209174
rect 136102 208938 136186 209174
rect 136422 208938 136454 209174
rect 135834 173494 136454 208938
rect 135834 173258 135866 173494
rect 136102 173258 136186 173494
rect 136422 173258 136454 173494
rect 135834 173174 136454 173258
rect 135834 172938 135866 173174
rect 136102 172938 136186 173174
rect 136422 172938 136454 173174
rect 135834 137494 136454 172938
rect 135834 137258 135866 137494
rect 136102 137258 136186 137494
rect 136422 137258 136454 137494
rect 135834 137174 136454 137258
rect 135834 136938 135866 137174
rect 136102 136938 136186 137174
rect 136422 136938 136454 137174
rect 43568 115174 43888 115206
rect 43568 114938 43610 115174
rect 43846 114938 43888 115174
rect 43568 114854 43888 114938
rect 43568 114618 43610 114854
rect 43846 114618 43888 114854
rect 43568 114586 43888 114618
rect 74288 115174 74608 115206
rect 74288 114938 74330 115174
rect 74566 114938 74608 115174
rect 74288 114854 74608 114938
rect 74288 114618 74330 114854
rect 74566 114618 74608 114854
rect 74288 114586 74608 114618
rect 105008 115174 105328 115206
rect 105008 114938 105050 115174
rect 105286 114938 105328 115174
rect 105008 114854 105328 114938
rect 105008 114618 105050 114854
rect 105286 114618 105328 114854
rect 105008 114586 105328 114618
rect 28208 111454 28528 111486
rect 28208 111218 28250 111454
rect 28486 111218 28528 111454
rect 28208 111134 28528 111218
rect 28208 110898 28250 111134
rect 28486 110898 28528 111134
rect 28208 110866 28528 110898
rect 58928 111454 59248 111486
rect 58928 111218 58970 111454
rect 59206 111218 59248 111454
rect 58928 111134 59248 111218
rect 58928 110898 58970 111134
rect 59206 110898 59248 111134
rect 58928 110866 59248 110898
rect 89648 111454 89968 111486
rect 89648 111218 89690 111454
rect 89926 111218 89968 111454
rect 89648 111134 89968 111218
rect 89648 110898 89690 111134
rect 89926 110898 89968 111134
rect 89648 110866 89968 110898
rect 120368 111454 120688 111486
rect 120368 111218 120410 111454
rect 120646 111218 120688 111454
rect 120368 111134 120688 111218
rect 120368 110898 120410 111134
rect 120646 110898 120688 111134
rect 120368 110866 120688 110898
rect 24114 97538 24146 97774
rect 24382 97538 24466 97774
rect 24702 97538 24734 97774
rect 24114 97454 24734 97538
rect 24114 97218 24146 97454
rect 24382 97218 24466 97454
rect 24702 97218 24734 97454
rect 24114 61774 24734 97218
rect 135834 101494 136454 136938
rect 135834 101258 135866 101494
rect 136102 101258 136186 101494
rect 136422 101258 136454 101494
rect 135834 101174 136454 101258
rect 135834 100938 135866 101174
rect 136102 100938 136186 101174
rect 136422 100938 136454 101174
rect 43568 79174 43888 79206
rect 43568 78938 43610 79174
rect 43846 78938 43888 79174
rect 43568 78854 43888 78938
rect 43568 78618 43610 78854
rect 43846 78618 43888 78854
rect 43568 78586 43888 78618
rect 74288 79174 74608 79206
rect 74288 78938 74330 79174
rect 74566 78938 74608 79174
rect 74288 78854 74608 78938
rect 74288 78618 74330 78854
rect 74566 78618 74608 78854
rect 74288 78586 74608 78618
rect 105008 79174 105328 79206
rect 105008 78938 105050 79174
rect 105286 78938 105328 79174
rect 105008 78854 105328 78938
rect 105008 78618 105050 78854
rect 105286 78618 105328 78854
rect 105008 78586 105328 78618
rect 28208 75454 28528 75486
rect 28208 75218 28250 75454
rect 28486 75218 28528 75454
rect 28208 75134 28528 75218
rect 28208 74898 28250 75134
rect 28486 74898 28528 75134
rect 28208 74866 28528 74898
rect 58928 75454 59248 75486
rect 58928 75218 58970 75454
rect 59206 75218 59248 75454
rect 58928 75134 59248 75218
rect 58928 74898 58970 75134
rect 59206 74898 59248 75134
rect 58928 74866 59248 74898
rect 89648 75454 89968 75486
rect 89648 75218 89690 75454
rect 89926 75218 89968 75454
rect 89648 75134 89968 75218
rect 89648 74898 89690 75134
rect 89926 74898 89968 75134
rect 89648 74866 89968 74898
rect 120368 75454 120688 75486
rect 120368 75218 120410 75454
rect 120646 75218 120688 75454
rect 120368 75134 120688 75218
rect 120368 74898 120410 75134
rect 120646 74898 120688 75134
rect 120368 74866 120688 74898
rect 24114 61538 24146 61774
rect 24382 61538 24466 61774
rect 24702 61538 24734 61774
rect 24114 61454 24734 61538
rect 24114 61218 24146 61454
rect 24382 61218 24466 61454
rect 24702 61218 24734 61454
rect 24114 25774 24734 61218
rect 135834 65494 136454 100938
rect 135834 65258 135866 65494
rect 136102 65258 136186 65494
rect 136422 65258 136454 65494
rect 135834 65174 136454 65258
rect 135834 64938 135866 65174
rect 136102 64938 136186 65174
rect 136422 64938 136454 65174
rect 43568 43174 43888 43206
rect 43568 42938 43610 43174
rect 43846 42938 43888 43174
rect 43568 42854 43888 42938
rect 43568 42618 43610 42854
rect 43846 42618 43888 42854
rect 43568 42586 43888 42618
rect 74288 43174 74608 43206
rect 74288 42938 74330 43174
rect 74566 42938 74608 43174
rect 74288 42854 74608 42938
rect 74288 42618 74330 42854
rect 74566 42618 74608 42854
rect 74288 42586 74608 42618
rect 105008 43174 105328 43206
rect 105008 42938 105050 43174
rect 105286 42938 105328 43174
rect 105008 42854 105328 42938
rect 105008 42618 105050 42854
rect 105286 42618 105328 42854
rect 105008 42586 105328 42618
rect 28208 39454 28528 39486
rect 28208 39218 28250 39454
rect 28486 39218 28528 39454
rect 28208 39134 28528 39218
rect 28208 38898 28250 39134
rect 28486 38898 28528 39134
rect 28208 38866 28528 38898
rect 58928 39454 59248 39486
rect 58928 39218 58970 39454
rect 59206 39218 59248 39454
rect 58928 39134 59248 39218
rect 58928 38898 58970 39134
rect 59206 38898 59248 39134
rect 58928 38866 59248 38898
rect 89648 39454 89968 39486
rect 89648 39218 89690 39454
rect 89926 39218 89968 39454
rect 89648 39134 89968 39218
rect 89648 38898 89690 39134
rect 89926 38898 89968 39134
rect 89648 38866 89968 38898
rect 120368 39454 120688 39486
rect 120368 39218 120410 39454
rect 120646 39218 120688 39454
rect 120368 39134 120688 39218
rect 120368 38898 120410 39134
rect 120646 38898 120688 39134
rect 120368 38866 120688 38898
rect 24114 25538 24146 25774
rect 24382 25538 24466 25774
rect 24702 25538 24734 25774
rect 24114 25454 24734 25538
rect 24114 25218 24146 25454
rect 24382 25218 24466 25454
rect 24702 25218 24734 25454
rect 24114 -6106 24734 25218
rect 135834 29494 136454 64938
rect 135834 29258 135866 29494
rect 136102 29258 136186 29494
rect 136422 29258 136454 29494
rect 135834 29174 136454 29258
rect 135834 28938 135866 29174
rect 136102 28938 136186 29174
rect 136422 28938 136454 29174
rect 24114 -6342 24146 -6106
rect 24382 -6342 24466 -6106
rect 24702 -6342 24734 -6106
rect 24114 -6426 24734 -6342
rect 24114 -6662 24146 -6426
rect 24382 -6662 24466 -6426
rect 24702 -6662 24734 -6426
rect 24114 -7654 24734 -6662
rect 37794 3454 38414 24559
rect 37794 3218 37826 3454
rect 38062 3218 38146 3454
rect 38382 3218 38414 3454
rect 37794 3134 38414 3218
rect 37794 2898 37826 3134
rect 38062 2898 38146 3134
rect 38382 2898 38414 3134
rect 37794 -346 38414 2898
rect 37794 -582 37826 -346
rect 38062 -582 38146 -346
rect 38382 -582 38414 -346
rect 37794 -666 38414 -582
rect 37794 -902 37826 -666
rect 38062 -902 38146 -666
rect 38382 -902 38414 -666
rect 37794 -7654 38414 -902
rect 41514 7174 42134 24559
rect 41514 6938 41546 7174
rect 41782 6938 41866 7174
rect 42102 6938 42134 7174
rect 41514 6854 42134 6938
rect 41514 6618 41546 6854
rect 41782 6618 41866 6854
rect 42102 6618 42134 6854
rect 41514 -1306 42134 6618
rect 41514 -1542 41546 -1306
rect 41782 -1542 41866 -1306
rect 42102 -1542 42134 -1306
rect 41514 -1626 42134 -1542
rect 41514 -1862 41546 -1626
rect 41782 -1862 41866 -1626
rect 42102 -1862 42134 -1626
rect 41514 -7654 42134 -1862
rect 45234 10894 45854 24559
rect 45234 10658 45266 10894
rect 45502 10658 45586 10894
rect 45822 10658 45854 10894
rect 45234 10574 45854 10658
rect 45234 10338 45266 10574
rect 45502 10338 45586 10574
rect 45822 10338 45854 10574
rect 45234 -2266 45854 10338
rect 45234 -2502 45266 -2266
rect 45502 -2502 45586 -2266
rect 45822 -2502 45854 -2266
rect 45234 -2586 45854 -2502
rect 45234 -2822 45266 -2586
rect 45502 -2822 45586 -2586
rect 45822 -2822 45854 -2586
rect 45234 -7654 45854 -2822
rect 48954 14614 49574 24559
rect 48954 14378 48986 14614
rect 49222 14378 49306 14614
rect 49542 14378 49574 14614
rect 48954 14294 49574 14378
rect 48954 14058 48986 14294
rect 49222 14058 49306 14294
rect 49542 14058 49574 14294
rect 48954 -3226 49574 14058
rect 48954 -3462 48986 -3226
rect 49222 -3462 49306 -3226
rect 49542 -3462 49574 -3226
rect 48954 -3546 49574 -3462
rect 48954 -3782 48986 -3546
rect 49222 -3782 49306 -3546
rect 49542 -3782 49574 -3546
rect 48954 -7654 49574 -3782
rect 52674 18334 53294 24559
rect 52674 18098 52706 18334
rect 52942 18098 53026 18334
rect 53262 18098 53294 18334
rect 52674 18014 53294 18098
rect 52674 17778 52706 18014
rect 52942 17778 53026 18014
rect 53262 17778 53294 18014
rect 52674 -4186 53294 17778
rect 52674 -4422 52706 -4186
rect 52942 -4422 53026 -4186
rect 53262 -4422 53294 -4186
rect 52674 -4506 53294 -4422
rect 52674 -4742 52706 -4506
rect 52942 -4742 53026 -4506
rect 53262 -4742 53294 -4506
rect 52674 -7654 53294 -4742
rect 56394 22054 57014 24559
rect 56394 21818 56426 22054
rect 56662 21818 56746 22054
rect 56982 21818 57014 22054
rect 56394 21734 57014 21818
rect 56394 21498 56426 21734
rect 56662 21498 56746 21734
rect 56982 21498 57014 21734
rect 56394 -5146 57014 21498
rect 56394 -5382 56426 -5146
rect 56662 -5382 56746 -5146
rect 56982 -5382 57014 -5146
rect 56394 -5466 57014 -5382
rect 56394 -5702 56426 -5466
rect 56662 -5702 56746 -5466
rect 56982 -5702 57014 -5466
rect 56394 -7654 57014 -5702
rect 73794 3454 74414 24068
rect 73794 3218 73826 3454
rect 74062 3218 74146 3454
rect 74382 3218 74414 3454
rect 73794 3134 74414 3218
rect 73794 2898 73826 3134
rect 74062 2898 74146 3134
rect 74382 2898 74414 3134
rect 73794 -346 74414 2898
rect 73794 -582 73826 -346
rect 74062 -582 74146 -346
rect 74382 -582 74414 -346
rect 73794 -666 74414 -582
rect 73794 -902 73826 -666
rect 74062 -902 74146 -666
rect 74382 -902 74414 -666
rect 73794 -7654 74414 -902
rect 77514 7174 78134 24559
rect 77514 6938 77546 7174
rect 77782 6938 77866 7174
rect 78102 6938 78134 7174
rect 77514 6854 78134 6938
rect 77514 6618 77546 6854
rect 77782 6618 77866 6854
rect 78102 6618 78134 6854
rect 77514 -1306 78134 6618
rect 77514 -1542 77546 -1306
rect 77782 -1542 77866 -1306
rect 78102 -1542 78134 -1306
rect 77514 -1626 78134 -1542
rect 77514 -1862 77546 -1626
rect 77782 -1862 77866 -1626
rect 78102 -1862 78134 -1626
rect 77514 -7654 78134 -1862
rect 81234 10894 81854 24559
rect 81234 10658 81266 10894
rect 81502 10658 81586 10894
rect 81822 10658 81854 10894
rect 81234 10574 81854 10658
rect 81234 10338 81266 10574
rect 81502 10338 81586 10574
rect 81822 10338 81854 10574
rect 81234 -2266 81854 10338
rect 81234 -2502 81266 -2266
rect 81502 -2502 81586 -2266
rect 81822 -2502 81854 -2266
rect 81234 -2586 81854 -2502
rect 81234 -2822 81266 -2586
rect 81502 -2822 81586 -2586
rect 81822 -2822 81854 -2586
rect 81234 -7654 81854 -2822
rect 84954 14614 85574 24559
rect 84954 14378 84986 14614
rect 85222 14378 85306 14614
rect 85542 14378 85574 14614
rect 84954 14294 85574 14378
rect 84954 14058 84986 14294
rect 85222 14058 85306 14294
rect 85542 14058 85574 14294
rect 84954 -3226 85574 14058
rect 84954 -3462 84986 -3226
rect 85222 -3462 85306 -3226
rect 85542 -3462 85574 -3226
rect 84954 -3546 85574 -3462
rect 84954 -3782 84986 -3546
rect 85222 -3782 85306 -3546
rect 85542 -3782 85574 -3546
rect 84954 -7654 85574 -3782
rect 88674 18334 89294 24559
rect 88674 18098 88706 18334
rect 88942 18098 89026 18334
rect 89262 18098 89294 18334
rect 88674 18014 89294 18098
rect 88674 17778 88706 18014
rect 88942 17778 89026 18014
rect 89262 17778 89294 18014
rect 88674 -4186 89294 17778
rect 88674 -4422 88706 -4186
rect 88942 -4422 89026 -4186
rect 89262 -4422 89294 -4186
rect 88674 -4506 89294 -4422
rect 88674 -4742 88706 -4506
rect 88942 -4742 89026 -4506
rect 89262 -4742 89294 -4506
rect 88674 -7654 89294 -4742
rect 92394 22054 93014 24559
rect 92394 21818 92426 22054
rect 92662 21818 92746 22054
rect 92982 21818 93014 22054
rect 92394 21734 93014 21818
rect 92394 21498 92426 21734
rect 92662 21498 92746 21734
rect 92982 21498 93014 21734
rect 92394 -5146 93014 21498
rect 92394 -5382 92426 -5146
rect 92662 -5382 92746 -5146
rect 92982 -5382 93014 -5146
rect 92394 -5466 93014 -5382
rect 92394 -5702 92426 -5466
rect 92662 -5702 92746 -5466
rect 92982 -5702 93014 -5466
rect 92394 -7654 93014 -5702
rect 109794 3454 110414 24559
rect 109794 3218 109826 3454
rect 110062 3218 110146 3454
rect 110382 3218 110414 3454
rect 109794 3134 110414 3218
rect 109794 2898 109826 3134
rect 110062 2898 110146 3134
rect 110382 2898 110414 3134
rect 109794 -346 110414 2898
rect 109794 -582 109826 -346
rect 110062 -582 110146 -346
rect 110382 -582 110414 -346
rect 109794 -666 110414 -582
rect 109794 -902 109826 -666
rect 110062 -902 110146 -666
rect 110382 -902 110414 -666
rect 109794 -7654 110414 -902
rect 113514 7174 114134 24559
rect 113514 6938 113546 7174
rect 113782 6938 113866 7174
rect 114102 6938 114134 7174
rect 113514 6854 114134 6938
rect 113514 6618 113546 6854
rect 113782 6618 113866 6854
rect 114102 6618 114134 6854
rect 113514 -1306 114134 6618
rect 113514 -1542 113546 -1306
rect 113782 -1542 113866 -1306
rect 114102 -1542 114134 -1306
rect 113514 -1626 114134 -1542
rect 113514 -1862 113546 -1626
rect 113782 -1862 113866 -1626
rect 114102 -1862 114134 -1626
rect 113514 -7654 114134 -1862
rect 117234 10894 117854 24559
rect 117234 10658 117266 10894
rect 117502 10658 117586 10894
rect 117822 10658 117854 10894
rect 117234 10574 117854 10658
rect 117234 10338 117266 10574
rect 117502 10338 117586 10574
rect 117822 10338 117854 10574
rect 117234 -2266 117854 10338
rect 117234 -2502 117266 -2266
rect 117502 -2502 117586 -2266
rect 117822 -2502 117854 -2266
rect 117234 -2586 117854 -2502
rect 117234 -2822 117266 -2586
rect 117502 -2822 117586 -2586
rect 117822 -2822 117854 -2586
rect 117234 -7654 117854 -2822
rect 120954 14614 121574 24559
rect 120954 14378 120986 14614
rect 121222 14378 121306 14614
rect 121542 14378 121574 14614
rect 120954 14294 121574 14378
rect 120954 14058 120986 14294
rect 121222 14058 121306 14294
rect 121542 14058 121574 14294
rect 120954 -3226 121574 14058
rect 120954 -3462 120986 -3226
rect 121222 -3462 121306 -3226
rect 121542 -3462 121574 -3226
rect 120954 -3546 121574 -3462
rect 120954 -3782 120986 -3546
rect 121222 -3782 121306 -3546
rect 121542 -3782 121574 -3546
rect 120954 -7654 121574 -3782
rect 124674 18334 125294 24559
rect 124674 18098 124706 18334
rect 124942 18098 125026 18334
rect 125262 18098 125294 18334
rect 124674 18014 125294 18098
rect 124674 17778 124706 18014
rect 124942 17778 125026 18014
rect 125262 17778 125294 18014
rect 124674 -4186 125294 17778
rect 124674 -4422 124706 -4186
rect 124942 -4422 125026 -4186
rect 125262 -4422 125294 -4186
rect 124674 -4506 125294 -4422
rect 124674 -4742 124706 -4506
rect 124942 -4742 125026 -4506
rect 125262 -4742 125294 -4506
rect 124674 -7654 125294 -4742
rect 128394 22054 129014 24559
rect 128394 21818 128426 22054
rect 128662 21818 128746 22054
rect 128982 21818 129014 22054
rect 128394 21734 129014 21818
rect 128394 21498 128426 21734
rect 128662 21498 128746 21734
rect 128982 21498 129014 21734
rect 128394 -5146 129014 21498
rect 128394 -5382 128426 -5146
rect 128662 -5382 128746 -5146
rect 128982 -5382 129014 -5146
rect 128394 -5466 129014 -5382
rect 128394 -5702 128426 -5466
rect 128662 -5702 128746 -5466
rect 128982 -5702 129014 -5466
rect 128394 -7654 129014 -5702
rect 135834 -7066 136454 28938
rect 135834 -7302 135866 -7066
rect 136102 -7302 136186 -7066
rect 136422 -7302 136454 -7066
rect 135834 -7386 136454 -7302
rect 135834 -7622 135866 -7386
rect 136102 -7622 136186 -7386
rect 136422 -7622 136454 -7386
rect 135834 -7654 136454 -7622
rect 145794 704838 146414 711590
rect 145794 704602 145826 704838
rect 146062 704602 146146 704838
rect 146382 704602 146414 704838
rect 145794 704518 146414 704602
rect 145794 704282 145826 704518
rect 146062 704282 146146 704518
rect 146382 704282 146414 704518
rect 145794 687454 146414 704282
rect 145794 687218 145826 687454
rect 146062 687218 146146 687454
rect 146382 687218 146414 687454
rect 145794 687134 146414 687218
rect 145794 686898 145826 687134
rect 146062 686898 146146 687134
rect 146382 686898 146414 687134
rect 145794 651454 146414 686898
rect 145794 651218 145826 651454
rect 146062 651218 146146 651454
rect 146382 651218 146414 651454
rect 145794 651134 146414 651218
rect 145794 650898 145826 651134
rect 146062 650898 146146 651134
rect 146382 650898 146414 651134
rect 145794 615454 146414 650898
rect 145794 615218 145826 615454
rect 146062 615218 146146 615454
rect 146382 615218 146414 615454
rect 145794 615134 146414 615218
rect 145794 614898 145826 615134
rect 146062 614898 146146 615134
rect 146382 614898 146414 615134
rect 145794 579454 146414 614898
rect 145794 579218 145826 579454
rect 146062 579218 146146 579454
rect 146382 579218 146414 579454
rect 145794 579134 146414 579218
rect 145794 578898 145826 579134
rect 146062 578898 146146 579134
rect 146382 578898 146414 579134
rect 145794 543454 146414 578898
rect 145794 543218 145826 543454
rect 146062 543218 146146 543454
rect 146382 543218 146414 543454
rect 145794 543134 146414 543218
rect 145794 542898 145826 543134
rect 146062 542898 146146 543134
rect 146382 542898 146414 543134
rect 145794 507454 146414 542898
rect 145794 507218 145826 507454
rect 146062 507218 146146 507454
rect 146382 507218 146414 507454
rect 145794 507134 146414 507218
rect 145794 506898 145826 507134
rect 146062 506898 146146 507134
rect 146382 506898 146414 507134
rect 145794 471454 146414 506898
rect 145794 471218 145826 471454
rect 146062 471218 146146 471454
rect 146382 471218 146414 471454
rect 145794 471134 146414 471218
rect 145794 470898 145826 471134
rect 146062 470898 146146 471134
rect 146382 470898 146414 471134
rect 145794 435454 146414 470898
rect 145794 435218 145826 435454
rect 146062 435218 146146 435454
rect 146382 435218 146414 435454
rect 145794 435134 146414 435218
rect 145794 434898 145826 435134
rect 146062 434898 146146 435134
rect 146382 434898 146414 435134
rect 145794 399454 146414 434898
rect 145794 399218 145826 399454
rect 146062 399218 146146 399454
rect 146382 399218 146414 399454
rect 145794 399134 146414 399218
rect 145794 398898 145826 399134
rect 146062 398898 146146 399134
rect 146382 398898 146414 399134
rect 145794 363454 146414 398898
rect 145794 363218 145826 363454
rect 146062 363218 146146 363454
rect 146382 363218 146414 363454
rect 145794 363134 146414 363218
rect 145794 362898 145826 363134
rect 146062 362898 146146 363134
rect 146382 362898 146414 363134
rect 145794 327454 146414 362898
rect 145794 327218 145826 327454
rect 146062 327218 146146 327454
rect 146382 327218 146414 327454
rect 145794 327134 146414 327218
rect 145794 326898 145826 327134
rect 146062 326898 146146 327134
rect 146382 326898 146414 327134
rect 145794 291454 146414 326898
rect 145794 291218 145826 291454
rect 146062 291218 146146 291454
rect 146382 291218 146414 291454
rect 145794 291134 146414 291218
rect 145794 290898 145826 291134
rect 146062 290898 146146 291134
rect 146382 290898 146414 291134
rect 145794 255454 146414 290898
rect 145794 255218 145826 255454
rect 146062 255218 146146 255454
rect 146382 255218 146414 255454
rect 145794 255134 146414 255218
rect 145794 254898 145826 255134
rect 146062 254898 146146 255134
rect 146382 254898 146414 255134
rect 145794 219454 146414 254898
rect 145794 219218 145826 219454
rect 146062 219218 146146 219454
rect 146382 219218 146414 219454
rect 145794 219134 146414 219218
rect 145794 218898 145826 219134
rect 146062 218898 146146 219134
rect 146382 218898 146414 219134
rect 145794 183454 146414 218898
rect 145794 183218 145826 183454
rect 146062 183218 146146 183454
rect 146382 183218 146414 183454
rect 145794 183134 146414 183218
rect 145794 182898 145826 183134
rect 146062 182898 146146 183134
rect 146382 182898 146414 183134
rect 145794 147454 146414 182898
rect 145794 147218 145826 147454
rect 146062 147218 146146 147454
rect 146382 147218 146414 147454
rect 145794 147134 146414 147218
rect 145794 146898 145826 147134
rect 146062 146898 146146 147134
rect 146382 146898 146414 147134
rect 145794 111454 146414 146898
rect 145794 111218 145826 111454
rect 146062 111218 146146 111454
rect 146382 111218 146414 111454
rect 145794 111134 146414 111218
rect 145794 110898 145826 111134
rect 146062 110898 146146 111134
rect 146382 110898 146414 111134
rect 145794 75454 146414 110898
rect 145794 75218 145826 75454
rect 146062 75218 146146 75454
rect 146382 75218 146414 75454
rect 145794 75134 146414 75218
rect 145794 74898 145826 75134
rect 146062 74898 146146 75134
rect 146382 74898 146414 75134
rect 145794 39454 146414 74898
rect 145794 39218 145826 39454
rect 146062 39218 146146 39454
rect 146382 39218 146414 39454
rect 145794 39134 146414 39218
rect 145794 38898 145826 39134
rect 146062 38898 146146 39134
rect 146382 38898 146414 39134
rect 145794 3454 146414 38898
rect 145794 3218 145826 3454
rect 146062 3218 146146 3454
rect 146382 3218 146414 3454
rect 145794 3134 146414 3218
rect 145794 2898 145826 3134
rect 146062 2898 146146 3134
rect 146382 2898 146414 3134
rect 145794 -346 146414 2898
rect 145794 -582 145826 -346
rect 146062 -582 146146 -346
rect 146382 -582 146414 -346
rect 145794 -666 146414 -582
rect 145794 -902 145826 -666
rect 146062 -902 146146 -666
rect 146382 -902 146414 -666
rect 145794 -7654 146414 -902
rect 149514 705798 150134 711590
rect 149514 705562 149546 705798
rect 149782 705562 149866 705798
rect 150102 705562 150134 705798
rect 149514 705478 150134 705562
rect 149514 705242 149546 705478
rect 149782 705242 149866 705478
rect 150102 705242 150134 705478
rect 149514 691174 150134 705242
rect 149514 690938 149546 691174
rect 149782 690938 149866 691174
rect 150102 690938 150134 691174
rect 149514 690854 150134 690938
rect 149514 690618 149546 690854
rect 149782 690618 149866 690854
rect 150102 690618 150134 690854
rect 149514 655174 150134 690618
rect 149514 654938 149546 655174
rect 149782 654938 149866 655174
rect 150102 654938 150134 655174
rect 149514 654854 150134 654938
rect 149514 654618 149546 654854
rect 149782 654618 149866 654854
rect 150102 654618 150134 654854
rect 149514 619174 150134 654618
rect 149514 618938 149546 619174
rect 149782 618938 149866 619174
rect 150102 618938 150134 619174
rect 149514 618854 150134 618938
rect 149514 618618 149546 618854
rect 149782 618618 149866 618854
rect 150102 618618 150134 618854
rect 149514 583174 150134 618618
rect 149514 582938 149546 583174
rect 149782 582938 149866 583174
rect 150102 582938 150134 583174
rect 149514 582854 150134 582938
rect 149514 582618 149546 582854
rect 149782 582618 149866 582854
rect 150102 582618 150134 582854
rect 149514 547174 150134 582618
rect 149514 546938 149546 547174
rect 149782 546938 149866 547174
rect 150102 546938 150134 547174
rect 149514 546854 150134 546938
rect 149514 546618 149546 546854
rect 149782 546618 149866 546854
rect 150102 546618 150134 546854
rect 149514 511174 150134 546618
rect 149514 510938 149546 511174
rect 149782 510938 149866 511174
rect 150102 510938 150134 511174
rect 149514 510854 150134 510938
rect 149514 510618 149546 510854
rect 149782 510618 149866 510854
rect 150102 510618 150134 510854
rect 149514 475174 150134 510618
rect 149514 474938 149546 475174
rect 149782 474938 149866 475174
rect 150102 474938 150134 475174
rect 149514 474854 150134 474938
rect 149514 474618 149546 474854
rect 149782 474618 149866 474854
rect 150102 474618 150134 474854
rect 149514 439174 150134 474618
rect 149514 438938 149546 439174
rect 149782 438938 149866 439174
rect 150102 438938 150134 439174
rect 149514 438854 150134 438938
rect 149514 438618 149546 438854
rect 149782 438618 149866 438854
rect 150102 438618 150134 438854
rect 149514 403174 150134 438618
rect 149514 402938 149546 403174
rect 149782 402938 149866 403174
rect 150102 402938 150134 403174
rect 149514 402854 150134 402938
rect 149514 402618 149546 402854
rect 149782 402618 149866 402854
rect 150102 402618 150134 402854
rect 149514 367174 150134 402618
rect 149514 366938 149546 367174
rect 149782 366938 149866 367174
rect 150102 366938 150134 367174
rect 149514 366854 150134 366938
rect 149514 366618 149546 366854
rect 149782 366618 149866 366854
rect 150102 366618 150134 366854
rect 149514 331174 150134 366618
rect 149514 330938 149546 331174
rect 149782 330938 149866 331174
rect 150102 330938 150134 331174
rect 149514 330854 150134 330938
rect 149514 330618 149546 330854
rect 149782 330618 149866 330854
rect 150102 330618 150134 330854
rect 149514 295174 150134 330618
rect 149514 294938 149546 295174
rect 149782 294938 149866 295174
rect 150102 294938 150134 295174
rect 149514 294854 150134 294938
rect 149514 294618 149546 294854
rect 149782 294618 149866 294854
rect 150102 294618 150134 294854
rect 149514 259174 150134 294618
rect 149514 258938 149546 259174
rect 149782 258938 149866 259174
rect 150102 258938 150134 259174
rect 149514 258854 150134 258938
rect 149514 258618 149546 258854
rect 149782 258618 149866 258854
rect 150102 258618 150134 258854
rect 149514 223174 150134 258618
rect 149514 222938 149546 223174
rect 149782 222938 149866 223174
rect 150102 222938 150134 223174
rect 149514 222854 150134 222938
rect 149514 222618 149546 222854
rect 149782 222618 149866 222854
rect 150102 222618 150134 222854
rect 149514 187174 150134 222618
rect 149514 186938 149546 187174
rect 149782 186938 149866 187174
rect 150102 186938 150134 187174
rect 149514 186854 150134 186938
rect 149514 186618 149546 186854
rect 149782 186618 149866 186854
rect 150102 186618 150134 186854
rect 149514 151174 150134 186618
rect 149514 150938 149546 151174
rect 149782 150938 149866 151174
rect 150102 150938 150134 151174
rect 149514 150854 150134 150938
rect 149514 150618 149546 150854
rect 149782 150618 149866 150854
rect 150102 150618 150134 150854
rect 149514 115174 150134 150618
rect 149514 114938 149546 115174
rect 149782 114938 149866 115174
rect 150102 114938 150134 115174
rect 149514 114854 150134 114938
rect 149514 114618 149546 114854
rect 149782 114618 149866 114854
rect 150102 114618 150134 114854
rect 149514 79174 150134 114618
rect 149514 78938 149546 79174
rect 149782 78938 149866 79174
rect 150102 78938 150134 79174
rect 149514 78854 150134 78938
rect 149514 78618 149546 78854
rect 149782 78618 149866 78854
rect 150102 78618 150134 78854
rect 149514 43174 150134 78618
rect 149514 42938 149546 43174
rect 149782 42938 149866 43174
rect 150102 42938 150134 43174
rect 149514 42854 150134 42938
rect 149514 42618 149546 42854
rect 149782 42618 149866 42854
rect 150102 42618 150134 42854
rect 149514 7174 150134 42618
rect 149514 6938 149546 7174
rect 149782 6938 149866 7174
rect 150102 6938 150134 7174
rect 149514 6854 150134 6938
rect 149514 6618 149546 6854
rect 149782 6618 149866 6854
rect 150102 6618 150134 6854
rect 149514 -1306 150134 6618
rect 149514 -1542 149546 -1306
rect 149782 -1542 149866 -1306
rect 150102 -1542 150134 -1306
rect 149514 -1626 150134 -1542
rect 149514 -1862 149546 -1626
rect 149782 -1862 149866 -1626
rect 150102 -1862 150134 -1626
rect 149514 -7654 150134 -1862
rect 153234 706758 153854 711590
rect 153234 706522 153266 706758
rect 153502 706522 153586 706758
rect 153822 706522 153854 706758
rect 153234 706438 153854 706522
rect 153234 706202 153266 706438
rect 153502 706202 153586 706438
rect 153822 706202 153854 706438
rect 153234 694894 153854 706202
rect 153234 694658 153266 694894
rect 153502 694658 153586 694894
rect 153822 694658 153854 694894
rect 153234 694574 153854 694658
rect 153234 694338 153266 694574
rect 153502 694338 153586 694574
rect 153822 694338 153854 694574
rect 153234 658894 153854 694338
rect 153234 658658 153266 658894
rect 153502 658658 153586 658894
rect 153822 658658 153854 658894
rect 153234 658574 153854 658658
rect 153234 658338 153266 658574
rect 153502 658338 153586 658574
rect 153822 658338 153854 658574
rect 153234 622894 153854 658338
rect 153234 622658 153266 622894
rect 153502 622658 153586 622894
rect 153822 622658 153854 622894
rect 153234 622574 153854 622658
rect 153234 622338 153266 622574
rect 153502 622338 153586 622574
rect 153822 622338 153854 622574
rect 153234 586894 153854 622338
rect 153234 586658 153266 586894
rect 153502 586658 153586 586894
rect 153822 586658 153854 586894
rect 153234 586574 153854 586658
rect 153234 586338 153266 586574
rect 153502 586338 153586 586574
rect 153822 586338 153854 586574
rect 153234 550894 153854 586338
rect 153234 550658 153266 550894
rect 153502 550658 153586 550894
rect 153822 550658 153854 550894
rect 153234 550574 153854 550658
rect 153234 550338 153266 550574
rect 153502 550338 153586 550574
rect 153822 550338 153854 550574
rect 153234 514894 153854 550338
rect 153234 514658 153266 514894
rect 153502 514658 153586 514894
rect 153822 514658 153854 514894
rect 153234 514574 153854 514658
rect 153234 514338 153266 514574
rect 153502 514338 153586 514574
rect 153822 514338 153854 514574
rect 153234 478894 153854 514338
rect 153234 478658 153266 478894
rect 153502 478658 153586 478894
rect 153822 478658 153854 478894
rect 153234 478574 153854 478658
rect 153234 478338 153266 478574
rect 153502 478338 153586 478574
rect 153822 478338 153854 478574
rect 153234 442894 153854 478338
rect 153234 442658 153266 442894
rect 153502 442658 153586 442894
rect 153822 442658 153854 442894
rect 153234 442574 153854 442658
rect 153234 442338 153266 442574
rect 153502 442338 153586 442574
rect 153822 442338 153854 442574
rect 153234 406894 153854 442338
rect 156954 707718 157574 711590
rect 156954 707482 156986 707718
rect 157222 707482 157306 707718
rect 157542 707482 157574 707718
rect 156954 707398 157574 707482
rect 156954 707162 156986 707398
rect 157222 707162 157306 707398
rect 157542 707162 157574 707398
rect 156954 698614 157574 707162
rect 156954 698378 156986 698614
rect 157222 698378 157306 698614
rect 157542 698378 157574 698614
rect 156954 698294 157574 698378
rect 156954 698058 156986 698294
rect 157222 698058 157306 698294
rect 157542 698058 157574 698294
rect 156954 662614 157574 698058
rect 156954 662378 156986 662614
rect 157222 662378 157306 662614
rect 157542 662378 157574 662614
rect 156954 662294 157574 662378
rect 156954 662058 156986 662294
rect 157222 662058 157306 662294
rect 157542 662058 157574 662294
rect 156954 626614 157574 662058
rect 156954 626378 156986 626614
rect 157222 626378 157306 626614
rect 157542 626378 157574 626614
rect 156954 626294 157574 626378
rect 156954 626058 156986 626294
rect 157222 626058 157306 626294
rect 157542 626058 157574 626294
rect 156954 590614 157574 626058
rect 156954 590378 156986 590614
rect 157222 590378 157306 590614
rect 157542 590378 157574 590614
rect 156954 590294 157574 590378
rect 156954 590058 156986 590294
rect 157222 590058 157306 590294
rect 157542 590058 157574 590294
rect 156954 554614 157574 590058
rect 156954 554378 156986 554614
rect 157222 554378 157306 554614
rect 157542 554378 157574 554614
rect 156954 554294 157574 554378
rect 156954 554058 156986 554294
rect 157222 554058 157306 554294
rect 157542 554058 157574 554294
rect 156954 518614 157574 554058
rect 156954 518378 156986 518614
rect 157222 518378 157306 518614
rect 157542 518378 157574 518614
rect 156954 518294 157574 518378
rect 156954 518058 156986 518294
rect 157222 518058 157306 518294
rect 157542 518058 157574 518294
rect 156954 482614 157574 518058
rect 156954 482378 156986 482614
rect 157222 482378 157306 482614
rect 157542 482378 157574 482614
rect 156954 482294 157574 482378
rect 156954 482058 156986 482294
rect 157222 482058 157306 482294
rect 157542 482058 157574 482294
rect 156954 446614 157574 482058
rect 156954 446378 156986 446614
rect 157222 446378 157306 446614
rect 157542 446378 157574 446614
rect 156954 446294 157574 446378
rect 156954 446058 156986 446294
rect 157222 446058 157306 446294
rect 157542 446058 157574 446294
rect 156954 423529 157574 446058
rect 160674 708678 161294 711590
rect 160674 708442 160706 708678
rect 160942 708442 161026 708678
rect 161262 708442 161294 708678
rect 160674 708358 161294 708442
rect 160674 708122 160706 708358
rect 160942 708122 161026 708358
rect 161262 708122 161294 708358
rect 160674 666334 161294 708122
rect 160674 666098 160706 666334
rect 160942 666098 161026 666334
rect 161262 666098 161294 666334
rect 160674 666014 161294 666098
rect 160674 665778 160706 666014
rect 160942 665778 161026 666014
rect 161262 665778 161294 666014
rect 160674 630334 161294 665778
rect 160674 630098 160706 630334
rect 160942 630098 161026 630334
rect 161262 630098 161294 630334
rect 160674 630014 161294 630098
rect 160674 629778 160706 630014
rect 160942 629778 161026 630014
rect 161262 629778 161294 630014
rect 160674 594334 161294 629778
rect 160674 594098 160706 594334
rect 160942 594098 161026 594334
rect 161262 594098 161294 594334
rect 160674 594014 161294 594098
rect 160674 593778 160706 594014
rect 160942 593778 161026 594014
rect 161262 593778 161294 594014
rect 160674 558334 161294 593778
rect 160674 558098 160706 558334
rect 160942 558098 161026 558334
rect 161262 558098 161294 558334
rect 160674 558014 161294 558098
rect 160674 557778 160706 558014
rect 160942 557778 161026 558014
rect 161262 557778 161294 558014
rect 160674 522334 161294 557778
rect 160674 522098 160706 522334
rect 160942 522098 161026 522334
rect 161262 522098 161294 522334
rect 160674 522014 161294 522098
rect 160674 521778 160706 522014
rect 160942 521778 161026 522014
rect 161262 521778 161294 522014
rect 160674 486334 161294 521778
rect 160674 486098 160706 486334
rect 160942 486098 161026 486334
rect 161262 486098 161294 486334
rect 160674 486014 161294 486098
rect 160674 485778 160706 486014
rect 160942 485778 161026 486014
rect 161262 485778 161294 486014
rect 160674 450334 161294 485778
rect 160674 450098 160706 450334
rect 160942 450098 161026 450334
rect 161262 450098 161294 450334
rect 160674 450014 161294 450098
rect 160674 449778 160706 450014
rect 160942 449778 161026 450014
rect 161262 449778 161294 450014
rect 160674 423529 161294 449778
rect 164394 709638 165014 711590
rect 164394 709402 164426 709638
rect 164662 709402 164746 709638
rect 164982 709402 165014 709638
rect 164394 709318 165014 709402
rect 164394 709082 164426 709318
rect 164662 709082 164746 709318
rect 164982 709082 165014 709318
rect 164394 670054 165014 709082
rect 164394 669818 164426 670054
rect 164662 669818 164746 670054
rect 164982 669818 165014 670054
rect 164394 669734 165014 669818
rect 164394 669498 164426 669734
rect 164662 669498 164746 669734
rect 164982 669498 165014 669734
rect 164394 634054 165014 669498
rect 164394 633818 164426 634054
rect 164662 633818 164746 634054
rect 164982 633818 165014 634054
rect 164394 633734 165014 633818
rect 164394 633498 164426 633734
rect 164662 633498 164746 633734
rect 164982 633498 165014 633734
rect 164394 598054 165014 633498
rect 164394 597818 164426 598054
rect 164662 597818 164746 598054
rect 164982 597818 165014 598054
rect 164394 597734 165014 597818
rect 164394 597498 164426 597734
rect 164662 597498 164746 597734
rect 164982 597498 165014 597734
rect 164394 562054 165014 597498
rect 164394 561818 164426 562054
rect 164662 561818 164746 562054
rect 164982 561818 165014 562054
rect 164394 561734 165014 561818
rect 164394 561498 164426 561734
rect 164662 561498 164746 561734
rect 164982 561498 165014 561734
rect 164394 526054 165014 561498
rect 164394 525818 164426 526054
rect 164662 525818 164746 526054
rect 164982 525818 165014 526054
rect 164394 525734 165014 525818
rect 164394 525498 164426 525734
rect 164662 525498 164746 525734
rect 164982 525498 165014 525734
rect 164394 490054 165014 525498
rect 164394 489818 164426 490054
rect 164662 489818 164746 490054
rect 164982 489818 165014 490054
rect 164394 489734 165014 489818
rect 164394 489498 164426 489734
rect 164662 489498 164746 489734
rect 164982 489498 165014 489734
rect 164394 454054 165014 489498
rect 164394 453818 164426 454054
rect 164662 453818 164746 454054
rect 164982 453818 165014 454054
rect 164394 453734 165014 453818
rect 164394 453498 164426 453734
rect 164662 453498 164746 453734
rect 164982 453498 165014 453734
rect 164394 423529 165014 453498
rect 168114 710598 168734 711590
rect 168114 710362 168146 710598
rect 168382 710362 168466 710598
rect 168702 710362 168734 710598
rect 168114 710278 168734 710362
rect 168114 710042 168146 710278
rect 168382 710042 168466 710278
rect 168702 710042 168734 710278
rect 168114 673774 168734 710042
rect 168114 673538 168146 673774
rect 168382 673538 168466 673774
rect 168702 673538 168734 673774
rect 168114 673454 168734 673538
rect 168114 673218 168146 673454
rect 168382 673218 168466 673454
rect 168702 673218 168734 673454
rect 168114 637774 168734 673218
rect 168114 637538 168146 637774
rect 168382 637538 168466 637774
rect 168702 637538 168734 637774
rect 168114 637454 168734 637538
rect 168114 637218 168146 637454
rect 168382 637218 168466 637454
rect 168702 637218 168734 637454
rect 168114 601774 168734 637218
rect 168114 601538 168146 601774
rect 168382 601538 168466 601774
rect 168702 601538 168734 601774
rect 168114 601454 168734 601538
rect 168114 601218 168146 601454
rect 168382 601218 168466 601454
rect 168702 601218 168734 601454
rect 168114 565774 168734 601218
rect 168114 565538 168146 565774
rect 168382 565538 168466 565774
rect 168702 565538 168734 565774
rect 168114 565454 168734 565538
rect 168114 565218 168146 565454
rect 168382 565218 168466 565454
rect 168702 565218 168734 565454
rect 168114 529774 168734 565218
rect 168114 529538 168146 529774
rect 168382 529538 168466 529774
rect 168702 529538 168734 529774
rect 168114 529454 168734 529538
rect 168114 529218 168146 529454
rect 168382 529218 168466 529454
rect 168702 529218 168734 529454
rect 168114 493774 168734 529218
rect 168114 493538 168146 493774
rect 168382 493538 168466 493774
rect 168702 493538 168734 493774
rect 168114 493454 168734 493538
rect 168114 493218 168146 493454
rect 168382 493218 168466 493454
rect 168702 493218 168734 493454
rect 168114 457774 168734 493218
rect 168114 457538 168146 457774
rect 168382 457538 168466 457774
rect 168702 457538 168734 457774
rect 168114 457454 168734 457538
rect 168114 457218 168146 457454
rect 168382 457218 168466 457454
rect 168702 457218 168734 457454
rect 168114 423529 168734 457218
rect 171834 711558 172454 711590
rect 171834 711322 171866 711558
rect 172102 711322 172186 711558
rect 172422 711322 172454 711558
rect 171834 711238 172454 711322
rect 171834 711002 171866 711238
rect 172102 711002 172186 711238
rect 172422 711002 172454 711238
rect 171834 677494 172454 711002
rect 171834 677258 171866 677494
rect 172102 677258 172186 677494
rect 172422 677258 172454 677494
rect 171834 677174 172454 677258
rect 171834 676938 171866 677174
rect 172102 676938 172186 677174
rect 172422 676938 172454 677174
rect 171834 641494 172454 676938
rect 171834 641258 171866 641494
rect 172102 641258 172186 641494
rect 172422 641258 172454 641494
rect 171834 641174 172454 641258
rect 171834 640938 171866 641174
rect 172102 640938 172186 641174
rect 172422 640938 172454 641174
rect 171834 605494 172454 640938
rect 171834 605258 171866 605494
rect 172102 605258 172186 605494
rect 172422 605258 172454 605494
rect 171834 605174 172454 605258
rect 171834 604938 171866 605174
rect 172102 604938 172186 605174
rect 172422 604938 172454 605174
rect 171834 569494 172454 604938
rect 171834 569258 171866 569494
rect 172102 569258 172186 569494
rect 172422 569258 172454 569494
rect 171834 569174 172454 569258
rect 171834 568938 171866 569174
rect 172102 568938 172186 569174
rect 172422 568938 172454 569174
rect 171834 533494 172454 568938
rect 171834 533258 171866 533494
rect 172102 533258 172186 533494
rect 172422 533258 172454 533494
rect 171834 533174 172454 533258
rect 171834 532938 171866 533174
rect 172102 532938 172186 533174
rect 172422 532938 172454 533174
rect 171834 497494 172454 532938
rect 171834 497258 171866 497494
rect 172102 497258 172186 497494
rect 172422 497258 172454 497494
rect 171834 497174 172454 497258
rect 171834 496938 171866 497174
rect 172102 496938 172186 497174
rect 172422 496938 172454 497174
rect 171834 461494 172454 496938
rect 171834 461258 171866 461494
rect 172102 461258 172186 461494
rect 172422 461258 172454 461494
rect 171834 461174 172454 461258
rect 171834 460938 171866 461174
rect 172102 460938 172186 461174
rect 172422 460938 172454 461174
rect 171834 425494 172454 460938
rect 171834 425258 171866 425494
rect 172102 425258 172186 425494
rect 172422 425258 172454 425494
rect 171834 425174 172454 425258
rect 171834 424938 171866 425174
rect 172102 424938 172186 425174
rect 172422 424938 172454 425174
rect 171834 423529 172454 424938
rect 181794 704838 182414 711590
rect 181794 704602 181826 704838
rect 182062 704602 182146 704838
rect 182382 704602 182414 704838
rect 181794 704518 182414 704602
rect 181794 704282 181826 704518
rect 182062 704282 182146 704518
rect 182382 704282 182414 704518
rect 181794 687454 182414 704282
rect 181794 687218 181826 687454
rect 182062 687218 182146 687454
rect 182382 687218 182414 687454
rect 181794 687134 182414 687218
rect 181794 686898 181826 687134
rect 182062 686898 182146 687134
rect 182382 686898 182414 687134
rect 181794 651454 182414 686898
rect 181794 651218 181826 651454
rect 182062 651218 182146 651454
rect 182382 651218 182414 651454
rect 181794 651134 182414 651218
rect 181794 650898 181826 651134
rect 182062 650898 182146 651134
rect 182382 650898 182414 651134
rect 181794 615454 182414 650898
rect 181794 615218 181826 615454
rect 182062 615218 182146 615454
rect 182382 615218 182414 615454
rect 181794 615134 182414 615218
rect 181794 614898 181826 615134
rect 182062 614898 182146 615134
rect 182382 614898 182414 615134
rect 181794 579454 182414 614898
rect 181794 579218 181826 579454
rect 182062 579218 182146 579454
rect 182382 579218 182414 579454
rect 181794 579134 182414 579218
rect 181794 578898 181826 579134
rect 182062 578898 182146 579134
rect 182382 578898 182414 579134
rect 181794 543454 182414 578898
rect 181794 543218 181826 543454
rect 182062 543218 182146 543454
rect 182382 543218 182414 543454
rect 181794 543134 182414 543218
rect 181794 542898 181826 543134
rect 182062 542898 182146 543134
rect 182382 542898 182414 543134
rect 181794 507454 182414 542898
rect 181794 507218 181826 507454
rect 182062 507218 182146 507454
rect 182382 507218 182414 507454
rect 181794 507134 182414 507218
rect 181794 506898 181826 507134
rect 182062 506898 182146 507134
rect 182382 506898 182414 507134
rect 181794 471454 182414 506898
rect 181794 471218 181826 471454
rect 182062 471218 182146 471454
rect 182382 471218 182414 471454
rect 181794 471134 182414 471218
rect 181794 470898 181826 471134
rect 182062 470898 182146 471134
rect 182382 470898 182414 471134
rect 181794 435454 182414 470898
rect 181794 435218 181826 435454
rect 182062 435218 182146 435454
rect 182382 435218 182414 435454
rect 181794 435134 182414 435218
rect 181794 434898 181826 435134
rect 182062 434898 182146 435134
rect 182382 434898 182414 435134
rect 181794 423529 182414 434898
rect 185514 705798 186134 711590
rect 185514 705562 185546 705798
rect 185782 705562 185866 705798
rect 186102 705562 186134 705798
rect 185514 705478 186134 705562
rect 185514 705242 185546 705478
rect 185782 705242 185866 705478
rect 186102 705242 186134 705478
rect 185514 691174 186134 705242
rect 185514 690938 185546 691174
rect 185782 690938 185866 691174
rect 186102 690938 186134 691174
rect 185514 690854 186134 690938
rect 185514 690618 185546 690854
rect 185782 690618 185866 690854
rect 186102 690618 186134 690854
rect 185514 655174 186134 690618
rect 185514 654938 185546 655174
rect 185782 654938 185866 655174
rect 186102 654938 186134 655174
rect 185514 654854 186134 654938
rect 185514 654618 185546 654854
rect 185782 654618 185866 654854
rect 186102 654618 186134 654854
rect 185514 619174 186134 654618
rect 185514 618938 185546 619174
rect 185782 618938 185866 619174
rect 186102 618938 186134 619174
rect 185514 618854 186134 618938
rect 185514 618618 185546 618854
rect 185782 618618 185866 618854
rect 186102 618618 186134 618854
rect 185514 583174 186134 618618
rect 185514 582938 185546 583174
rect 185782 582938 185866 583174
rect 186102 582938 186134 583174
rect 185514 582854 186134 582938
rect 185514 582618 185546 582854
rect 185782 582618 185866 582854
rect 186102 582618 186134 582854
rect 185514 547174 186134 582618
rect 185514 546938 185546 547174
rect 185782 546938 185866 547174
rect 186102 546938 186134 547174
rect 185514 546854 186134 546938
rect 185514 546618 185546 546854
rect 185782 546618 185866 546854
rect 186102 546618 186134 546854
rect 185514 511174 186134 546618
rect 185514 510938 185546 511174
rect 185782 510938 185866 511174
rect 186102 510938 186134 511174
rect 185514 510854 186134 510938
rect 185514 510618 185546 510854
rect 185782 510618 185866 510854
rect 186102 510618 186134 510854
rect 185514 475174 186134 510618
rect 185514 474938 185546 475174
rect 185782 474938 185866 475174
rect 186102 474938 186134 475174
rect 185514 474854 186134 474938
rect 185514 474618 185546 474854
rect 185782 474618 185866 474854
rect 186102 474618 186134 474854
rect 185514 439174 186134 474618
rect 185514 438938 185546 439174
rect 185782 438938 185866 439174
rect 186102 438938 186134 439174
rect 185514 438854 186134 438938
rect 185514 438618 185546 438854
rect 185782 438618 185866 438854
rect 186102 438618 186134 438854
rect 185514 423529 186134 438618
rect 189234 706758 189854 711590
rect 189234 706522 189266 706758
rect 189502 706522 189586 706758
rect 189822 706522 189854 706758
rect 189234 706438 189854 706522
rect 189234 706202 189266 706438
rect 189502 706202 189586 706438
rect 189822 706202 189854 706438
rect 189234 694894 189854 706202
rect 189234 694658 189266 694894
rect 189502 694658 189586 694894
rect 189822 694658 189854 694894
rect 189234 694574 189854 694658
rect 189234 694338 189266 694574
rect 189502 694338 189586 694574
rect 189822 694338 189854 694574
rect 189234 658894 189854 694338
rect 189234 658658 189266 658894
rect 189502 658658 189586 658894
rect 189822 658658 189854 658894
rect 189234 658574 189854 658658
rect 189234 658338 189266 658574
rect 189502 658338 189586 658574
rect 189822 658338 189854 658574
rect 189234 622894 189854 658338
rect 189234 622658 189266 622894
rect 189502 622658 189586 622894
rect 189822 622658 189854 622894
rect 189234 622574 189854 622658
rect 189234 622338 189266 622574
rect 189502 622338 189586 622574
rect 189822 622338 189854 622574
rect 189234 586894 189854 622338
rect 189234 586658 189266 586894
rect 189502 586658 189586 586894
rect 189822 586658 189854 586894
rect 189234 586574 189854 586658
rect 189234 586338 189266 586574
rect 189502 586338 189586 586574
rect 189822 586338 189854 586574
rect 189234 550894 189854 586338
rect 189234 550658 189266 550894
rect 189502 550658 189586 550894
rect 189822 550658 189854 550894
rect 189234 550574 189854 550658
rect 189234 550338 189266 550574
rect 189502 550338 189586 550574
rect 189822 550338 189854 550574
rect 189234 514894 189854 550338
rect 189234 514658 189266 514894
rect 189502 514658 189586 514894
rect 189822 514658 189854 514894
rect 189234 514574 189854 514658
rect 189234 514338 189266 514574
rect 189502 514338 189586 514574
rect 189822 514338 189854 514574
rect 189234 478894 189854 514338
rect 189234 478658 189266 478894
rect 189502 478658 189586 478894
rect 189822 478658 189854 478894
rect 189234 478574 189854 478658
rect 189234 478338 189266 478574
rect 189502 478338 189586 478574
rect 189822 478338 189854 478574
rect 189234 442894 189854 478338
rect 189234 442658 189266 442894
rect 189502 442658 189586 442894
rect 189822 442658 189854 442894
rect 189234 442574 189854 442658
rect 189234 442338 189266 442574
rect 189502 442338 189586 442574
rect 189822 442338 189854 442574
rect 189234 423529 189854 442338
rect 192954 707718 193574 711590
rect 192954 707482 192986 707718
rect 193222 707482 193306 707718
rect 193542 707482 193574 707718
rect 192954 707398 193574 707482
rect 192954 707162 192986 707398
rect 193222 707162 193306 707398
rect 193542 707162 193574 707398
rect 192954 698614 193574 707162
rect 192954 698378 192986 698614
rect 193222 698378 193306 698614
rect 193542 698378 193574 698614
rect 192954 698294 193574 698378
rect 192954 698058 192986 698294
rect 193222 698058 193306 698294
rect 193542 698058 193574 698294
rect 192954 662614 193574 698058
rect 192954 662378 192986 662614
rect 193222 662378 193306 662614
rect 193542 662378 193574 662614
rect 192954 662294 193574 662378
rect 192954 662058 192986 662294
rect 193222 662058 193306 662294
rect 193542 662058 193574 662294
rect 192954 626614 193574 662058
rect 192954 626378 192986 626614
rect 193222 626378 193306 626614
rect 193542 626378 193574 626614
rect 192954 626294 193574 626378
rect 192954 626058 192986 626294
rect 193222 626058 193306 626294
rect 193542 626058 193574 626294
rect 192954 590614 193574 626058
rect 192954 590378 192986 590614
rect 193222 590378 193306 590614
rect 193542 590378 193574 590614
rect 192954 590294 193574 590378
rect 192954 590058 192986 590294
rect 193222 590058 193306 590294
rect 193542 590058 193574 590294
rect 192954 554614 193574 590058
rect 192954 554378 192986 554614
rect 193222 554378 193306 554614
rect 193542 554378 193574 554614
rect 192954 554294 193574 554378
rect 192954 554058 192986 554294
rect 193222 554058 193306 554294
rect 193542 554058 193574 554294
rect 192954 518614 193574 554058
rect 192954 518378 192986 518614
rect 193222 518378 193306 518614
rect 193542 518378 193574 518614
rect 192954 518294 193574 518378
rect 192954 518058 192986 518294
rect 193222 518058 193306 518294
rect 193542 518058 193574 518294
rect 192954 482614 193574 518058
rect 192954 482378 192986 482614
rect 193222 482378 193306 482614
rect 193542 482378 193574 482614
rect 192954 482294 193574 482378
rect 192954 482058 192986 482294
rect 193222 482058 193306 482294
rect 193542 482058 193574 482294
rect 192954 446614 193574 482058
rect 192954 446378 192986 446614
rect 193222 446378 193306 446614
rect 193542 446378 193574 446614
rect 192954 446294 193574 446378
rect 192954 446058 192986 446294
rect 193222 446058 193306 446294
rect 193542 446058 193574 446294
rect 192954 429868 193574 446058
rect 196674 708678 197294 711590
rect 196674 708442 196706 708678
rect 196942 708442 197026 708678
rect 197262 708442 197294 708678
rect 196674 708358 197294 708442
rect 196674 708122 196706 708358
rect 196942 708122 197026 708358
rect 197262 708122 197294 708358
rect 196674 666334 197294 708122
rect 196674 666098 196706 666334
rect 196942 666098 197026 666334
rect 197262 666098 197294 666334
rect 196674 666014 197294 666098
rect 196674 665778 196706 666014
rect 196942 665778 197026 666014
rect 197262 665778 197294 666014
rect 196674 630334 197294 665778
rect 196674 630098 196706 630334
rect 196942 630098 197026 630334
rect 197262 630098 197294 630334
rect 196674 630014 197294 630098
rect 196674 629778 196706 630014
rect 196942 629778 197026 630014
rect 197262 629778 197294 630014
rect 196674 594334 197294 629778
rect 196674 594098 196706 594334
rect 196942 594098 197026 594334
rect 197262 594098 197294 594334
rect 196674 594014 197294 594098
rect 196674 593778 196706 594014
rect 196942 593778 197026 594014
rect 197262 593778 197294 594014
rect 196674 558334 197294 593778
rect 196674 558098 196706 558334
rect 196942 558098 197026 558334
rect 197262 558098 197294 558334
rect 196674 558014 197294 558098
rect 196674 557778 196706 558014
rect 196942 557778 197026 558014
rect 197262 557778 197294 558014
rect 196674 522334 197294 557778
rect 196674 522098 196706 522334
rect 196942 522098 197026 522334
rect 197262 522098 197294 522334
rect 196674 522014 197294 522098
rect 196674 521778 196706 522014
rect 196942 521778 197026 522014
rect 197262 521778 197294 522014
rect 196674 486334 197294 521778
rect 196674 486098 196706 486334
rect 196942 486098 197026 486334
rect 197262 486098 197294 486334
rect 196674 486014 197294 486098
rect 196674 485778 196706 486014
rect 196942 485778 197026 486014
rect 197262 485778 197294 486014
rect 196674 450334 197294 485778
rect 196674 450098 196706 450334
rect 196942 450098 197026 450334
rect 197262 450098 197294 450334
rect 196674 450014 197294 450098
rect 196674 449778 196706 450014
rect 196942 449778 197026 450014
rect 197262 449778 197294 450014
rect 196674 423529 197294 449778
rect 200394 709638 201014 711590
rect 200394 709402 200426 709638
rect 200662 709402 200746 709638
rect 200982 709402 201014 709638
rect 200394 709318 201014 709402
rect 200394 709082 200426 709318
rect 200662 709082 200746 709318
rect 200982 709082 201014 709318
rect 200394 670054 201014 709082
rect 200394 669818 200426 670054
rect 200662 669818 200746 670054
rect 200982 669818 201014 670054
rect 200394 669734 201014 669818
rect 200394 669498 200426 669734
rect 200662 669498 200746 669734
rect 200982 669498 201014 669734
rect 200394 634054 201014 669498
rect 200394 633818 200426 634054
rect 200662 633818 200746 634054
rect 200982 633818 201014 634054
rect 200394 633734 201014 633818
rect 200394 633498 200426 633734
rect 200662 633498 200746 633734
rect 200982 633498 201014 633734
rect 200394 598054 201014 633498
rect 200394 597818 200426 598054
rect 200662 597818 200746 598054
rect 200982 597818 201014 598054
rect 200394 597734 201014 597818
rect 200394 597498 200426 597734
rect 200662 597498 200746 597734
rect 200982 597498 201014 597734
rect 200394 562054 201014 597498
rect 200394 561818 200426 562054
rect 200662 561818 200746 562054
rect 200982 561818 201014 562054
rect 200394 561734 201014 561818
rect 200394 561498 200426 561734
rect 200662 561498 200746 561734
rect 200982 561498 201014 561734
rect 200394 526054 201014 561498
rect 200394 525818 200426 526054
rect 200662 525818 200746 526054
rect 200982 525818 201014 526054
rect 200394 525734 201014 525818
rect 200394 525498 200426 525734
rect 200662 525498 200746 525734
rect 200982 525498 201014 525734
rect 200394 490054 201014 525498
rect 200394 489818 200426 490054
rect 200662 489818 200746 490054
rect 200982 489818 201014 490054
rect 200394 489734 201014 489818
rect 200394 489498 200426 489734
rect 200662 489498 200746 489734
rect 200982 489498 201014 489734
rect 200394 454054 201014 489498
rect 200394 453818 200426 454054
rect 200662 453818 200746 454054
rect 200982 453818 201014 454054
rect 200394 453734 201014 453818
rect 200394 453498 200426 453734
rect 200662 453498 200746 453734
rect 200982 453498 201014 453734
rect 200394 423529 201014 453498
rect 204114 710598 204734 711590
rect 204114 710362 204146 710598
rect 204382 710362 204466 710598
rect 204702 710362 204734 710598
rect 204114 710278 204734 710362
rect 204114 710042 204146 710278
rect 204382 710042 204466 710278
rect 204702 710042 204734 710278
rect 204114 673774 204734 710042
rect 204114 673538 204146 673774
rect 204382 673538 204466 673774
rect 204702 673538 204734 673774
rect 204114 673454 204734 673538
rect 204114 673218 204146 673454
rect 204382 673218 204466 673454
rect 204702 673218 204734 673454
rect 204114 637774 204734 673218
rect 204114 637538 204146 637774
rect 204382 637538 204466 637774
rect 204702 637538 204734 637774
rect 204114 637454 204734 637538
rect 204114 637218 204146 637454
rect 204382 637218 204466 637454
rect 204702 637218 204734 637454
rect 204114 601774 204734 637218
rect 204114 601538 204146 601774
rect 204382 601538 204466 601774
rect 204702 601538 204734 601774
rect 204114 601454 204734 601538
rect 204114 601218 204146 601454
rect 204382 601218 204466 601454
rect 204702 601218 204734 601454
rect 204114 565774 204734 601218
rect 204114 565538 204146 565774
rect 204382 565538 204466 565774
rect 204702 565538 204734 565774
rect 204114 565454 204734 565538
rect 204114 565218 204146 565454
rect 204382 565218 204466 565454
rect 204702 565218 204734 565454
rect 204114 529774 204734 565218
rect 204114 529538 204146 529774
rect 204382 529538 204466 529774
rect 204702 529538 204734 529774
rect 204114 529454 204734 529538
rect 204114 529218 204146 529454
rect 204382 529218 204466 529454
rect 204702 529218 204734 529454
rect 204114 493774 204734 529218
rect 204114 493538 204146 493774
rect 204382 493538 204466 493774
rect 204702 493538 204734 493774
rect 204114 493454 204734 493538
rect 204114 493218 204146 493454
rect 204382 493218 204466 493454
rect 204702 493218 204734 493454
rect 204114 457774 204734 493218
rect 204114 457538 204146 457774
rect 204382 457538 204466 457774
rect 204702 457538 204734 457774
rect 204114 457454 204734 457538
rect 204114 457218 204146 457454
rect 204382 457218 204466 457454
rect 204702 457218 204734 457454
rect 204114 423529 204734 457218
rect 207834 711558 208454 711590
rect 207834 711322 207866 711558
rect 208102 711322 208186 711558
rect 208422 711322 208454 711558
rect 207834 711238 208454 711322
rect 207834 711002 207866 711238
rect 208102 711002 208186 711238
rect 208422 711002 208454 711238
rect 207834 677494 208454 711002
rect 207834 677258 207866 677494
rect 208102 677258 208186 677494
rect 208422 677258 208454 677494
rect 207834 677174 208454 677258
rect 207834 676938 207866 677174
rect 208102 676938 208186 677174
rect 208422 676938 208454 677174
rect 207834 641494 208454 676938
rect 207834 641258 207866 641494
rect 208102 641258 208186 641494
rect 208422 641258 208454 641494
rect 207834 641174 208454 641258
rect 207834 640938 207866 641174
rect 208102 640938 208186 641174
rect 208422 640938 208454 641174
rect 207834 605494 208454 640938
rect 207834 605258 207866 605494
rect 208102 605258 208186 605494
rect 208422 605258 208454 605494
rect 207834 605174 208454 605258
rect 207834 604938 207866 605174
rect 208102 604938 208186 605174
rect 208422 604938 208454 605174
rect 207834 569494 208454 604938
rect 207834 569258 207866 569494
rect 208102 569258 208186 569494
rect 208422 569258 208454 569494
rect 207834 569174 208454 569258
rect 207834 568938 207866 569174
rect 208102 568938 208186 569174
rect 208422 568938 208454 569174
rect 207834 533494 208454 568938
rect 207834 533258 207866 533494
rect 208102 533258 208186 533494
rect 208422 533258 208454 533494
rect 207834 533174 208454 533258
rect 207834 532938 207866 533174
rect 208102 532938 208186 533174
rect 208422 532938 208454 533174
rect 207834 497494 208454 532938
rect 207834 497258 207866 497494
rect 208102 497258 208186 497494
rect 208422 497258 208454 497494
rect 207834 497174 208454 497258
rect 207834 496938 207866 497174
rect 208102 496938 208186 497174
rect 208422 496938 208454 497174
rect 207834 461494 208454 496938
rect 207834 461258 207866 461494
rect 208102 461258 208186 461494
rect 208422 461258 208454 461494
rect 207834 461174 208454 461258
rect 207834 460938 207866 461174
rect 208102 460938 208186 461174
rect 208422 460938 208454 461174
rect 207834 429868 208454 460938
rect 217794 704838 218414 711590
rect 217794 704602 217826 704838
rect 218062 704602 218146 704838
rect 218382 704602 218414 704838
rect 217794 704518 218414 704602
rect 217794 704282 217826 704518
rect 218062 704282 218146 704518
rect 218382 704282 218414 704518
rect 217794 687454 218414 704282
rect 217794 687218 217826 687454
rect 218062 687218 218146 687454
rect 218382 687218 218414 687454
rect 217794 687134 218414 687218
rect 217794 686898 217826 687134
rect 218062 686898 218146 687134
rect 218382 686898 218414 687134
rect 217794 651454 218414 686898
rect 217794 651218 217826 651454
rect 218062 651218 218146 651454
rect 218382 651218 218414 651454
rect 217794 651134 218414 651218
rect 217794 650898 217826 651134
rect 218062 650898 218146 651134
rect 218382 650898 218414 651134
rect 217794 615454 218414 650898
rect 217794 615218 217826 615454
rect 218062 615218 218146 615454
rect 218382 615218 218414 615454
rect 217794 615134 218414 615218
rect 217794 614898 217826 615134
rect 218062 614898 218146 615134
rect 218382 614898 218414 615134
rect 217794 579454 218414 614898
rect 217794 579218 217826 579454
rect 218062 579218 218146 579454
rect 218382 579218 218414 579454
rect 217794 579134 218414 579218
rect 217794 578898 217826 579134
rect 218062 578898 218146 579134
rect 218382 578898 218414 579134
rect 217794 543454 218414 578898
rect 217794 543218 217826 543454
rect 218062 543218 218146 543454
rect 218382 543218 218414 543454
rect 217794 543134 218414 543218
rect 217794 542898 217826 543134
rect 218062 542898 218146 543134
rect 218382 542898 218414 543134
rect 217794 507454 218414 542898
rect 217794 507218 217826 507454
rect 218062 507218 218146 507454
rect 218382 507218 218414 507454
rect 217794 507134 218414 507218
rect 217794 506898 217826 507134
rect 218062 506898 218146 507134
rect 218382 506898 218414 507134
rect 217794 471454 218414 506898
rect 217794 471218 217826 471454
rect 218062 471218 218146 471454
rect 218382 471218 218414 471454
rect 217794 471134 218414 471218
rect 217794 470898 217826 471134
rect 218062 470898 218146 471134
rect 218382 470898 218414 471134
rect 217794 435454 218414 470898
rect 217794 435218 217826 435454
rect 218062 435218 218146 435454
rect 218382 435218 218414 435454
rect 217794 435134 218414 435218
rect 217794 434898 217826 435134
rect 218062 434898 218146 435134
rect 218382 434898 218414 435134
rect 153234 406658 153266 406894
rect 153502 406658 153586 406894
rect 153822 406658 153854 406894
rect 153234 406574 153854 406658
rect 153234 406338 153266 406574
rect 153502 406338 153586 406574
rect 153822 406338 153854 406574
rect 153234 370894 153854 406338
rect 177568 403174 177888 403206
rect 177568 402938 177610 403174
rect 177846 402938 177888 403174
rect 177568 402854 177888 402938
rect 177568 402618 177610 402854
rect 177846 402618 177888 402854
rect 177568 402586 177888 402618
rect 208288 403174 208608 403206
rect 208288 402938 208330 403174
rect 208566 402938 208608 403174
rect 208288 402854 208608 402938
rect 208288 402618 208330 402854
rect 208566 402618 208608 402854
rect 208288 402586 208608 402618
rect 162208 399454 162528 399486
rect 162208 399218 162250 399454
rect 162486 399218 162528 399454
rect 162208 399134 162528 399218
rect 162208 398898 162250 399134
rect 162486 398898 162528 399134
rect 162208 398866 162528 398898
rect 192928 399454 193248 399486
rect 192928 399218 192970 399454
rect 193206 399218 193248 399454
rect 192928 399134 193248 399218
rect 192928 398898 192970 399134
rect 193206 398898 193248 399134
rect 192928 398866 193248 398898
rect 217794 399454 218414 434898
rect 217794 399218 217826 399454
rect 218062 399218 218146 399454
rect 218382 399218 218414 399454
rect 217794 399134 218414 399218
rect 217794 398898 217826 399134
rect 218062 398898 218146 399134
rect 218382 398898 218414 399134
rect 153234 370658 153266 370894
rect 153502 370658 153586 370894
rect 153822 370658 153854 370894
rect 153234 370574 153854 370658
rect 153234 370338 153266 370574
rect 153502 370338 153586 370574
rect 153822 370338 153854 370574
rect 153234 334894 153854 370338
rect 177568 367174 177888 367206
rect 177568 366938 177610 367174
rect 177846 366938 177888 367174
rect 177568 366854 177888 366938
rect 177568 366618 177610 366854
rect 177846 366618 177888 366854
rect 177568 366586 177888 366618
rect 208288 367174 208608 367206
rect 208288 366938 208330 367174
rect 208566 366938 208608 367174
rect 208288 366854 208608 366938
rect 208288 366618 208330 366854
rect 208566 366618 208608 366854
rect 208288 366586 208608 366618
rect 162208 363454 162528 363486
rect 162208 363218 162250 363454
rect 162486 363218 162528 363454
rect 162208 363134 162528 363218
rect 162208 362898 162250 363134
rect 162486 362898 162528 363134
rect 162208 362866 162528 362898
rect 192928 363454 193248 363486
rect 192928 363218 192970 363454
rect 193206 363218 193248 363454
rect 192928 363134 193248 363218
rect 192928 362898 192970 363134
rect 193206 362898 193248 363134
rect 192928 362866 193248 362898
rect 217794 363454 218414 398898
rect 217794 363218 217826 363454
rect 218062 363218 218146 363454
rect 218382 363218 218414 363454
rect 217794 363134 218414 363218
rect 217794 362898 217826 363134
rect 218062 362898 218146 363134
rect 218382 362898 218414 363134
rect 153234 334658 153266 334894
rect 153502 334658 153586 334894
rect 153822 334658 153854 334894
rect 153234 334574 153854 334658
rect 153234 334338 153266 334574
rect 153502 334338 153586 334574
rect 153822 334338 153854 334574
rect 153234 298894 153854 334338
rect 177568 331174 177888 331206
rect 177568 330938 177610 331174
rect 177846 330938 177888 331174
rect 177568 330854 177888 330938
rect 177568 330618 177610 330854
rect 177846 330618 177888 330854
rect 177568 330586 177888 330618
rect 208288 331174 208608 331206
rect 208288 330938 208330 331174
rect 208566 330938 208608 331174
rect 208288 330854 208608 330938
rect 208288 330618 208330 330854
rect 208566 330618 208608 330854
rect 208288 330586 208608 330618
rect 162208 327454 162528 327486
rect 162208 327218 162250 327454
rect 162486 327218 162528 327454
rect 162208 327134 162528 327218
rect 162208 326898 162250 327134
rect 162486 326898 162528 327134
rect 162208 326866 162528 326898
rect 192928 327454 193248 327486
rect 192928 327218 192970 327454
rect 193206 327218 193248 327454
rect 192928 327134 193248 327218
rect 192928 326898 192970 327134
rect 193206 326898 193248 327134
rect 192928 326866 193248 326898
rect 217794 327454 218414 362898
rect 217794 327218 217826 327454
rect 218062 327218 218146 327454
rect 218382 327218 218414 327454
rect 217794 327134 218414 327218
rect 217794 326898 217826 327134
rect 218062 326898 218146 327134
rect 218382 326898 218414 327134
rect 153234 298658 153266 298894
rect 153502 298658 153586 298894
rect 153822 298658 153854 298894
rect 153234 298574 153854 298658
rect 153234 298338 153266 298574
rect 153502 298338 153586 298574
rect 153822 298338 153854 298574
rect 153234 262894 153854 298338
rect 177568 295174 177888 295206
rect 177568 294938 177610 295174
rect 177846 294938 177888 295174
rect 177568 294854 177888 294938
rect 177568 294618 177610 294854
rect 177846 294618 177888 294854
rect 177568 294586 177888 294618
rect 208288 295174 208608 295206
rect 208288 294938 208330 295174
rect 208566 294938 208608 295174
rect 208288 294854 208608 294938
rect 208288 294618 208330 294854
rect 208566 294618 208608 294854
rect 208288 294586 208608 294618
rect 155355 293180 155421 293181
rect 155355 293116 155356 293180
rect 155420 293116 155421 293180
rect 155355 293115 155421 293116
rect 153234 262658 153266 262894
rect 153502 262658 153586 262894
rect 153822 262658 153854 262894
rect 153234 262574 153854 262658
rect 153234 262338 153266 262574
rect 153502 262338 153586 262574
rect 153822 262338 153854 262574
rect 153234 226894 153854 262338
rect 153234 226658 153266 226894
rect 153502 226658 153586 226894
rect 153822 226658 153854 226894
rect 153234 226574 153854 226658
rect 153234 226338 153266 226574
rect 153502 226338 153586 226574
rect 153822 226338 153854 226574
rect 153234 190894 153854 226338
rect 153234 190658 153266 190894
rect 153502 190658 153586 190894
rect 153822 190658 153854 190894
rect 153234 190574 153854 190658
rect 153234 190338 153266 190574
rect 153502 190338 153586 190574
rect 153822 190338 153854 190574
rect 153234 154894 153854 190338
rect 155358 171189 155418 293115
rect 162208 291454 162528 291486
rect 162208 291218 162250 291454
rect 162486 291218 162528 291454
rect 162208 291134 162528 291218
rect 162208 290898 162250 291134
rect 162486 290898 162528 291134
rect 162208 290866 162528 290898
rect 192928 291454 193248 291486
rect 192928 291218 192970 291454
rect 193206 291218 193248 291454
rect 192928 291134 193248 291218
rect 192928 290898 192970 291134
rect 193206 290898 193248 291134
rect 192928 290866 193248 290898
rect 217794 291454 218414 326898
rect 217794 291218 217826 291454
rect 218062 291218 218146 291454
rect 218382 291218 218414 291454
rect 217794 291134 218414 291218
rect 217794 290898 217826 291134
rect 218062 290898 218146 291134
rect 218382 290898 218414 291134
rect 156954 266614 157574 270287
rect 156954 266378 156986 266614
rect 157222 266378 157306 266614
rect 157542 266378 157574 266614
rect 156954 266294 157574 266378
rect 156954 266058 156986 266294
rect 157222 266058 157306 266294
rect 157542 266058 157574 266294
rect 156954 230614 157574 266058
rect 156954 230378 156986 230614
rect 157222 230378 157306 230614
rect 157542 230378 157574 230614
rect 156954 230294 157574 230378
rect 156954 230058 156986 230294
rect 157222 230058 157306 230294
rect 157542 230058 157574 230294
rect 156954 194614 157574 230058
rect 156954 194378 156986 194614
rect 157222 194378 157306 194614
rect 157542 194378 157574 194614
rect 156954 194294 157574 194378
rect 156954 194058 156986 194294
rect 157222 194058 157306 194294
rect 157542 194058 157574 194294
rect 155355 171188 155421 171189
rect 155355 171124 155356 171188
rect 155420 171124 155421 171188
rect 155355 171123 155421 171124
rect 153234 154658 153266 154894
rect 153502 154658 153586 154894
rect 153822 154658 153854 154894
rect 153234 154574 153854 154658
rect 153234 154338 153266 154574
rect 153502 154338 153586 154574
rect 153822 154338 153854 154574
rect 153234 118894 153854 154338
rect 153234 118658 153266 118894
rect 153502 118658 153586 118894
rect 153822 118658 153854 118894
rect 153234 118574 153854 118658
rect 153234 118338 153266 118574
rect 153502 118338 153586 118574
rect 153822 118338 153854 118574
rect 153234 82894 153854 118338
rect 153234 82658 153266 82894
rect 153502 82658 153586 82894
rect 153822 82658 153854 82894
rect 153234 82574 153854 82658
rect 153234 82338 153266 82574
rect 153502 82338 153586 82574
rect 153822 82338 153854 82574
rect 153234 46894 153854 82338
rect 153234 46658 153266 46894
rect 153502 46658 153586 46894
rect 153822 46658 153854 46894
rect 153234 46574 153854 46658
rect 153234 46338 153266 46574
rect 153502 46338 153586 46574
rect 153822 46338 153854 46574
rect 153234 10894 153854 46338
rect 153234 10658 153266 10894
rect 153502 10658 153586 10894
rect 153822 10658 153854 10894
rect 153234 10574 153854 10658
rect 153234 10338 153266 10574
rect 153502 10338 153586 10574
rect 153822 10338 153854 10574
rect 153234 -2266 153854 10338
rect 153234 -2502 153266 -2266
rect 153502 -2502 153586 -2266
rect 153822 -2502 153854 -2266
rect 153234 -2586 153854 -2502
rect 153234 -2822 153266 -2586
rect 153502 -2822 153586 -2586
rect 153822 -2822 153854 -2586
rect 153234 -7654 153854 -2822
rect 156954 158614 157574 194058
rect 156954 158378 156986 158614
rect 157222 158378 157306 158614
rect 157542 158378 157574 158614
rect 156954 158294 157574 158378
rect 156954 158058 156986 158294
rect 157222 158058 157306 158294
rect 157542 158058 157574 158294
rect 156954 122614 157574 158058
rect 160674 234334 161294 270287
rect 160674 234098 160706 234334
rect 160942 234098 161026 234334
rect 161262 234098 161294 234334
rect 160674 234014 161294 234098
rect 160674 233778 160706 234014
rect 160942 233778 161026 234014
rect 161262 233778 161294 234014
rect 160674 198334 161294 233778
rect 160674 198098 160706 198334
rect 160942 198098 161026 198334
rect 161262 198098 161294 198334
rect 160674 198014 161294 198098
rect 160674 197778 160706 198014
rect 160942 197778 161026 198014
rect 161262 197778 161294 198014
rect 160674 162334 161294 197778
rect 160674 162098 160706 162334
rect 160942 162098 161026 162334
rect 161262 162098 161294 162334
rect 160674 162014 161294 162098
rect 160674 161778 160706 162014
rect 160942 161778 161026 162014
rect 161262 161778 161294 162014
rect 160674 131409 161294 161778
rect 164394 238054 165014 270287
rect 164394 237818 164426 238054
rect 164662 237818 164746 238054
rect 164982 237818 165014 238054
rect 164394 237734 165014 237818
rect 164394 237498 164426 237734
rect 164662 237498 164746 237734
rect 164982 237498 165014 237734
rect 164394 202054 165014 237498
rect 164394 201818 164426 202054
rect 164662 201818 164746 202054
rect 164982 201818 165014 202054
rect 164394 201734 165014 201818
rect 164394 201498 164426 201734
rect 164662 201498 164746 201734
rect 164982 201498 165014 201734
rect 164394 166054 165014 201498
rect 164394 165818 164426 166054
rect 164662 165818 164746 166054
rect 164982 165818 165014 166054
rect 164394 165734 165014 165818
rect 164394 165498 164426 165734
rect 164662 165498 164746 165734
rect 164982 165498 165014 165734
rect 164394 131409 165014 165498
rect 168114 241774 168734 270287
rect 168114 241538 168146 241774
rect 168382 241538 168466 241774
rect 168702 241538 168734 241774
rect 168114 241454 168734 241538
rect 168114 241218 168146 241454
rect 168382 241218 168466 241454
rect 168702 241218 168734 241454
rect 168114 205774 168734 241218
rect 168114 205538 168146 205774
rect 168382 205538 168466 205774
rect 168702 205538 168734 205774
rect 168114 205454 168734 205538
rect 168114 205218 168146 205454
rect 168382 205218 168466 205454
rect 168702 205218 168734 205454
rect 168114 169774 168734 205218
rect 168114 169538 168146 169774
rect 168382 169538 168466 169774
rect 168702 169538 168734 169774
rect 168114 169454 168734 169538
rect 168114 169218 168146 169454
rect 168382 169218 168466 169454
rect 168702 169218 168734 169454
rect 168114 133774 168734 169218
rect 168114 133538 168146 133774
rect 168382 133538 168466 133774
rect 168702 133538 168734 133774
rect 168114 133454 168734 133538
rect 168114 133218 168146 133454
rect 168382 133218 168466 133454
rect 168702 133218 168734 133454
rect 168114 131409 168734 133218
rect 171834 245494 172454 270287
rect 171834 245258 171866 245494
rect 172102 245258 172186 245494
rect 172422 245258 172454 245494
rect 171834 245174 172454 245258
rect 171834 244938 171866 245174
rect 172102 244938 172186 245174
rect 172422 244938 172454 245174
rect 171834 209494 172454 244938
rect 171834 209258 171866 209494
rect 172102 209258 172186 209494
rect 172422 209258 172454 209494
rect 171834 209174 172454 209258
rect 171834 208938 171866 209174
rect 172102 208938 172186 209174
rect 172422 208938 172454 209174
rect 171834 173494 172454 208938
rect 171834 173258 171866 173494
rect 172102 173258 172186 173494
rect 172422 173258 172454 173494
rect 171834 173174 172454 173258
rect 171834 172938 171866 173174
rect 172102 172938 172186 173174
rect 172422 172938 172454 173174
rect 171834 137494 172454 172938
rect 171834 137258 171866 137494
rect 172102 137258 172186 137494
rect 172422 137258 172454 137494
rect 171834 137174 172454 137258
rect 171834 136938 171866 137174
rect 172102 136938 172186 137174
rect 172422 136938 172454 137174
rect 171834 131409 172454 136938
rect 181794 255454 182414 270287
rect 181794 255218 181826 255454
rect 182062 255218 182146 255454
rect 182382 255218 182414 255454
rect 181794 255134 182414 255218
rect 181794 254898 181826 255134
rect 182062 254898 182146 255134
rect 182382 254898 182414 255134
rect 181794 219454 182414 254898
rect 181794 219218 181826 219454
rect 182062 219218 182146 219454
rect 182382 219218 182414 219454
rect 181794 219134 182414 219218
rect 181794 218898 181826 219134
rect 182062 218898 182146 219134
rect 182382 218898 182414 219134
rect 181794 183454 182414 218898
rect 181794 183218 181826 183454
rect 182062 183218 182146 183454
rect 182382 183218 182414 183454
rect 181794 183134 182414 183218
rect 181794 182898 181826 183134
rect 182062 182898 182146 183134
rect 182382 182898 182414 183134
rect 181794 147454 182414 182898
rect 181794 147218 181826 147454
rect 182062 147218 182146 147454
rect 182382 147218 182414 147454
rect 181794 147134 182414 147218
rect 181794 146898 181826 147134
rect 182062 146898 182146 147134
rect 182382 146898 182414 147134
rect 181794 131409 182414 146898
rect 185514 259174 186134 270287
rect 185514 258938 185546 259174
rect 185782 258938 185866 259174
rect 186102 258938 186134 259174
rect 185514 258854 186134 258938
rect 185514 258618 185546 258854
rect 185782 258618 185866 258854
rect 186102 258618 186134 258854
rect 185514 223174 186134 258618
rect 185514 222938 185546 223174
rect 185782 222938 185866 223174
rect 186102 222938 186134 223174
rect 185514 222854 186134 222938
rect 185514 222618 185546 222854
rect 185782 222618 185866 222854
rect 186102 222618 186134 222854
rect 185514 187174 186134 222618
rect 185514 186938 185546 187174
rect 185782 186938 185866 187174
rect 186102 186938 186134 187174
rect 185514 186854 186134 186938
rect 185514 186618 185546 186854
rect 185782 186618 185866 186854
rect 186102 186618 186134 186854
rect 185514 151174 186134 186618
rect 185514 150938 185546 151174
rect 185782 150938 185866 151174
rect 186102 150938 186134 151174
rect 185514 150854 186134 150938
rect 185514 150618 185546 150854
rect 185782 150618 185866 150854
rect 186102 150618 186134 150854
rect 185514 131409 186134 150618
rect 189234 262894 189854 270287
rect 189234 262658 189266 262894
rect 189502 262658 189586 262894
rect 189822 262658 189854 262894
rect 189234 262574 189854 262658
rect 189234 262338 189266 262574
rect 189502 262338 189586 262574
rect 189822 262338 189854 262574
rect 189234 226894 189854 262338
rect 189234 226658 189266 226894
rect 189502 226658 189586 226894
rect 189822 226658 189854 226894
rect 189234 226574 189854 226658
rect 189234 226338 189266 226574
rect 189502 226338 189586 226574
rect 189822 226338 189854 226574
rect 189234 190894 189854 226338
rect 189234 190658 189266 190894
rect 189502 190658 189586 190894
rect 189822 190658 189854 190894
rect 189234 190574 189854 190658
rect 189234 190338 189266 190574
rect 189502 190338 189586 190574
rect 189822 190338 189854 190574
rect 189234 154894 189854 190338
rect 189234 154658 189266 154894
rect 189502 154658 189586 154894
rect 189822 154658 189854 154894
rect 189234 154574 189854 154658
rect 189234 154338 189266 154574
rect 189502 154338 189586 154574
rect 189822 154338 189854 154574
rect 189234 131409 189854 154338
rect 192954 266614 193574 270068
rect 192954 266378 192986 266614
rect 193222 266378 193306 266614
rect 193542 266378 193574 266614
rect 192954 266294 193574 266378
rect 192954 266058 192986 266294
rect 193222 266058 193306 266294
rect 193542 266058 193574 266294
rect 192954 230614 193574 266058
rect 192954 230378 192986 230614
rect 193222 230378 193306 230614
rect 193542 230378 193574 230614
rect 192954 230294 193574 230378
rect 192954 230058 192986 230294
rect 193222 230058 193306 230294
rect 193542 230058 193574 230294
rect 192954 194614 193574 230058
rect 192954 194378 192986 194614
rect 193222 194378 193306 194614
rect 193542 194378 193574 194614
rect 192954 194294 193574 194378
rect 192954 194058 192986 194294
rect 193222 194058 193306 194294
rect 193542 194058 193574 194294
rect 192954 158614 193574 194058
rect 192954 158378 192986 158614
rect 193222 158378 193306 158614
rect 193542 158378 193574 158614
rect 192954 158294 193574 158378
rect 192954 158058 192986 158294
rect 193222 158058 193306 158294
rect 193542 158058 193574 158294
rect 192954 131900 193574 158058
rect 196674 234334 197294 270287
rect 196674 234098 196706 234334
rect 196942 234098 197026 234334
rect 197262 234098 197294 234334
rect 196674 234014 197294 234098
rect 196674 233778 196706 234014
rect 196942 233778 197026 234014
rect 197262 233778 197294 234014
rect 196674 198334 197294 233778
rect 196674 198098 196706 198334
rect 196942 198098 197026 198334
rect 197262 198098 197294 198334
rect 196674 198014 197294 198098
rect 196674 197778 196706 198014
rect 196942 197778 197026 198014
rect 197262 197778 197294 198014
rect 196674 162334 197294 197778
rect 196674 162098 196706 162334
rect 196942 162098 197026 162334
rect 197262 162098 197294 162334
rect 196674 162014 197294 162098
rect 196674 161778 196706 162014
rect 196942 161778 197026 162014
rect 197262 161778 197294 162014
rect 156954 122378 156986 122614
rect 157222 122378 157306 122614
rect 157542 122378 157574 122614
rect 156954 122294 157574 122378
rect 156954 122058 156986 122294
rect 157222 122058 157306 122294
rect 157542 122058 157574 122294
rect 156954 86614 157574 122058
rect 196674 126334 197294 161778
rect 196674 126098 196706 126334
rect 196942 126098 197026 126334
rect 197262 126098 197294 126334
rect 196674 126014 197294 126098
rect 196674 125778 196706 126014
rect 196942 125778 197026 126014
rect 197262 125778 197294 126014
rect 177568 115174 177888 115206
rect 177568 114938 177610 115174
rect 177846 114938 177888 115174
rect 177568 114854 177888 114938
rect 177568 114618 177610 114854
rect 177846 114618 177888 114854
rect 177568 114586 177888 114618
rect 162208 111454 162528 111486
rect 162208 111218 162250 111454
rect 162486 111218 162528 111454
rect 162208 111134 162528 111218
rect 162208 110898 162250 111134
rect 162486 110898 162528 111134
rect 162208 110866 162528 110898
rect 192928 111454 193248 111486
rect 192928 111218 192970 111454
rect 193206 111218 193248 111454
rect 192928 111134 193248 111218
rect 192928 110898 192970 111134
rect 193206 110898 193248 111134
rect 192928 110866 193248 110898
rect 156954 86378 156986 86614
rect 157222 86378 157306 86614
rect 157542 86378 157574 86614
rect 156954 86294 157574 86378
rect 156954 86058 156986 86294
rect 157222 86058 157306 86294
rect 157542 86058 157574 86294
rect 156954 50614 157574 86058
rect 196674 90334 197294 125778
rect 196674 90098 196706 90334
rect 196942 90098 197026 90334
rect 197262 90098 197294 90334
rect 196674 90014 197294 90098
rect 196674 89778 196706 90014
rect 196942 89778 197026 90014
rect 197262 89778 197294 90014
rect 177568 79174 177888 79206
rect 177568 78938 177610 79174
rect 177846 78938 177888 79174
rect 177568 78854 177888 78938
rect 177568 78618 177610 78854
rect 177846 78618 177888 78854
rect 177568 78586 177888 78618
rect 162208 75454 162528 75486
rect 162208 75218 162250 75454
rect 162486 75218 162528 75454
rect 162208 75134 162528 75218
rect 162208 74898 162250 75134
rect 162486 74898 162528 75134
rect 162208 74866 162528 74898
rect 192928 75454 193248 75486
rect 192928 75218 192970 75454
rect 193206 75218 193248 75454
rect 192928 75134 193248 75218
rect 192928 74898 192970 75134
rect 193206 74898 193248 75134
rect 192928 74866 193248 74898
rect 196674 54334 197294 89778
rect 196674 54098 196706 54334
rect 196942 54098 197026 54334
rect 197262 54098 197294 54334
rect 196674 54014 197294 54098
rect 196674 53778 196706 54014
rect 196942 53778 197026 54014
rect 197262 53778 197294 54014
rect 173571 52732 173637 52733
rect 173571 52668 173572 52732
rect 173636 52668 173637 52732
rect 173571 52667 173637 52668
rect 169891 52324 169957 52325
rect 169891 52260 169892 52324
rect 169956 52260 169957 52324
rect 169891 52259 169957 52260
rect 161795 52052 161861 52053
rect 161795 51988 161796 52052
rect 161860 51988 161861 52052
rect 161795 51987 161861 51988
rect 163635 52052 163701 52053
rect 163635 51988 163636 52052
rect 163700 51988 163701 52052
rect 163635 51987 163701 51988
rect 169155 52052 169221 52053
rect 169155 51988 169156 52052
rect 169220 51988 169221 52052
rect 169155 51987 169221 51988
rect 160323 51916 160389 51917
rect 160323 51852 160324 51916
rect 160388 51852 160389 51916
rect 160323 51851 160389 51852
rect 161427 51916 161493 51917
rect 161427 51852 161428 51916
rect 161492 51852 161493 51916
rect 161427 51851 161493 51852
rect 160139 51780 160205 51781
rect 160139 51716 160140 51780
rect 160204 51716 160205 51780
rect 160139 51715 160205 51716
rect 156954 50378 156986 50614
rect 157222 50378 157306 50614
rect 157542 50378 157574 50614
rect 156954 50294 157574 50378
rect 156954 50058 156986 50294
rect 157222 50058 157306 50294
rect 157542 50058 157574 50294
rect 156954 14614 157574 50058
rect 156954 14378 156986 14614
rect 157222 14378 157306 14614
rect 157542 14378 157574 14614
rect 156954 14294 157574 14378
rect 156954 14058 156986 14294
rect 157222 14058 157306 14294
rect 157542 14058 157574 14294
rect 156954 -3226 157574 14058
rect 160142 11661 160202 51715
rect 160326 21317 160386 51851
rect 160323 21316 160389 21317
rect 160323 21252 160324 21316
rect 160388 21252 160389 21316
rect 160323 21251 160389 21252
rect 160674 18334 161294 50791
rect 161430 46069 161490 51851
rect 161611 51644 161677 51645
rect 161611 51580 161612 51644
rect 161676 51580 161677 51644
rect 161611 51579 161677 51580
rect 161427 46068 161493 46069
rect 161427 46004 161428 46068
rect 161492 46004 161493 46068
rect 161427 46003 161493 46004
rect 160674 18098 160706 18334
rect 160942 18098 161026 18334
rect 161262 18098 161294 18334
rect 160674 18014 161294 18098
rect 160674 17778 160706 18014
rect 160942 17778 161026 18014
rect 161262 17778 161294 18014
rect 160139 11660 160205 11661
rect 160139 11596 160140 11660
rect 160204 11596 160205 11660
rect 160139 11595 160205 11596
rect 156954 -3462 156986 -3226
rect 157222 -3462 157306 -3226
rect 157542 -3462 157574 -3226
rect 156954 -3546 157574 -3462
rect 156954 -3782 156986 -3546
rect 157222 -3782 157306 -3546
rect 157542 -3782 157574 -3546
rect 156954 -7654 157574 -3782
rect 160674 -4186 161294 17778
rect 161614 8941 161674 51579
rect 161798 18597 161858 51987
rect 162163 51916 162229 51917
rect 162163 51852 162164 51916
rect 162228 51852 162229 51916
rect 162163 51851 162229 51852
rect 162715 51916 162781 51917
rect 162715 51852 162716 51916
rect 162780 51852 162781 51916
rect 162715 51851 162781 51852
rect 161979 48924 162045 48925
rect 161979 48860 161980 48924
rect 162044 48860 162045 48924
rect 161979 48859 162045 48860
rect 161982 22677 162042 48859
rect 162166 46341 162226 51851
rect 162163 46340 162229 46341
rect 162163 46276 162164 46340
rect 162228 46276 162229 46340
rect 162163 46275 162229 46276
rect 162718 45933 162778 51851
rect 162899 51780 162965 51781
rect 162899 51716 162900 51780
rect 162964 51716 162965 51780
rect 162899 51715 162965 51716
rect 162715 45932 162781 45933
rect 162715 45868 162716 45932
rect 162780 45868 162781 45932
rect 162715 45867 162781 45868
rect 161979 22676 162045 22677
rect 161979 22612 161980 22676
rect 162044 22612 162045 22676
rect 161979 22611 162045 22612
rect 161795 18596 161861 18597
rect 161795 18532 161796 18596
rect 161860 18532 161861 18596
rect 161795 18531 161861 18532
rect 161611 8940 161677 8941
rect 161611 8876 161612 8940
rect 161676 8876 161677 8940
rect 161611 8875 161677 8876
rect 162902 6221 162962 51715
rect 163267 48924 163333 48925
rect 163267 48860 163268 48924
rect 163332 48860 163333 48924
rect 163267 48859 163333 48860
rect 163083 48788 163149 48789
rect 163083 48724 163084 48788
rect 163148 48724 163149 48788
rect 163083 48723 163149 48724
rect 163086 6357 163146 48723
rect 163270 10301 163330 48859
rect 163451 48788 163517 48789
rect 163451 48724 163452 48788
rect 163516 48724 163517 48788
rect 163451 48723 163517 48724
rect 163454 15877 163514 48723
rect 163638 46885 163698 51987
rect 165843 51916 165909 51917
rect 165843 51852 165844 51916
rect 165908 51852 165909 51916
rect 165843 51851 165909 51852
rect 167499 51916 167565 51917
rect 167499 51852 167500 51916
rect 167564 51852 167565 51916
rect 167499 51851 167565 51852
rect 163819 51508 163885 51509
rect 163819 51444 163820 51508
rect 163884 51444 163885 51508
rect 163819 51443 163885 51444
rect 163822 47565 163882 51443
rect 163819 47564 163885 47565
rect 163819 47500 163820 47564
rect 163884 47500 163885 47564
rect 163819 47499 163885 47500
rect 163635 46884 163701 46885
rect 163635 46820 163636 46884
rect 163700 46820 163701 46884
rect 163635 46819 163701 46820
rect 164394 22054 165014 50791
rect 165659 49468 165725 49469
rect 165659 49404 165660 49468
rect 165724 49404 165725 49468
rect 165659 49403 165725 49404
rect 165291 48652 165357 48653
rect 165291 48588 165292 48652
rect 165356 48588 165357 48652
rect 165291 48587 165357 48588
rect 164394 21818 164426 22054
rect 164662 21818 164746 22054
rect 164982 21818 165014 22054
rect 164394 21734 165014 21818
rect 164394 21498 164426 21734
rect 164662 21498 164746 21734
rect 164982 21498 165014 21734
rect 163451 15876 163517 15877
rect 163451 15812 163452 15876
rect 163516 15812 163517 15876
rect 163451 15811 163517 15812
rect 163267 10300 163333 10301
rect 163267 10236 163268 10300
rect 163332 10236 163333 10300
rect 163267 10235 163333 10236
rect 163083 6356 163149 6357
rect 163083 6292 163084 6356
rect 163148 6292 163149 6356
rect 163083 6291 163149 6292
rect 162899 6220 162965 6221
rect 162899 6156 162900 6220
rect 162964 6156 162965 6220
rect 162899 6155 162965 6156
rect 160674 -4422 160706 -4186
rect 160942 -4422 161026 -4186
rect 161262 -4422 161294 -4186
rect 160674 -4506 161294 -4422
rect 160674 -4742 160706 -4506
rect 160942 -4742 161026 -4506
rect 161262 -4742 161294 -4506
rect 160674 -7654 161294 -4742
rect 164394 -5146 165014 21498
rect 165294 4861 165354 48587
rect 165662 4997 165722 49403
rect 165846 13021 165906 51851
rect 166027 51780 166093 51781
rect 166027 51716 166028 51780
rect 166092 51716 166093 51780
rect 166027 51715 166093 51716
rect 166763 51780 166829 51781
rect 166763 51716 166764 51780
rect 166828 51716 166829 51780
rect 166763 51715 166829 51716
rect 166030 14517 166090 51715
rect 166211 49468 166277 49469
rect 166211 49404 166212 49468
rect 166276 49404 166277 49468
rect 166211 49403 166277 49404
rect 166214 17237 166274 49403
rect 166766 47429 166826 51715
rect 167315 47564 167381 47565
rect 167315 47500 167316 47564
rect 167380 47500 167381 47564
rect 167315 47499 167381 47500
rect 166763 47428 166829 47429
rect 166763 47364 166764 47428
rect 166828 47364 166829 47428
rect 166763 47363 166829 47364
rect 167131 47428 167197 47429
rect 167131 47364 167132 47428
rect 167196 47364 167197 47428
rect 167131 47363 167197 47364
rect 166947 41444 167013 41445
rect 166947 41380 166948 41444
rect 167012 41380 167013 41444
rect 166947 41379 167013 41380
rect 166211 17236 166277 17237
rect 166211 17172 166212 17236
rect 166276 17172 166277 17236
rect 166211 17171 166277 17172
rect 166027 14516 166093 14517
rect 166027 14452 166028 14516
rect 166092 14452 166093 14516
rect 166027 14451 166093 14452
rect 166950 13157 167010 41379
rect 167134 14653 167194 47363
rect 167318 21453 167378 47499
rect 167502 45797 167562 51851
rect 168971 51508 169037 51509
rect 168971 51444 168972 51508
rect 169036 51444 169037 51508
rect 168971 51443 169037 51444
rect 167683 47700 167749 47701
rect 167683 47636 167684 47700
rect 167748 47636 167749 47700
rect 167683 47635 167749 47636
rect 167499 45796 167565 45797
rect 167499 45732 167500 45796
rect 167564 45732 167565 45796
rect 167499 45731 167565 45732
rect 167686 41445 167746 47635
rect 167683 41444 167749 41445
rect 167683 41380 167684 41444
rect 167748 41380 167749 41444
rect 167683 41379 167749 41380
rect 168114 25774 168734 50791
rect 168114 25538 168146 25774
rect 168382 25538 168466 25774
rect 168702 25538 168734 25774
rect 168114 25454 168734 25538
rect 168114 25218 168146 25454
rect 168382 25218 168466 25454
rect 168702 25218 168734 25454
rect 167315 21452 167381 21453
rect 167315 21388 167316 21452
rect 167380 21388 167381 21452
rect 167315 21387 167381 21388
rect 167131 14652 167197 14653
rect 167131 14588 167132 14652
rect 167196 14588 167197 14652
rect 167131 14587 167197 14588
rect 166947 13156 167013 13157
rect 166947 13092 166948 13156
rect 167012 13092 167013 13156
rect 166947 13091 167013 13092
rect 165843 13020 165909 13021
rect 165843 12956 165844 13020
rect 165908 12956 165909 13020
rect 165843 12955 165909 12956
rect 165659 4996 165725 4997
rect 165659 4932 165660 4996
rect 165724 4932 165725 4996
rect 165659 4931 165725 4932
rect 165291 4860 165357 4861
rect 165291 4796 165292 4860
rect 165356 4796 165357 4860
rect 165291 4795 165357 4796
rect 164394 -5382 164426 -5146
rect 164662 -5382 164746 -5146
rect 164982 -5382 165014 -5146
rect 164394 -5466 165014 -5382
rect 164394 -5702 164426 -5466
rect 164662 -5702 164746 -5466
rect 164982 -5702 165014 -5466
rect 164394 -7654 165014 -5702
rect 168114 -6106 168734 25218
rect 168974 5133 169034 51443
rect 169158 9213 169218 51987
rect 169707 51916 169773 51917
rect 169707 51852 169708 51916
rect 169772 51852 169773 51916
rect 169707 51851 169773 51852
rect 169710 50285 169770 51851
rect 169894 51509 169954 52259
rect 170443 51916 170509 51917
rect 170443 51852 170444 51916
rect 170508 51852 170509 51916
rect 170443 51851 170509 51852
rect 173387 51916 173453 51917
rect 173387 51852 173388 51916
rect 173452 51852 173453 51916
rect 173387 51851 173453 51852
rect 170075 51780 170141 51781
rect 170075 51716 170076 51780
rect 170140 51716 170141 51780
rect 170075 51715 170141 51716
rect 169891 51508 169957 51509
rect 169891 51444 169892 51508
rect 169956 51444 169957 51508
rect 169891 51443 169957 51444
rect 169707 50284 169773 50285
rect 169707 50220 169708 50284
rect 169772 50220 169773 50284
rect 169707 50219 169773 50220
rect 170078 48925 170138 51715
rect 170075 48924 170141 48925
rect 170075 48860 170076 48924
rect 170140 48860 170141 48924
rect 170075 48859 170141 48860
rect 170446 48653 170506 51851
rect 173019 51780 173085 51781
rect 173019 51716 173020 51780
rect 173084 51716 173085 51780
rect 173019 51715 173085 51716
rect 170811 50828 170877 50829
rect 170811 50764 170812 50828
rect 170876 50764 170877 50828
rect 170811 50763 170877 50764
rect 170627 50284 170693 50285
rect 170627 50220 170628 50284
rect 170692 50220 170693 50284
rect 170627 50219 170693 50220
rect 170443 48652 170509 48653
rect 170443 48588 170444 48652
rect 170508 48588 170509 48652
rect 170443 48587 170509 48588
rect 169339 48108 169405 48109
rect 169339 48044 169340 48108
rect 169404 48044 169405 48108
rect 169339 48043 169405 48044
rect 169155 9212 169221 9213
rect 169155 9148 169156 9212
rect 169220 9148 169221 9212
rect 169155 9147 169221 9148
rect 169342 9077 169402 48043
rect 170630 41989 170690 50219
rect 170627 41988 170693 41989
rect 170627 41924 170628 41988
rect 170692 41924 170693 41988
rect 170627 41923 170693 41924
rect 170814 41309 170874 50763
rect 170995 48788 171061 48789
rect 170995 48724 170996 48788
rect 171060 48724 171061 48788
rect 170995 48723 171061 48724
rect 170811 41308 170877 41309
rect 170811 41244 170812 41308
rect 170876 41244 170877 41308
rect 170811 41243 170877 41244
rect 170998 41173 171058 48723
rect 170995 41172 171061 41173
rect 170995 41108 170996 41172
rect 171060 41108 171061 41172
rect 170995 41107 171061 41108
rect 171834 29494 172454 50791
rect 173022 50285 173082 51715
rect 173203 51644 173269 51645
rect 173203 51580 173204 51644
rect 173268 51580 173269 51644
rect 173203 51579 173269 51580
rect 173206 51373 173266 51579
rect 173203 51372 173269 51373
rect 173203 51308 173204 51372
rect 173268 51308 173269 51372
rect 173203 51307 173269 51308
rect 173390 50965 173450 51851
rect 173574 51509 173634 52667
rect 194363 52324 194429 52325
rect 194363 52260 194364 52324
rect 194428 52260 194429 52324
rect 194363 52259 194429 52260
rect 194547 52324 194613 52325
rect 194547 52260 194548 52324
rect 194612 52260 194613 52324
rect 194547 52259 194613 52260
rect 194915 52324 194981 52325
rect 194915 52260 194916 52324
rect 194980 52260 194981 52324
rect 194915 52259 194981 52260
rect 193811 52188 193877 52189
rect 193811 52124 193812 52188
rect 193876 52124 193877 52188
rect 193811 52123 193877 52124
rect 174307 52052 174373 52053
rect 174307 51988 174308 52052
rect 174372 51988 174373 52052
rect 174307 51987 174373 51988
rect 175963 52052 176029 52053
rect 175963 51988 175964 52052
rect 176028 51988 176029 52052
rect 175963 51987 176029 51988
rect 173755 51916 173821 51917
rect 173755 51852 173756 51916
rect 173820 51852 173821 51916
rect 173755 51851 173821 51852
rect 174123 51916 174189 51917
rect 174123 51852 174124 51916
rect 174188 51852 174189 51916
rect 174123 51851 174189 51852
rect 173571 51508 173637 51509
rect 173571 51444 173572 51508
rect 173636 51444 173637 51508
rect 173571 51443 173637 51444
rect 173387 50964 173453 50965
rect 173387 50900 173388 50964
rect 173452 50900 173453 50964
rect 173387 50899 173453 50900
rect 173758 50693 173818 51851
rect 173755 50692 173821 50693
rect 173755 50628 173756 50692
rect 173820 50628 173821 50692
rect 173755 50627 173821 50628
rect 173019 50284 173085 50285
rect 173019 50220 173020 50284
rect 173084 50220 173085 50284
rect 173019 50219 173085 50220
rect 174126 50013 174186 51851
rect 174310 50013 174370 51987
rect 174859 51916 174925 51917
rect 174859 51852 174860 51916
rect 174924 51852 174925 51916
rect 174859 51851 174925 51852
rect 174491 51780 174557 51781
rect 174491 51716 174492 51780
rect 174556 51716 174557 51780
rect 174491 51715 174557 51716
rect 174494 51237 174554 51715
rect 174491 51236 174557 51237
rect 174491 51172 174492 51236
rect 174556 51172 174557 51236
rect 174491 51171 174557 51172
rect 174862 51101 174922 51851
rect 175411 51780 175477 51781
rect 175411 51716 175412 51780
rect 175476 51716 175477 51780
rect 175411 51715 175477 51716
rect 175414 51101 175474 51715
rect 174859 51100 174925 51101
rect 174859 51036 174860 51100
rect 174924 51036 174925 51100
rect 174859 51035 174925 51036
rect 175411 51100 175477 51101
rect 175411 51036 175412 51100
rect 175476 51036 175477 51100
rect 175411 51035 175477 51036
rect 175966 50421 176026 51987
rect 176331 51916 176397 51917
rect 176331 51852 176332 51916
rect 176396 51852 176397 51916
rect 176331 51851 176397 51852
rect 177987 51916 178053 51917
rect 177987 51852 177988 51916
rect 178052 51852 178053 51916
rect 177987 51851 178053 51852
rect 178907 51916 178973 51917
rect 178907 51852 178908 51916
rect 178972 51852 178973 51916
rect 178907 51851 178973 51852
rect 180011 51916 180077 51917
rect 180011 51852 180012 51916
rect 180076 51852 180077 51916
rect 180011 51851 180077 51852
rect 180379 51916 180445 51917
rect 180379 51852 180380 51916
rect 180444 51852 180445 51916
rect 180379 51851 180445 51852
rect 180931 51916 180997 51917
rect 180931 51852 180932 51916
rect 180996 51852 180997 51916
rect 180931 51851 180997 51852
rect 181299 51916 181365 51917
rect 181299 51852 181300 51916
rect 181364 51852 181365 51916
rect 181299 51851 181365 51852
rect 182771 51916 182837 51917
rect 182771 51852 182772 51916
rect 182836 51852 182837 51916
rect 182771 51851 182837 51852
rect 182955 51916 183021 51917
rect 182955 51852 182956 51916
rect 183020 51852 183021 51916
rect 183875 51916 183941 51917
rect 183875 51914 183876 51916
rect 182955 51851 183021 51852
rect 183694 51854 183876 51914
rect 175963 50420 176029 50421
rect 175963 50356 175964 50420
rect 176028 50356 176029 50420
rect 175963 50355 176029 50356
rect 174123 50012 174189 50013
rect 174123 49948 174124 50012
rect 174188 49948 174189 50012
rect 174123 49947 174189 49948
rect 174307 50012 174373 50013
rect 174307 49948 174308 50012
rect 174372 49948 174373 50012
rect 174307 49947 174373 49948
rect 176334 49605 176394 51851
rect 177990 50013 178050 51851
rect 178910 50149 178970 51851
rect 178907 50148 178973 50149
rect 178907 50084 178908 50148
rect 178972 50084 178973 50148
rect 178907 50083 178973 50084
rect 177987 50012 178053 50013
rect 177987 49948 177988 50012
rect 178052 49948 178053 50012
rect 177987 49947 178053 49948
rect 176331 49604 176397 49605
rect 176331 49540 176332 49604
rect 176396 49540 176397 49604
rect 176331 49539 176397 49540
rect 180014 47973 180074 51851
rect 180011 47972 180077 47973
rect 180011 47908 180012 47972
rect 180076 47908 180077 47972
rect 180011 47907 180077 47908
rect 180195 47972 180261 47973
rect 180195 47908 180196 47972
rect 180260 47908 180261 47972
rect 180195 47907 180261 47908
rect 171834 29258 171866 29494
rect 172102 29258 172186 29494
rect 172422 29258 172454 29494
rect 171834 29174 172454 29258
rect 171834 28938 171866 29174
rect 172102 28938 172186 29174
rect 172422 28938 172454 29174
rect 169339 9076 169405 9077
rect 169339 9012 169340 9076
rect 169404 9012 169405 9076
rect 169339 9011 169405 9012
rect 168971 5132 169037 5133
rect 168971 5068 168972 5132
rect 169036 5068 169037 5132
rect 168971 5067 169037 5068
rect 168114 -6342 168146 -6106
rect 168382 -6342 168466 -6106
rect 168702 -6342 168734 -6106
rect 168114 -6426 168734 -6342
rect 168114 -6662 168146 -6426
rect 168382 -6662 168466 -6426
rect 168702 -6662 168734 -6426
rect 168114 -7654 168734 -6662
rect 171834 -7066 172454 28938
rect 180198 25533 180258 47907
rect 180195 25532 180261 25533
rect 180195 25468 180196 25532
rect 180260 25468 180261 25532
rect 180195 25467 180261 25468
rect 180382 21317 180442 51851
rect 180563 47972 180629 47973
rect 180563 47908 180564 47972
rect 180628 47908 180629 47972
rect 180563 47907 180629 47908
rect 180379 21316 180445 21317
rect 180379 21252 180380 21316
rect 180444 21252 180445 21316
rect 180379 21251 180445 21252
rect 180566 14789 180626 47907
rect 180934 18733 180994 51851
rect 181302 48517 181362 51851
rect 181299 48516 181365 48517
rect 181299 48452 181300 48516
rect 181364 48452 181365 48516
rect 181299 48451 181365 48452
rect 181115 48380 181181 48381
rect 181115 48316 181116 48380
rect 181180 48316 181181 48380
rect 181115 48315 181181 48316
rect 181118 18869 181178 48315
rect 181299 47972 181365 47973
rect 181299 47908 181300 47972
rect 181364 47908 181365 47972
rect 181299 47907 181365 47908
rect 181115 18868 181181 18869
rect 181115 18804 181116 18868
rect 181180 18804 181181 18868
rect 181115 18803 181181 18804
rect 180931 18732 180997 18733
rect 180931 18668 180932 18732
rect 180996 18668 180997 18732
rect 180931 18667 180997 18668
rect 181302 17373 181362 47907
rect 181794 39454 182414 50791
rect 182587 48516 182653 48517
rect 182587 48452 182588 48516
rect 182652 48452 182653 48516
rect 182587 48451 182653 48452
rect 181794 39218 181826 39454
rect 182062 39218 182146 39454
rect 182382 39218 182414 39454
rect 181794 39134 182414 39218
rect 181794 38898 181826 39134
rect 182062 38898 182146 39134
rect 182382 38898 182414 39134
rect 181299 17372 181365 17373
rect 181299 17308 181300 17372
rect 181364 17308 181365 17372
rect 181299 17307 181365 17308
rect 180563 14788 180629 14789
rect 180563 14724 180564 14788
rect 180628 14724 180629 14788
rect 180563 14723 180629 14724
rect 171834 -7302 171866 -7066
rect 172102 -7302 172186 -7066
rect 172422 -7302 172454 -7066
rect 171834 -7386 172454 -7302
rect 171834 -7622 171866 -7386
rect 172102 -7622 172186 -7386
rect 172422 -7622 172454 -7386
rect 171834 -7654 172454 -7622
rect 181794 3454 182414 38898
rect 182590 35189 182650 48451
rect 182774 37909 182834 51851
rect 182958 49741 183018 51851
rect 182955 49740 183021 49741
rect 182955 49676 182956 49740
rect 183020 49676 183021 49740
rect 182955 49675 183021 49676
rect 182955 49060 183021 49061
rect 182955 48996 182956 49060
rect 183020 48996 183021 49060
rect 182955 48995 183021 48996
rect 182958 44981 183018 48995
rect 183139 48788 183205 48789
rect 183139 48724 183140 48788
rect 183204 48724 183205 48788
rect 183139 48723 183205 48724
rect 182955 44980 183021 44981
rect 182955 44916 182956 44980
rect 183020 44916 183021 44980
rect 182955 44915 183021 44916
rect 183142 43485 183202 48723
rect 183139 43484 183205 43485
rect 183139 43420 183140 43484
rect 183204 43420 183205 43484
rect 183139 43419 183205 43420
rect 182771 37908 182837 37909
rect 182771 37844 182772 37908
rect 182836 37844 182837 37908
rect 182771 37843 182837 37844
rect 182587 35188 182653 35189
rect 182587 35124 182588 35188
rect 182652 35124 182653 35188
rect 182587 35123 182653 35124
rect 183694 6221 183754 51854
rect 183875 51852 183876 51854
rect 183940 51852 183941 51916
rect 183875 51851 183941 51852
rect 184427 51916 184493 51917
rect 184427 51852 184428 51916
rect 184492 51852 184493 51916
rect 184427 51851 184493 51852
rect 184611 51916 184677 51917
rect 184611 51852 184612 51916
rect 184676 51852 184677 51916
rect 185347 51916 185413 51917
rect 185347 51914 185348 51916
rect 184611 51851 184677 51852
rect 185166 51854 185348 51914
rect 183875 49740 183941 49741
rect 183875 49676 183876 49740
rect 183940 49676 183941 49740
rect 183875 49675 183941 49676
rect 183691 6220 183757 6221
rect 183691 6156 183692 6220
rect 183756 6156 183757 6220
rect 183691 6155 183757 6156
rect 183878 4861 183938 49675
rect 184430 48789 184490 51851
rect 184427 48788 184493 48789
rect 184427 48724 184428 48788
rect 184492 48724 184493 48788
rect 184427 48723 184493 48724
rect 184614 48517 184674 51851
rect 185166 48517 185226 51854
rect 185347 51852 185348 51854
rect 185412 51852 185413 51916
rect 185347 51851 185413 51852
rect 187003 51916 187069 51917
rect 187003 51852 187004 51916
rect 187068 51852 187069 51916
rect 187003 51851 187069 51852
rect 188475 51916 188541 51917
rect 188475 51852 188476 51916
rect 188540 51852 188541 51916
rect 189027 51916 189093 51917
rect 189027 51914 189028 51916
rect 188475 51851 188541 51852
rect 188846 51854 189028 51914
rect 184611 48516 184677 48517
rect 184611 48452 184612 48516
rect 184676 48452 184677 48516
rect 184611 48451 184677 48452
rect 185163 48516 185229 48517
rect 185163 48452 185164 48516
rect 185228 48452 185229 48516
rect 185163 48451 185229 48452
rect 185347 48516 185413 48517
rect 185347 48452 185348 48516
rect 185412 48452 185413 48516
rect 185347 48451 185413 48452
rect 185163 48380 185229 48381
rect 185163 48316 185164 48380
rect 185228 48316 185229 48380
rect 185163 48315 185229 48316
rect 185166 21453 185226 48315
rect 185350 44437 185410 48451
rect 185347 44436 185413 44437
rect 185347 44372 185348 44436
rect 185412 44372 185413 44436
rect 185347 44371 185413 44372
rect 185514 43174 186134 50791
rect 187006 50149 187066 51851
rect 187003 50148 187069 50149
rect 187003 50084 187004 50148
rect 187068 50084 187069 50148
rect 187003 50083 187069 50084
rect 187003 48788 187069 48789
rect 187003 48724 187004 48788
rect 187068 48724 187069 48788
rect 187003 48723 187069 48724
rect 187006 45525 187066 48723
rect 187187 48652 187253 48653
rect 187187 48588 187188 48652
rect 187252 48588 187253 48652
rect 187187 48587 187253 48588
rect 187003 45524 187069 45525
rect 187003 45460 187004 45524
rect 187068 45460 187069 45524
rect 187003 45459 187069 45460
rect 185514 42938 185546 43174
rect 185782 42938 185866 43174
rect 186102 42938 186134 43174
rect 185514 42854 186134 42938
rect 185514 42618 185546 42854
rect 185782 42618 185866 42854
rect 186102 42618 186134 42854
rect 185163 21452 185229 21453
rect 185163 21388 185164 21452
rect 185228 21388 185229 21452
rect 185163 21387 185229 21388
rect 185514 7174 186134 42618
rect 187190 17781 187250 48587
rect 187555 48516 187621 48517
rect 187555 48452 187556 48516
rect 187620 48452 187621 48516
rect 187555 48451 187621 48452
rect 187371 48380 187437 48381
rect 187371 48316 187372 48380
rect 187436 48316 187437 48380
rect 187371 48315 187437 48316
rect 187187 17780 187253 17781
rect 187187 17716 187188 17780
rect 187252 17716 187253 17780
rect 187187 17715 187253 17716
rect 187374 17237 187434 48315
rect 187371 17236 187437 17237
rect 187371 17172 187372 17236
rect 187436 17172 187437 17236
rect 187371 17171 187437 17172
rect 185514 6938 185546 7174
rect 185782 6938 185866 7174
rect 186102 6938 186134 7174
rect 185514 6854 186134 6938
rect 185514 6618 185546 6854
rect 185782 6618 185866 6854
rect 186102 6618 186134 6854
rect 183875 4860 183941 4861
rect 183875 4796 183876 4860
rect 183940 4796 183941 4860
rect 183875 4795 183941 4796
rect 181794 3218 181826 3454
rect 182062 3218 182146 3454
rect 182382 3218 182414 3454
rect 181794 3134 182414 3218
rect 181794 2898 181826 3134
rect 182062 2898 182146 3134
rect 182382 2898 182414 3134
rect 181794 -346 182414 2898
rect 181794 -582 181826 -346
rect 182062 -582 182146 -346
rect 182382 -582 182414 -346
rect 181794 -666 182414 -582
rect 181794 -902 181826 -666
rect 182062 -902 182146 -666
rect 182382 -902 182414 -666
rect 181794 -7654 182414 -902
rect 185514 -1306 186134 6618
rect 187558 4861 187618 48451
rect 188478 42125 188538 51851
rect 188659 48380 188725 48381
rect 188659 48316 188660 48380
rect 188724 48316 188725 48380
rect 188659 48315 188725 48316
rect 188475 42124 188541 42125
rect 188475 42060 188476 42124
rect 188540 42060 188541 42124
rect 188475 42059 188541 42060
rect 188662 6085 188722 48315
rect 188659 6084 188725 6085
rect 188659 6020 188660 6084
rect 188724 6020 188725 6084
rect 188659 6019 188725 6020
rect 187555 4860 187621 4861
rect 187555 4796 187556 4860
rect 187620 4796 187621 4860
rect 187555 4795 187621 4796
rect 188846 3637 188906 51854
rect 189027 51852 189028 51854
rect 189092 51852 189093 51916
rect 189027 51851 189093 51852
rect 192707 51916 192773 51917
rect 192707 51852 192708 51916
rect 192772 51852 192773 51916
rect 192707 51851 192773 51852
rect 189027 48652 189093 48653
rect 189027 48588 189028 48652
rect 189092 48588 189093 48652
rect 189027 48587 189093 48588
rect 189030 46341 189090 48587
rect 189234 46894 189854 50791
rect 191419 50148 191485 50149
rect 191419 50084 191420 50148
rect 191484 50084 191485 50148
rect 191419 50083 191485 50084
rect 190131 50012 190197 50013
rect 190131 49948 190132 50012
rect 190196 49948 190197 50012
rect 190131 49947 190197 49948
rect 191051 50012 191117 50013
rect 191051 49948 191052 50012
rect 191116 49948 191117 50012
rect 191051 49947 191117 49948
rect 189234 46658 189266 46894
rect 189502 46658 189586 46894
rect 189822 46658 189854 46894
rect 189234 46574 189854 46658
rect 189027 46340 189093 46341
rect 189027 46276 189028 46340
rect 189092 46276 189093 46340
rect 189027 46275 189093 46276
rect 189234 46338 189266 46574
rect 189502 46338 189586 46574
rect 189822 46338 189854 46574
rect 189234 10894 189854 46338
rect 190134 43485 190194 49947
rect 190315 48380 190381 48381
rect 190315 48316 190316 48380
rect 190380 48316 190381 48380
rect 190315 48315 190381 48316
rect 190131 43484 190197 43485
rect 190131 43420 190132 43484
rect 190196 43420 190197 43484
rect 190131 43419 190197 43420
rect 189234 10658 189266 10894
rect 189502 10658 189586 10894
rect 189822 10658 189854 10894
rect 189234 10574 189854 10658
rect 189234 10338 189266 10574
rect 189502 10338 189586 10574
rect 189822 10338 189854 10574
rect 188843 3636 188909 3637
rect 188843 3572 188844 3636
rect 188908 3572 188909 3636
rect 188843 3571 188909 3572
rect 185514 -1542 185546 -1306
rect 185782 -1542 185866 -1306
rect 186102 -1542 186134 -1306
rect 185514 -1626 186134 -1542
rect 185514 -1862 185546 -1626
rect 185782 -1862 185866 -1626
rect 186102 -1862 186134 -1626
rect 185514 -7654 186134 -1862
rect 189234 -2266 189854 10338
rect 190318 6901 190378 48315
rect 191054 36549 191114 49947
rect 191235 49876 191301 49877
rect 191235 49812 191236 49876
rect 191300 49812 191301 49876
rect 191235 49811 191301 49812
rect 191051 36548 191117 36549
rect 191051 36484 191052 36548
rect 191116 36484 191117 36548
rect 191051 36483 191117 36484
rect 191238 13565 191298 49811
rect 191235 13564 191301 13565
rect 191235 13500 191236 13564
rect 191300 13500 191301 13564
rect 191235 13499 191301 13500
rect 191422 13429 191482 50083
rect 191603 50012 191669 50013
rect 191603 49948 191604 50012
rect 191668 49948 191669 50012
rect 191603 49947 191669 49948
rect 191419 13428 191485 13429
rect 191419 13364 191420 13428
rect 191484 13364 191485 13428
rect 191419 13363 191485 13364
rect 190315 6900 190381 6901
rect 190315 6836 190316 6900
rect 190380 6836 190381 6900
rect 190315 6835 190381 6836
rect 191606 3773 191666 49947
rect 192155 48788 192221 48789
rect 192155 48724 192156 48788
rect 192220 48724 192221 48788
rect 192155 48723 192221 48724
rect 192158 35597 192218 48723
rect 192339 48652 192405 48653
rect 192339 48588 192340 48652
rect 192404 48588 192405 48652
rect 192339 48587 192405 48588
rect 192155 35596 192221 35597
rect 192155 35532 192156 35596
rect 192220 35532 192221 35596
rect 192155 35531 192221 35532
rect 192342 24445 192402 48587
rect 192523 48516 192589 48517
rect 192523 48452 192524 48516
rect 192588 48452 192589 48516
rect 192523 48451 192589 48452
rect 192339 24444 192405 24445
rect 192339 24380 192340 24444
rect 192404 24380 192405 24444
rect 192339 24379 192405 24380
rect 192526 17645 192586 48451
rect 192523 17644 192589 17645
rect 192523 17580 192524 17644
rect 192588 17580 192589 17644
rect 192523 17579 192589 17580
rect 192710 13293 192770 51851
rect 192954 50614 193574 52068
rect 192954 50378 192986 50614
rect 193222 50378 193306 50614
rect 193542 50378 193574 50614
rect 192954 50294 193574 50378
rect 192954 50058 192986 50294
rect 193222 50058 193306 50294
rect 193542 50058 193574 50294
rect 192954 14614 193574 50058
rect 193814 47429 193874 52123
rect 194179 51916 194245 51917
rect 194179 51852 194180 51916
rect 194244 51852 194245 51916
rect 194179 51851 194245 51852
rect 193995 50148 194061 50149
rect 193995 50084 193996 50148
rect 194060 50084 194061 50148
rect 193995 50083 194061 50084
rect 193811 47428 193877 47429
rect 193811 47364 193812 47428
rect 193876 47364 193877 47428
rect 193811 47363 193877 47364
rect 193998 34237 194058 50083
rect 194182 50013 194242 51851
rect 194179 50012 194245 50013
rect 194179 49948 194180 50012
rect 194244 49948 194245 50012
rect 194179 49947 194245 49948
rect 194366 49741 194426 52259
rect 194550 52053 194610 52259
rect 194731 52188 194797 52189
rect 194731 52124 194732 52188
rect 194796 52124 194797 52188
rect 194731 52123 194797 52124
rect 194547 52052 194613 52053
rect 194547 51988 194548 52052
rect 194612 51988 194613 52052
rect 194547 51987 194613 51988
rect 194363 49740 194429 49741
rect 194363 49676 194364 49740
rect 194428 49676 194429 49740
rect 194363 49675 194429 49676
rect 194363 47564 194429 47565
rect 194363 47500 194364 47564
rect 194428 47500 194429 47564
rect 194363 47499 194429 47500
rect 194179 47428 194245 47429
rect 194179 47364 194180 47428
rect 194244 47364 194245 47428
rect 194179 47363 194245 47364
rect 193995 34236 194061 34237
rect 193995 34172 193996 34236
rect 194060 34172 194061 34236
rect 193995 34171 194061 34172
rect 194182 18597 194242 47363
rect 194179 18596 194245 18597
rect 194179 18532 194180 18596
rect 194244 18532 194245 18596
rect 194179 18531 194245 18532
rect 192954 14378 192986 14614
rect 193222 14378 193306 14614
rect 193542 14378 193574 14614
rect 192954 14294 193574 14378
rect 192954 14058 192986 14294
rect 193222 14058 193306 14294
rect 193542 14058 193574 14294
rect 192707 13292 192773 13293
rect 192707 13228 192708 13292
rect 192772 13228 192773 13292
rect 192707 13227 192773 13228
rect 191603 3772 191669 3773
rect 191603 3708 191604 3772
rect 191668 3708 191669 3772
rect 191603 3707 191669 3708
rect 189234 -2502 189266 -2266
rect 189502 -2502 189586 -2266
rect 189822 -2502 189854 -2266
rect 189234 -2586 189854 -2502
rect 189234 -2822 189266 -2586
rect 189502 -2822 189586 -2586
rect 189822 -2822 189854 -2586
rect 189234 -7654 189854 -2822
rect 192954 -3226 193574 14058
rect 194366 6765 194426 47499
rect 194734 47429 194794 52123
rect 194731 47428 194797 47429
rect 194731 47364 194732 47428
rect 194796 47364 194797 47428
rect 194731 47363 194797 47364
rect 194918 47293 194978 52259
rect 196203 52052 196269 52053
rect 196203 51988 196204 52052
rect 196268 51988 196269 52052
rect 196203 51987 196269 51988
rect 195099 51916 195165 51917
rect 195099 51852 195100 51916
rect 195164 51852 195165 51916
rect 195099 51851 195165 51852
rect 195651 51916 195717 51917
rect 195651 51852 195652 51916
rect 195716 51852 195717 51916
rect 195651 51851 195717 51852
rect 195102 47565 195162 51851
rect 195654 51090 195714 51851
rect 195470 51030 195714 51090
rect 195099 47564 195165 47565
rect 195099 47500 195100 47564
rect 195164 47500 195165 47564
rect 195099 47499 195165 47500
rect 195283 47428 195349 47429
rect 195283 47364 195284 47428
rect 195348 47364 195349 47428
rect 195283 47363 195349 47364
rect 194915 47292 194981 47293
rect 194915 47228 194916 47292
rect 194980 47228 194981 47292
rect 194915 47227 194981 47228
rect 195286 37909 195346 47363
rect 195283 37908 195349 37909
rect 195283 37844 195284 37908
rect 195348 37844 195349 37908
rect 195283 37843 195349 37844
rect 195470 29885 195530 51030
rect 196206 49330 196266 51987
rect 196387 51916 196453 51917
rect 196387 51852 196388 51916
rect 196452 51852 196453 51916
rect 196387 51851 196453 51852
rect 196390 49741 196450 51851
rect 196387 49740 196453 49741
rect 196387 49676 196388 49740
rect 196452 49676 196453 49740
rect 196387 49675 196453 49676
rect 196206 49270 196450 49330
rect 196203 48652 196269 48653
rect 196203 48588 196204 48652
rect 196268 48588 196269 48652
rect 196203 48587 196269 48588
rect 195651 47700 195717 47701
rect 195651 47636 195652 47700
rect 195716 47636 195717 47700
rect 195651 47635 195717 47636
rect 195467 29884 195533 29885
rect 195467 29820 195468 29884
rect 195532 29820 195533 29884
rect 195467 29819 195533 29820
rect 195654 14653 195714 47635
rect 195835 47564 195901 47565
rect 195835 47500 195836 47564
rect 195900 47500 195901 47564
rect 195835 47499 195901 47500
rect 195651 14652 195717 14653
rect 195651 14588 195652 14652
rect 195716 14588 195717 14652
rect 195651 14587 195717 14588
rect 195838 13157 195898 47499
rect 196206 29749 196266 48587
rect 196203 29748 196269 29749
rect 196203 29684 196204 29748
rect 196268 29684 196269 29748
rect 196203 29683 196269 29684
rect 196390 21861 196450 49270
rect 196387 21860 196453 21861
rect 196387 21796 196388 21860
rect 196452 21796 196453 21860
rect 196387 21795 196453 21796
rect 196674 18334 197294 53778
rect 200394 238054 201014 270287
rect 200394 237818 200426 238054
rect 200662 237818 200746 238054
rect 200982 237818 201014 238054
rect 200394 237734 201014 237818
rect 200394 237498 200426 237734
rect 200662 237498 200746 237734
rect 200982 237498 201014 237734
rect 200394 202054 201014 237498
rect 200394 201818 200426 202054
rect 200662 201818 200746 202054
rect 200982 201818 201014 202054
rect 200394 201734 201014 201818
rect 200394 201498 200426 201734
rect 200662 201498 200746 201734
rect 200982 201498 201014 201734
rect 200394 166054 201014 201498
rect 200394 165818 200426 166054
rect 200662 165818 200746 166054
rect 200982 165818 201014 166054
rect 200394 165734 201014 165818
rect 200394 165498 200426 165734
rect 200662 165498 200746 165734
rect 200982 165498 201014 165734
rect 200394 130054 201014 165498
rect 200394 129818 200426 130054
rect 200662 129818 200746 130054
rect 200982 129818 201014 130054
rect 200394 129734 201014 129818
rect 200394 129498 200426 129734
rect 200662 129498 200746 129734
rect 200982 129498 201014 129734
rect 200394 94054 201014 129498
rect 200394 93818 200426 94054
rect 200662 93818 200746 94054
rect 200982 93818 201014 94054
rect 200394 93734 201014 93818
rect 200394 93498 200426 93734
rect 200662 93498 200746 93734
rect 200982 93498 201014 93734
rect 200394 58054 201014 93498
rect 200394 57818 200426 58054
rect 200662 57818 200746 58054
rect 200982 57818 201014 58054
rect 200394 57734 201014 57818
rect 200394 57498 200426 57734
rect 200662 57498 200746 57734
rect 200982 57498 201014 57734
rect 198227 51916 198293 51917
rect 198227 51852 198228 51916
rect 198292 51852 198293 51916
rect 198227 51851 198293 51852
rect 198595 51916 198661 51917
rect 198595 51852 198596 51916
rect 198660 51852 198661 51916
rect 198595 51851 198661 51852
rect 200067 51916 200133 51917
rect 200067 51852 200068 51916
rect 200132 51852 200133 51916
rect 200067 51851 200133 51852
rect 198043 48652 198109 48653
rect 198043 48588 198044 48652
rect 198108 48588 198109 48652
rect 198043 48587 198109 48588
rect 198046 32741 198106 48587
rect 198043 32740 198109 32741
rect 198043 32676 198044 32740
rect 198108 32676 198109 32740
rect 198043 32675 198109 32676
rect 198230 21725 198290 51851
rect 198411 48924 198477 48925
rect 198411 48860 198412 48924
rect 198476 48860 198477 48924
rect 198411 48859 198477 48860
rect 198227 21724 198293 21725
rect 198227 21660 198228 21724
rect 198292 21660 198293 21724
rect 198227 21659 198293 21660
rect 196674 18098 196706 18334
rect 196942 18098 197026 18334
rect 197262 18098 197294 18334
rect 196674 18014 197294 18098
rect 196674 17778 196706 18014
rect 196942 17778 197026 18014
rect 197262 17778 197294 18014
rect 195835 13156 195901 13157
rect 195835 13092 195836 13156
rect 195900 13092 195901 13156
rect 195835 13091 195901 13092
rect 194363 6764 194429 6765
rect 194363 6700 194364 6764
rect 194428 6700 194429 6764
rect 194363 6699 194429 6700
rect 192954 -3462 192986 -3226
rect 193222 -3462 193306 -3226
rect 193542 -3462 193574 -3226
rect 192954 -3546 193574 -3462
rect 192954 -3782 192986 -3546
rect 193222 -3782 193306 -3546
rect 193542 -3782 193574 -3546
rect 192954 -7654 193574 -3782
rect 196674 -4186 197294 17778
rect 198414 16013 198474 48859
rect 198411 16012 198477 16013
rect 198411 15948 198412 16012
rect 198476 15948 198477 16012
rect 198411 15947 198477 15948
rect 198598 6629 198658 51851
rect 199331 48652 199397 48653
rect 199331 48588 199332 48652
rect 199396 48588 199397 48652
rect 199331 48587 199397 48588
rect 199334 31109 199394 48587
rect 199699 48516 199765 48517
rect 199699 48452 199700 48516
rect 199764 48452 199765 48516
rect 199699 48451 199765 48452
rect 199515 48380 199581 48381
rect 199515 48316 199516 48380
rect 199580 48316 199581 48380
rect 199515 48315 199581 48316
rect 199331 31108 199397 31109
rect 199331 31044 199332 31108
rect 199396 31044 199397 31108
rect 199331 31043 199397 31044
rect 199518 28525 199578 48315
rect 199515 28524 199581 28525
rect 199515 28460 199516 28524
rect 199580 28460 199581 28524
rect 199515 28459 199581 28460
rect 199702 21589 199762 48451
rect 199883 48380 199949 48381
rect 199883 48316 199884 48380
rect 199948 48316 199949 48380
rect 199883 48315 199949 48316
rect 199699 21588 199765 21589
rect 199699 21524 199700 21588
rect 199764 21524 199765 21588
rect 199699 21523 199765 21524
rect 198595 6628 198661 6629
rect 198595 6564 198596 6628
rect 198660 6564 198661 6628
rect 198595 6563 198661 6564
rect 199886 6493 199946 48315
rect 200070 41445 200130 51851
rect 200067 41444 200133 41445
rect 200067 41380 200068 41444
rect 200132 41380 200133 41444
rect 200067 41379 200133 41380
rect 200067 36004 200133 36005
rect 200067 35940 200068 36004
rect 200132 35940 200133 36004
rect 200067 35939 200133 35940
rect 200070 35461 200130 35939
rect 200067 35460 200133 35461
rect 200067 35396 200068 35460
rect 200132 35396 200133 35460
rect 200067 35395 200133 35396
rect 200394 22054 201014 57498
rect 204114 241774 204734 270287
rect 204114 241538 204146 241774
rect 204382 241538 204466 241774
rect 204702 241538 204734 241774
rect 204114 241454 204734 241538
rect 204114 241218 204146 241454
rect 204382 241218 204466 241454
rect 204702 241218 204734 241454
rect 204114 205774 204734 241218
rect 204114 205538 204146 205774
rect 204382 205538 204466 205774
rect 204702 205538 204734 205774
rect 204114 205454 204734 205538
rect 204114 205218 204146 205454
rect 204382 205218 204466 205454
rect 204702 205218 204734 205454
rect 204114 169774 204734 205218
rect 204114 169538 204146 169774
rect 204382 169538 204466 169774
rect 204702 169538 204734 169774
rect 204114 169454 204734 169538
rect 204114 169218 204146 169454
rect 204382 169218 204466 169454
rect 204702 169218 204734 169454
rect 204114 133774 204734 169218
rect 204114 133538 204146 133774
rect 204382 133538 204466 133774
rect 204702 133538 204734 133774
rect 204114 133454 204734 133538
rect 204114 133218 204146 133454
rect 204382 133218 204466 133454
rect 204702 133218 204734 133454
rect 204114 97774 204734 133218
rect 207834 245494 208454 270068
rect 207834 245258 207866 245494
rect 208102 245258 208186 245494
rect 208422 245258 208454 245494
rect 207834 245174 208454 245258
rect 207834 244938 207866 245174
rect 208102 244938 208186 245174
rect 208422 244938 208454 245174
rect 207834 209494 208454 244938
rect 207834 209258 207866 209494
rect 208102 209258 208186 209494
rect 208422 209258 208454 209494
rect 207834 209174 208454 209258
rect 207834 208938 207866 209174
rect 208102 208938 208186 209174
rect 208422 208938 208454 209174
rect 207834 173494 208454 208938
rect 207834 173258 207866 173494
rect 208102 173258 208186 173494
rect 208422 173258 208454 173494
rect 207834 173174 208454 173258
rect 207834 172938 207866 173174
rect 208102 172938 208186 173174
rect 208422 172938 208454 173174
rect 207834 137494 208454 172938
rect 207834 137258 207866 137494
rect 208102 137258 208186 137494
rect 208422 137258 208454 137494
rect 207834 137174 208454 137258
rect 207834 136938 207866 137174
rect 208102 136938 208186 137174
rect 208422 136938 208454 137174
rect 207834 131900 208454 136938
rect 217794 255454 218414 290898
rect 217794 255218 217826 255454
rect 218062 255218 218146 255454
rect 218382 255218 218414 255454
rect 217794 255134 218414 255218
rect 217794 254898 217826 255134
rect 218062 254898 218146 255134
rect 218382 254898 218414 255134
rect 217794 219454 218414 254898
rect 217794 219218 217826 219454
rect 218062 219218 218146 219454
rect 218382 219218 218414 219454
rect 217794 219134 218414 219218
rect 217794 218898 217826 219134
rect 218062 218898 218146 219134
rect 218382 218898 218414 219134
rect 217794 183454 218414 218898
rect 217794 183218 217826 183454
rect 218062 183218 218146 183454
rect 218382 183218 218414 183454
rect 217794 183134 218414 183218
rect 217794 182898 217826 183134
rect 218062 182898 218146 183134
rect 218382 182898 218414 183134
rect 217794 147454 218414 182898
rect 217794 147218 217826 147454
rect 218062 147218 218146 147454
rect 218382 147218 218414 147454
rect 217794 147134 218414 147218
rect 217794 146898 217826 147134
rect 218062 146898 218146 147134
rect 218382 146898 218414 147134
rect 208288 115174 208608 115206
rect 208288 114938 208330 115174
rect 208566 114938 208608 115174
rect 208288 114854 208608 114938
rect 208288 114618 208330 114854
rect 208566 114618 208608 114854
rect 208288 114586 208608 114618
rect 204114 97538 204146 97774
rect 204382 97538 204466 97774
rect 204702 97538 204734 97774
rect 204114 97454 204734 97538
rect 204114 97218 204146 97454
rect 204382 97218 204466 97454
rect 204702 97218 204734 97454
rect 204114 61774 204734 97218
rect 217794 111454 218414 146898
rect 217794 111218 217826 111454
rect 218062 111218 218146 111454
rect 218382 111218 218414 111454
rect 217794 111134 218414 111218
rect 217794 110898 217826 111134
rect 218062 110898 218146 111134
rect 218382 110898 218414 111134
rect 208288 79174 208608 79206
rect 208288 78938 208330 79174
rect 208566 78938 208608 79174
rect 208288 78854 208608 78938
rect 208288 78618 208330 78854
rect 208566 78618 208608 78854
rect 208288 78586 208608 78618
rect 204114 61538 204146 61774
rect 204382 61538 204466 61774
rect 204702 61538 204734 61774
rect 204114 61454 204734 61538
rect 204114 61218 204146 61454
rect 204382 61218 204466 61454
rect 204702 61218 204734 61454
rect 202091 51916 202157 51917
rect 202091 51852 202092 51916
rect 202156 51852 202157 51916
rect 202091 51851 202157 51852
rect 203379 51916 203445 51917
rect 203379 51852 203380 51916
rect 203444 51852 203445 51916
rect 203379 51851 203445 51852
rect 202094 49741 202154 51851
rect 202091 49740 202157 49741
rect 202091 49676 202092 49740
rect 202156 49676 202157 49740
rect 202091 49675 202157 49676
rect 202091 48924 202157 48925
rect 202091 48860 202092 48924
rect 202156 48860 202157 48924
rect 202091 48859 202157 48860
rect 203195 48924 203261 48925
rect 203195 48860 203196 48924
rect 203260 48860 203261 48924
rect 203195 48859 203261 48860
rect 201355 48380 201421 48381
rect 201355 48316 201356 48380
rect 201420 48316 201421 48380
rect 201355 48315 201421 48316
rect 200394 21818 200426 22054
rect 200662 21818 200746 22054
rect 200982 21818 201014 22054
rect 200394 21734 201014 21818
rect 200394 21498 200426 21734
rect 200662 21498 200746 21734
rect 200982 21498 201014 21734
rect 199883 6492 199949 6493
rect 199883 6428 199884 6492
rect 199948 6428 199949 6492
rect 199883 6427 199949 6428
rect 196674 -4422 196706 -4186
rect 196942 -4422 197026 -4186
rect 197262 -4422 197294 -4186
rect 196674 -4506 197294 -4422
rect 196674 -4742 196706 -4506
rect 196942 -4742 197026 -4506
rect 197262 -4742 197294 -4506
rect 196674 -7654 197294 -4742
rect 200394 -5146 201014 21498
rect 201358 13021 201418 48315
rect 202094 34101 202154 48859
rect 202275 48652 202341 48653
rect 202275 48588 202276 48652
rect 202340 48588 202341 48652
rect 202275 48587 202341 48588
rect 202091 34100 202157 34101
rect 202091 34036 202092 34100
rect 202156 34036 202157 34100
rect 202091 34035 202157 34036
rect 202278 20093 202338 48587
rect 202459 48516 202525 48517
rect 202459 48452 202460 48516
rect 202524 48452 202525 48516
rect 202459 48451 202525 48452
rect 202275 20092 202341 20093
rect 202275 20028 202276 20092
rect 202340 20028 202341 20092
rect 202275 20027 202341 20028
rect 202462 14517 202522 48451
rect 202643 48380 202709 48381
rect 202643 48316 202644 48380
rect 202708 48316 202709 48380
rect 202643 48315 202709 48316
rect 202459 14516 202525 14517
rect 202459 14452 202460 14516
rect 202524 14452 202525 14516
rect 202459 14451 202525 14452
rect 201355 13020 201421 13021
rect 201355 12956 201356 13020
rect 201420 12956 201421 13020
rect 201355 12955 201421 12956
rect 202646 6357 202706 48315
rect 203198 29613 203258 48859
rect 203195 29612 203261 29613
rect 203195 29548 203196 29612
rect 203260 29548 203261 29612
rect 203195 29547 203261 29548
rect 203382 21453 203442 51851
rect 203563 50148 203629 50149
rect 203563 50084 203564 50148
rect 203628 50084 203629 50148
rect 203563 50083 203629 50084
rect 203379 21452 203445 21453
rect 203379 21388 203380 21452
rect 203444 21388 203445 21452
rect 203379 21387 203445 21388
rect 203566 15877 203626 50083
rect 203747 48380 203813 48381
rect 203747 48316 203748 48380
rect 203812 48316 203813 48380
rect 203747 48315 203813 48316
rect 203563 15876 203629 15877
rect 203563 15812 203564 15876
rect 203628 15812 203629 15876
rect 203563 15811 203629 15812
rect 202643 6356 202709 6357
rect 202643 6292 202644 6356
rect 202708 6292 202709 6356
rect 202643 6291 202709 6292
rect 203750 4997 203810 48315
rect 204114 25774 204734 61218
rect 217794 75454 218414 110898
rect 217794 75218 217826 75454
rect 218062 75218 218146 75454
rect 218382 75218 218414 75454
rect 217794 75134 218414 75218
rect 217794 74898 217826 75134
rect 218062 74898 218146 75134
rect 218382 74898 218414 75134
rect 208715 52868 208781 52869
rect 208715 52804 208716 52868
rect 208780 52804 208781 52868
rect 208715 52803 208781 52804
rect 208718 52325 208778 52803
rect 208715 52324 208781 52325
rect 208715 52260 208716 52324
rect 208780 52260 208781 52324
rect 208715 52259 208781 52260
rect 204851 52188 204917 52189
rect 204851 52124 204852 52188
rect 204916 52124 204917 52188
rect 204851 52123 204917 52124
rect 205587 52188 205653 52189
rect 205587 52124 205588 52188
rect 205652 52124 205653 52188
rect 205587 52123 205653 52124
rect 204854 49877 204914 52123
rect 205035 51916 205101 51917
rect 205035 51852 205036 51916
rect 205100 51852 205101 51916
rect 205403 51916 205469 51917
rect 205403 51914 205404 51916
rect 205035 51851 205101 51852
rect 205222 51854 205404 51914
rect 205038 50149 205098 51851
rect 205035 50148 205101 50149
rect 205035 50084 205036 50148
rect 205100 50084 205101 50148
rect 205035 50083 205101 50084
rect 204851 49876 204917 49877
rect 204851 49812 204852 49876
rect 204916 49812 204917 49876
rect 204851 49811 204917 49812
rect 205035 48380 205101 48381
rect 205035 48316 205036 48380
rect 205100 48316 205101 48380
rect 205035 48315 205101 48316
rect 205038 27029 205098 48315
rect 205035 27028 205101 27029
rect 205035 26964 205036 27028
rect 205100 26964 205101 27028
rect 205035 26963 205101 26964
rect 204114 25538 204146 25774
rect 204382 25538 204466 25774
rect 204702 25538 204734 25774
rect 204114 25454 204734 25538
rect 204114 25218 204146 25454
rect 204382 25218 204466 25454
rect 204702 25218 204734 25454
rect 203747 4996 203813 4997
rect 203747 4932 203748 4996
rect 203812 4932 203813 4996
rect 203747 4931 203813 4932
rect 200394 -5382 200426 -5146
rect 200662 -5382 200746 -5146
rect 200982 -5382 201014 -5146
rect 200394 -5466 201014 -5382
rect 200394 -5702 200426 -5466
rect 200662 -5702 200746 -5466
rect 200982 -5702 201014 -5466
rect 200394 -7654 201014 -5702
rect 204114 -6106 204734 25218
rect 205222 19957 205282 51854
rect 205403 51852 205404 51854
rect 205468 51852 205469 51916
rect 205403 51851 205469 51852
rect 205590 51781 205650 52123
rect 207243 52052 207309 52053
rect 207243 51988 207244 52052
rect 207308 51988 207309 52052
rect 207243 51987 207309 51988
rect 205771 51950 205837 51951
rect 205771 51886 205772 51950
rect 205836 51914 205837 51950
rect 206323 51916 206389 51917
rect 206323 51914 206324 51916
rect 205836 51886 206018 51914
rect 205771 51885 206018 51886
rect 205774 51854 206018 51885
rect 205587 51780 205653 51781
rect 205587 51716 205588 51780
rect 205652 51716 205653 51780
rect 205587 51715 205653 51716
rect 205403 50148 205469 50149
rect 205403 50084 205404 50148
rect 205468 50084 205469 50148
rect 205403 50083 205469 50084
rect 205219 19956 205285 19957
rect 205219 19892 205220 19956
rect 205284 19892 205285 19956
rect 205219 19891 205285 19892
rect 205406 9077 205466 50083
rect 205958 50013 206018 51854
rect 206142 51854 206324 51914
rect 205955 50012 206021 50013
rect 205955 49948 205956 50012
rect 206020 49948 206021 50012
rect 205955 49947 206021 49948
rect 206142 48381 206202 51854
rect 206323 51852 206324 51854
rect 206388 51852 206389 51916
rect 206323 51851 206389 51852
rect 206691 51916 206757 51917
rect 206691 51852 206692 51916
rect 206756 51852 206757 51916
rect 207059 51916 207125 51917
rect 207059 51914 207060 51916
rect 206691 51851 206757 51852
rect 206878 51854 207060 51914
rect 206507 51780 206573 51781
rect 206507 51778 206508 51780
rect 206326 51718 206508 51778
rect 206139 48380 206205 48381
rect 206139 48316 206140 48380
rect 206204 48316 206205 48380
rect 206139 48315 206205 48316
rect 205403 9076 205469 9077
rect 205403 9012 205404 9076
rect 205468 9012 205469 9076
rect 205403 9011 205469 9012
rect 206326 3365 206386 51718
rect 206507 51716 206508 51718
rect 206572 51716 206573 51780
rect 206507 51715 206573 51716
rect 206507 50148 206573 50149
rect 206507 50084 206508 50148
rect 206572 50084 206573 50148
rect 206507 50083 206573 50084
rect 206510 17509 206570 50083
rect 206507 17508 206573 17509
rect 206507 17444 206508 17508
rect 206572 17444 206573 17508
rect 206507 17443 206573 17444
rect 206694 12069 206754 51851
rect 206878 49741 206938 51854
rect 207059 51852 207060 51854
rect 207124 51852 207125 51916
rect 207059 51851 207125 51852
rect 207059 50148 207125 50149
rect 207059 50084 207060 50148
rect 207124 50084 207125 50148
rect 207059 50083 207125 50084
rect 206875 49740 206941 49741
rect 206875 49676 206876 49740
rect 206940 49676 206941 49740
rect 206875 49675 206941 49676
rect 207062 48330 207122 50083
rect 206878 48270 207122 48330
rect 206878 46205 206938 48270
rect 206875 46204 206941 46205
rect 206875 46140 206876 46204
rect 206940 46140 206941 46204
rect 206875 46139 206941 46140
rect 207246 17373 207306 51987
rect 207427 51916 207493 51917
rect 207427 51852 207428 51916
rect 207492 51852 207493 51916
rect 207427 51851 207493 51852
rect 207430 50010 207490 51851
rect 207611 51780 207677 51781
rect 207611 51716 207612 51780
rect 207676 51716 207677 51780
rect 207611 51715 207677 51716
rect 207614 50149 207674 51715
rect 207611 50148 207677 50149
rect 207611 50084 207612 50148
rect 207676 50084 207677 50148
rect 207611 50083 207677 50084
rect 207430 49950 207674 50010
rect 207427 49876 207493 49877
rect 207427 49812 207428 49876
rect 207492 49812 207493 49876
rect 207427 49811 207493 49812
rect 207243 17372 207309 17373
rect 207243 17308 207244 17372
rect 207308 17308 207309 17372
rect 207243 17307 207309 17308
rect 206691 12068 206757 12069
rect 206691 12004 206692 12068
rect 206756 12004 206757 12068
rect 206691 12003 206757 12004
rect 207430 6221 207490 49811
rect 207614 47565 207674 49950
rect 207611 47564 207677 47565
rect 207611 47500 207612 47564
rect 207676 47500 207677 47564
rect 207611 47499 207677 47500
rect 207834 29494 208454 52068
rect 209083 52052 209149 52053
rect 209083 51988 209084 52052
rect 209148 51988 209149 52052
rect 209083 51987 209149 51988
rect 209086 35325 209146 51987
rect 209267 51916 209333 51917
rect 209267 51852 209268 51916
rect 209332 51852 209333 51916
rect 209267 51851 209333 51852
rect 209451 51916 209517 51917
rect 209451 51852 209452 51916
rect 209516 51852 209517 51916
rect 209451 51851 209517 51852
rect 210555 51916 210621 51917
rect 210555 51852 210556 51916
rect 210620 51914 210621 51916
rect 210923 51916 210989 51917
rect 210620 51854 210802 51914
rect 210620 51852 210621 51854
rect 210555 51851 210621 51852
rect 209270 50149 209330 51851
rect 209267 50148 209333 50149
rect 209267 50084 209268 50148
rect 209332 50084 209333 50148
rect 209267 50083 209333 50084
rect 209267 50012 209333 50013
rect 209267 49948 209268 50012
rect 209332 49948 209333 50012
rect 209267 49947 209333 49948
rect 209083 35324 209149 35325
rect 209083 35260 209084 35324
rect 209148 35260 209149 35324
rect 209083 35259 209149 35260
rect 207834 29258 207866 29494
rect 208102 29258 208186 29494
rect 208422 29258 208454 29494
rect 207834 29174 208454 29258
rect 207834 28938 207866 29174
rect 208102 28938 208186 29174
rect 208422 28938 208454 29174
rect 207427 6220 207493 6221
rect 207427 6156 207428 6220
rect 207492 6156 207493 6220
rect 207427 6155 207493 6156
rect 206323 3364 206389 3365
rect 206323 3300 206324 3364
rect 206388 3300 206389 3364
rect 206323 3299 206389 3300
rect 204114 -6342 204146 -6106
rect 204382 -6342 204466 -6106
rect 204702 -6342 204734 -6106
rect 204114 -6426 204734 -6342
rect 204114 -6662 204146 -6426
rect 204382 -6662 204466 -6426
rect 204702 -6662 204734 -6426
rect 204114 -7654 204734 -6662
rect 207834 -7066 208454 28938
rect 209270 26893 209330 49947
rect 209267 26892 209333 26893
rect 209267 26828 209268 26892
rect 209332 26828 209333 26892
rect 209267 26827 209333 26828
rect 209454 24309 209514 51851
rect 210187 51780 210253 51781
rect 210187 51716 210188 51780
rect 210252 51716 210253 51780
rect 210187 51715 210253 51716
rect 210555 51780 210621 51781
rect 210555 51716 210556 51780
rect 210620 51716 210621 51780
rect 210555 51715 210621 51716
rect 209635 50148 209701 50149
rect 209635 50084 209636 50148
rect 209700 50084 209701 50148
rect 209635 50083 209701 50084
rect 209451 24308 209517 24309
rect 209451 24244 209452 24308
rect 209516 24244 209517 24308
rect 209451 24243 209517 24244
rect 209638 10301 209698 50083
rect 210190 48789 210250 51715
rect 210371 50148 210437 50149
rect 210371 50084 210372 50148
rect 210436 50084 210437 50148
rect 210371 50083 210437 50084
rect 210187 48788 210253 48789
rect 210187 48724 210188 48788
rect 210252 48724 210253 48788
rect 210187 48723 210253 48724
rect 210374 33965 210434 50083
rect 210371 33964 210437 33965
rect 210371 33900 210372 33964
rect 210436 33900 210437 33964
rect 210371 33899 210437 33900
rect 210558 28253 210618 51715
rect 210742 49741 210802 51854
rect 210923 51852 210924 51916
rect 210988 51852 210989 51916
rect 210923 51851 210989 51852
rect 212027 51916 212093 51917
rect 212027 51852 212028 51916
rect 212092 51852 212093 51916
rect 213499 51916 213565 51917
rect 213499 51914 213500 51916
rect 212027 51851 212093 51852
rect 213318 51854 213500 51914
rect 210739 49740 210805 49741
rect 210739 49676 210740 49740
rect 210804 49676 210805 49740
rect 210739 49675 210805 49676
rect 210739 48788 210805 48789
rect 210739 48724 210740 48788
rect 210804 48724 210805 48788
rect 210739 48723 210805 48724
rect 210742 28389 210802 48723
rect 210739 28388 210805 28389
rect 210739 28324 210740 28388
rect 210804 28324 210805 28388
rect 210739 28323 210805 28324
rect 210555 28252 210621 28253
rect 210555 28188 210556 28252
rect 210620 28188 210621 28252
rect 210555 28187 210621 28188
rect 210926 17237 210986 51851
rect 211659 51780 211725 51781
rect 211659 51716 211660 51780
rect 211724 51716 211725 51780
rect 211659 51715 211725 51716
rect 211662 45797 211722 51715
rect 211843 48788 211909 48789
rect 211843 48724 211844 48788
rect 211908 48724 211909 48788
rect 211843 48723 211909 48724
rect 211659 45796 211725 45797
rect 211659 45732 211660 45796
rect 211724 45732 211725 45796
rect 211659 45731 211725 45732
rect 211846 33829 211906 48723
rect 211843 33828 211909 33829
rect 211843 33764 211844 33828
rect 211908 33764 211909 33828
rect 211843 33763 211909 33764
rect 212030 30973 212090 51851
rect 212211 51780 212277 51781
rect 212211 51716 212212 51780
rect 212276 51716 212277 51780
rect 212211 51715 212277 51716
rect 212395 51780 212461 51781
rect 212395 51716 212396 51780
rect 212460 51716 212461 51780
rect 212395 51715 212461 51716
rect 212027 30972 212093 30973
rect 212027 30908 212028 30972
rect 212092 30908 212093 30972
rect 212027 30907 212093 30908
rect 210923 17236 210989 17237
rect 210923 17172 210924 17236
rect 210988 17172 210989 17236
rect 210923 17171 210989 17172
rect 212214 11933 212274 51715
rect 212211 11932 212277 11933
rect 212211 11868 212212 11932
rect 212276 11868 212277 11932
rect 212211 11867 212277 11868
rect 212398 11797 212458 51715
rect 213131 48924 213197 48925
rect 213131 48860 213132 48924
rect 213196 48860 213197 48924
rect 213131 48859 213197 48860
rect 213134 35189 213194 48859
rect 213131 35188 213197 35189
rect 213131 35124 213132 35188
rect 213196 35124 213197 35188
rect 213131 35123 213197 35124
rect 213318 32469 213378 51854
rect 213499 51852 213500 51854
rect 213564 51852 213565 51916
rect 213499 51851 213565 51852
rect 214051 51916 214117 51917
rect 214051 51852 214052 51916
rect 214116 51852 214117 51916
rect 214051 51851 214117 51852
rect 215523 51916 215589 51917
rect 215523 51852 215524 51916
rect 215588 51852 215589 51916
rect 215523 51851 215589 51852
rect 213499 50012 213565 50013
rect 213499 49948 213500 50012
rect 213564 49948 213565 50012
rect 213499 49947 213565 49948
rect 213502 32605 213562 49947
rect 213683 49740 213749 49741
rect 213683 49676 213684 49740
rect 213748 49676 213749 49740
rect 213683 49675 213749 49676
rect 213499 32604 213565 32605
rect 213499 32540 213500 32604
rect 213564 32540 213565 32604
rect 213499 32539 213565 32540
rect 213315 32468 213381 32469
rect 213315 32404 213316 32468
rect 213380 32404 213381 32468
rect 213315 32403 213381 32404
rect 212395 11796 212461 11797
rect 212395 11732 212396 11796
rect 212460 11732 212461 11796
rect 212395 11731 212461 11732
rect 209635 10300 209701 10301
rect 209635 10236 209636 10300
rect 209700 10236 209701 10300
rect 209635 10235 209701 10236
rect 213686 8941 213746 49675
rect 214054 47973 214114 51851
rect 214235 51780 214301 51781
rect 214235 51716 214236 51780
rect 214300 51716 214301 51780
rect 214235 51715 214301 51716
rect 214238 48381 214298 51715
rect 215155 49060 215221 49061
rect 215155 48996 215156 49060
rect 215220 48996 215221 49060
rect 215155 48995 215221 48996
rect 214419 48924 214485 48925
rect 214419 48860 214420 48924
rect 214484 48860 214485 48924
rect 214419 48859 214485 48860
rect 214235 48380 214301 48381
rect 214235 48316 214236 48380
rect 214300 48316 214301 48380
rect 214235 48315 214301 48316
rect 214051 47972 214117 47973
rect 214051 47908 214052 47972
rect 214116 47908 214117 47972
rect 214051 47907 214117 47908
rect 213683 8940 213749 8941
rect 213683 8876 213684 8940
rect 213748 8876 213749 8940
rect 213683 8875 213749 8876
rect 214422 4861 214482 48859
rect 214787 48788 214853 48789
rect 214787 48724 214788 48788
rect 214852 48724 214853 48788
rect 214787 48723 214853 48724
rect 214603 48380 214669 48381
rect 214603 48316 214604 48380
rect 214668 48316 214669 48380
rect 214603 48315 214669 48316
rect 214606 25669 214666 48315
rect 214603 25668 214669 25669
rect 214603 25604 214604 25668
rect 214668 25604 214669 25668
rect 214603 25603 214669 25604
rect 214790 24173 214850 48723
rect 215158 48381 215218 48995
rect 215526 48789 215586 51851
rect 215523 48788 215589 48789
rect 215523 48724 215524 48788
rect 215588 48724 215589 48788
rect 215523 48723 215589 48724
rect 215155 48380 215221 48381
rect 215155 48316 215156 48380
rect 215220 48316 215221 48380
rect 215155 48315 215221 48316
rect 214971 47972 215037 47973
rect 214971 47908 214972 47972
rect 215036 47908 215037 47972
rect 214971 47907 215037 47908
rect 214787 24172 214853 24173
rect 214787 24108 214788 24172
rect 214852 24108 214853 24172
rect 214787 24107 214853 24108
rect 214974 11661 215034 47907
rect 217794 39454 218414 74898
rect 217794 39218 217826 39454
rect 218062 39218 218146 39454
rect 218382 39218 218414 39454
rect 217794 39134 218414 39218
rect 217794 38898 217826 39134
rect 218062 38898 218146 39134
rect 218382 38898 218414 39134
rect 214971 11660 215037 11661
rect 214971 11596 214972 11660
rect 215036 11596 215037 11660
rect 214971 11595 215037 11596
rect 214419 4860 214485 4861
rect 214419 4796 214420 4860
rect 214484 4796 214485 4860
rect 214419 4795 214485 4796
rect 207834 -7302 207866 -7066
rect 208102 -7302 208186 -7066
rect 208422 -7302 208454 -7066
rect 207834 -7386 208454 -7302
rect 207834 -7622 207866 -7386
rect 208102 -7622 208186 -7386
rect 208422 -7622 208454 -7386
rect 207834 -7654 208454 -7622
rect 217794 3454 218414 38898
rect 217794 3218 217826 3454
rect 218062 3218 218146 3454
rect 218382 3218 218414 3454
rect 217794 3134 218414 3218
rect 217794 2898 217826 3134
rect 218062 2898 218146 3134
rect 218382 2898 218414 3134
rect 217794 -346 218414 2898
rect 217794 -582 217826 -346
rect 218062 -582 218146 -346
rect 218382 -582 218414 -346
rect 217794 -666 218414 -582
rect 217794 -902 217826 -666
rect 218062 -902 218146 -666
rect 218382 -902 218414 -666
rect 217794 -7654 218414 -902
rect 221514 705798 222134 711590
rect 221514 705562 221546 705798
rect 221782 705562 221866 705798
rect 222102 705562 222134 705798
rect 221514 705478 222134 705562
rect 221514 705242 221546 705478
rect 221782 705242 221866 705478
rect 222102 705242 222134 705478
rect 221514 691174 222134 705242
rect 221514 690938 221546 691174
rect 221782 690938 221866 691174
rect 222102 690938 222134 691174
rect 221514 690854 222134 690938
rect 221514 690618 221546 690854
rect 221782 690618 221866 690854
rect 222102 690618 222134 690854
rect 221514 655174 222134 690618
rect 221514 654938 221546 655174
rect 221782 654938 221866 655174
rect 222102 654938 222134 655174
rect 221514 654854 222134 654938
rect 221514 654618 221546 654854
rect 221782 654618 221866 654854
rect 222102 654618 222134 654854
rect 221514 619174 222134 654618
rect 221514 618938 221546 619174
rect 221782 618938 221866 619174
rect 222102 618938 222134 619174
rect 221514 618854 222134 618938
rect 221514 618618 221546 618854
rect 221782 618618 221866 618854
rect 222102 618618 222134 618854
rect 221514 583174 222134 618618
rect 221514 582938 221546 583174
rect 221782 582938 221866 583174
rect 222102 582938 222134 583174
rect 221514 582854 222134 582938
rect 221514 582618 221546 582854
rect 221782 582618 221866 582854
rect 222102 582618 222134 582854
rect 221514 547174 222134 582618
rect 221514 546938 221546 547174
rect 221782 546938 221866 547174
rect 222102 546938 222134 547174
rect 221514 546854 222134 546938
rect 221514 546618 221546 546854
rect 221782 546618 221866 546854
rect 222102 546618 222134 546854
rect 221514 511174 222134 546618
rect 221514 510938 221546 511174
rect 221782 510938 221866 511174
rect 222102 510938 222134 511174
rect 221514 510854 222134 510938
rect 221514 510618 221546 510854
rect 221782 510618 221866 510854
rect 222102 510618 222134 510854
rect 221514 475174 222134 510618
rect 221514 474938 221546 475174
rect 221782 474938 221866 475174
rect 222102 474938 222134 475174
rect 221514 474854 222134 474938
rect 221514 474618 221546 474854
rect 221782 474618 221866 474854
rect 222102 474618 222134 474854
rect 221514 439174 222134 474618
rect 221514 438938 221546 439174
rect 221782 438938 221866 439174
rect 222102 438938 222134 439174
rect 221514 438854 222134 438938
rect 221514 438618 221546 438854
rect 221782 438618 221866 438854
rect 222102 438618 222134 438854
rect 221514 403174 222134 438618
rect 221514 402938 221546 403174
rect 221782 402938 221866 403174
rect 222102 402938 222134 403174
rect 221514 402854 222134 402938
rect 221514 402618 221546 402854
rect 221782 402618 221866 402854
rect 222102 402618 222134 402854
rect 221514 367174 222134 402618
rect 221514 366938 221546 367174
rect 221782 366938 221866 367174
rect 222102 366938 222134 367174
rect 221514 366854 222134 366938
rect 221514 366618 221546 366854
rect 221782 366618 221866 366854
rect 222102 366618 222134 366854
rect 221514 331174 222134 366618
rect 221514 330938 221546 331174
rect 221782 330938 221866 331174
rect 222102 330938 222134 331174
rect 221514 330854 222134 330938
rect 221514 330618 221546 330854
rect 221782 330618 221866 330854
rect 222102 330618 222134 330854
rect 221514 295174 222134 330618
rect 225234 706758 225854 711590
rect 225234 706522 225266 706758
rect 225502 706522 225586 706758
rect 225822 706522 225854 706758
rect 225234 706438 225854 706522
rect 225234 706202 225266 706438
rect 225502 706202 225586 706438
rect 225822 706202 225854 706438
rect 225234 694894 225854 706202
rect 225234 694658 225266 694894
rect 225502 694658 225586 694894
rect 225822 694658 225854 694894
rect 225234 694574 225854 694658
rect 225234 694338 225266 694574
rect 225502 694338 225586 694574
rect 225822 694338 225854 694574
rect 225234 658894 225854 694338
rect 225234 658658 225266 658894
rect 225502 658658 225586 658894
rect 225822 658658 225854 658894
rect 225234 658574 225854 658658
rect 225234 658338 225266 658574
rect 225502 658338 225586 658574
rect 225822 658338 225854 658574
rect 225234 622894 225854 658338
rect 225234 622658 225266 622894
rect 225502 622658 225586 622894
rect 225822 622658 225854 622894
rect 225234 622574 225854 622658
rect 225234 622338 225266 622574
rect 225502 622338 225586 622574
rect 225822 622338 225854 622574
rect 225234 586894 225854 622338
rect 225234 586658 225266 586894
rect 225502 586658 225586 586894
rect 225822 586658 225854 586894
rect 225234 586574 225854 586658
rect 225234 586338 225266 586574
rect 225502 586338 225586 586574
rect 225822 586338 225854 586574
rect 225234 550894 225854 586338
rect 225234 550658 225266 550894
rect 225502 550658 225586 550894
rect 225822 550658 225854 550894
rect 225234 550574 225854 550658
rect 225234 550338 225266 550574
rect 225502 550338 225586 550574
rect 225822 550338 225854 550574
rect 225234 514894 225854 550338
rect 225234 514658 225266 514894
rect 225502 514658 225586 514894
rect 225822 514658 225854 514894
rect 225234 514574 225854 514658
rect 225234 514338 225266 514574
rect 225502 514338 225586 514574
rect 225822 514338 225854 514574
rect 225234 478894 225854 514338
rect 225234 478658 225266 478894
rect 225502 478658 225586 478894
rect 225822 478658 225854 478894
rect 225234 478574 225854 478658
rect 225234 478338 225266 478574
rect 225502 478338 225586 478574
rect 225822 478338 225854 478574
rect 225234 442894 225854 478338
rect 225234 442658 225266 442894
rect 225502 442658 225586 442894
rect 225822 442658 225854 442894
rect 225234 442574 225854 442658
rect 225234 442338 225266 442574
rect 225502 442338 225586 442574
rect 225822 442338 225854 442574
rect 225234 406894 225854 442338
rect 225234 406658 225266 406894
rect 225502 406658 225586 406894
rect 225822 406658 225854 406894
rect 225234 406574 225854 406658
rect 225234 406338 225266 406574
rect 225502 406338 225586 406574
rect 225822 406338 225854 406574
rect 225234 370894 225854 406338
rect 225234 370658 225266 370894
rect 225502 370658 225586 370894
rect 225822 370658 225854 370894
rect 225234 370574 225854 370658
rect 225234 370338 225266 370574
rect 225502 370338 225586 370574
rect 225822 370338 225854 370574
rect 225234 334894 225854 370338
rect 225234 334658 225266 334894
rect 225502 334658 225586 334894
rect 225822 334658 225854 334894
rect 225234 334574 225854 334658
rect 225234 334338 225266 334574
rect 225502 334338 225586 334574
rect 225822 334338 225854 334574
rect 224171 300388 224237 300389
rect 224171 300324 224172 300388
rect 224236 300324 224237 300388
rect 224171 300323 224237 300324
rect 221514 294938 221546 295174
rect 221782 294938 221866 295174
rect 222102 294938 222134 295174
rect 221514 294854 222134 294938
rect 221514 294618 221546 294854
rect 221782 294618 221866 294854
rect 222102 294618 222134 294854
rect 221514 259174 222134 294618
rect 221514 258938 221546 259174
rect 221782 258938 221866 259174
rect 222102 258938 222134 259174
rect 221514 258854 222134 258938
rect 221514 258618 221546 258854
rect 221782 258618 221866 258854
rect 222102 258618 222134 258854
rect 221514 223174 222134 258618
rect 221514 222938 221546 223174
rect 221782 222938 221866 223174
rect 222102 222938 222134 223174
rect 221514 222854 222134 222938
rect 221514 222618 221546 222854
rect 221782 222618 221866 222854
rect 222102 222618 222134 222854
rect 221514 187174 222134 222618
rect 221514 186938 221546 187174
rect 221782 186938 221866 187174
rect 222102 186938 222134 187174
rect 221514 186854 222134 186938
rect 221514 186618 221546 186854
rect 221782 186618 221866 186854
rect 222102 186618 222134 186854
rect 221514 151174 222134 186618
rect 221514 150938 221546 151174
rect 221782 150938 221866 151174
rect 222102 150938 222134 151174
rect 221514 150854 222134 150938
rect 221514 150618 221546 150854
rect 221782 150618 221866 150854
rect 222102 150618 222134 150854
rect 221514 115174 222134 150618
rect 224174 122909 224234 300323
rect 225234 298894 225854 334338
rect 225234 298658 225266 298894
rect 225502 298658 225586 298894
rect 225822 298658 225854 298894
rect 225234 298574 225854 298658
rect 225234 298338 225266 298574
rect 225502 298338 225586 298574
rect 225822 298338 225854 298574
rect 225234 262894 225854 298338
rect 225234 262658 225266 262894
rect 225502 262658 225586 262894
rect 225822 262658 225854 262894
rect 225234 262574 225854 262658
rect 225234 262338 225266 262574
rect 225502 262338 225586 262574
rect 225822 262338 225854 262574
rect 225234 226894 225854 262338
rect 225234 226658 225266 226894
rect 225502 226658 225586 226894
rect 225822 226658 225854 226894
rect 225234 226574 225854 226658
rect 225234 226338 225266 226574
rect 225502 226338 225586 226574
rect 225822 226338 225854 226574
rect 225234 190894 225854 226338
rect 225234 190658 225266 190894
rect 225502 190658 225586 190894
rect 225822 190658 225854 190894
rect 225234 190574 225854 190658
rect 225234 190338 225266 190574
rect 225502 190338 225586 190574
rect 225822 190338 225854 190574
rect 225234 154894 225854 190338
rect 225234 154658 225266 154894
rect 225502 154658 225586 154894
rect 225822 154658 225854 154894
rect 225234 154574 225854 154658
rect 225234 154338 225266 154574
rect 225502 154338 225586 154574
rect 225822 154338 225854 154574
rect 224171 122908 224237 122909
rect 224171 122844 224172 122908
rect 224236 122844 224237 122908
rect 224171 122843 224237 122844
rect 221514 114938 221546 115174
rect 221782 114938 221866 115174
rect 222102 114938 222134 115174
rect 221514 114854 222134 114938
rect 221514 114618 221546 114854
rect 221782 114618 221866 114854
rect 222102 114618 222134 114854
rect 221514 79174 222134 114618
rect 221514 78938 221546 79174
rect 221782 78938 221866 79174
rect 222102 78938 222134 79174
rect 221514 78854 222134 78938
rect 221514 78618 221546 78854
rect 221782 78618 221866 78854
rect 222102 78618 222134 78854
rect 221514 43174 222134 78618
rect 221514 42938 221546 43174
rect 221782 42938 221866 43174
rect 222102 42938 222134 43174
rect 221514 42854 222134 42938
rect 221514 42618 221546 42854
rect 221782 42618 221866 42854
rect 222102 42618 222134 42854
rect 221514 7174 222134 42618
rect 221514 6938 221546 7174
rect 221782 6938 221866 7174
rect 222102 6938 222134 7174
rect 221514 6854 222134 6938
rect 221514 6618 221546 6854
rect 221782 6618 221866 6854
rect 222102 6618 222134 6854
rect 221514 -1306 222134 6618
rect 221514 -1542 221546 -1306
rect 221782 -1542 221866 -1306
rect 222102 -1542 222134 -1306
rect 221514 -1626 222134 -1542
rect 221514 -1862 221546 -1626
rect 221782 -1862 221866 -1626
rect 222102 -1862 222134 -1626
rect 221514 -7654 222134 -1862
rect 225234 118894 225854 154338
rect 225234 118658 225266 118894
rect 225502 118658 225586 118894
rect 225822 118658 225854 118894
rect 225234 118574 225854 118658
rect 225234 118338 225266 118574
rect 225502 118338 225586 118574
rect 225822 118338 225854 118574
rect 225234 82894 225854 118338
rect 225234 82658 225266 82894
rect 225502 82658 225586 82894
rect 225822 82658 225854 82894
rect 225234 82574 225854 82658
rect 225234 82338 225266 82574
rect 225502 82338 225586 82574
rect 225822 82338 225854 82574
rect 225234 46894 225854 82338
rect 225234 46658 225266 46894
rect 225502 46658 225586 46894
rect 225822 46658 225854 46894
rect 225234 46574 225854 46658
rect 225234 46338 225266 46574
rect 225502 46338 225586 46574
rect 225822 46338 225854 46574
rect 225234 10894 225854 46338
rect 225234 10658 225266 10894
rect 225502 10658 225586 10894
rect 225822 10658 225854 10894
rect 225234 10574 225854 10658
rect 225234 10338 225266 10574
rect 225502 10338 225586 10574
rect 225822 10338 225854 10574
rect 225234 -2266 225854 10338
rect 225234 -2502 225266 -2266
rect 225502 -2502 225586 -2266
rect 225822 -2502 225854 -2266
rect 225234 -2586 225854 -2502
rect 225234 -2822 225266 -2586
rect 225502 -2822 225586 -2586
rect 225822 -2822 225854 -2586
rect 225234 -7654 225854 -2822
rect 228954 707718 229574 711590
rect 228954 707482 228986 707718
rect 229222 707482 229306 707718
rect 229542 707482 229574 707718
rect 228954 707398 229574 707482
rect 228954 707162 228986 707398
rect 229222 707162 229306 707398
rect 229542 707162 229574 707398
rect 228954 698614 229574 707162
rect 228954 698378 228986 698614
rect 229222 698378 229306 698614
rect 229542 698378 229574 698614
rect 228954 698294 229574 698378
rect 228954 698058 228986 698294
rect 229222 698058 229306 698294
rect 229542 698058 229574 698294
rect 228954 662614 229574 698058
rect 228954 662378 228986 662614
rect 229222 662378 229306 662614
rect 229542 662378 229574 662614
rect 228954 662294 229574 662378
rect 228954 662058 228986 662294
rect 229222 662058 229306 662294
rect 229542 662058 229574 662294
rect 228954 626614 229574 662058
rect 228954 626378 228986 626614
rect 229222 626378 229306 626614
rect 229542 626378 229574 626614
rect 228954 626294 229574 626378
rect 228954 626058 228986 626294
rect 229222 626058 229306 626294
rect 229542 626058 229574 626294
rect 228954 590614 229574 626058
rect 228954 590378 228986 590614
rect 229222 590378 229306 590614
rect 229542 590378 229574 590614
rect 228954 590294 229574 590378
rect 228954 590058 228986 590294
rect 229222 590058 229306 590294
rect 229542 590058 229574 590294
rect 228954 554614 229574 590058
rect 228954 554378 228986 554614
rect 229222 554378 229306 554614
rect 229542 554378 229574 554614
rect 228954 554294 229574 554378
rect 228954 554058 228986 554294
rect 229222 554058 229306 554294
rect 229542 554058 229574 554294
rect 228954 518614 229574 554058
rect 228954 518378 228986 518614
rect 229222 518378 229306 518614
rect 229542 518378 229574 518614
rect 228954 518294 229574 518378
rect 228954 518058 228986 518294
rect 229222 518058 229306 518294
rect 229542 518058 229574 518294
rect 228954 482614 229574 518058
rect 228954 482378 228986 482614
rect 229222 482378 229306 482614
rect 229542 482378 229574 482614
rect 228954 482294 229574 482378
rect 228954 482058 228986 482294
rect 229222 482058 229306 482294
rect 229542 482058 229574 482294
rect 228954 446614 229574 482058
rect 228954 446378 228986 446614
rect 229222 446378 229306 446614
rect 229542 446378 229574 446614
rect 228954 446294 229574 446378
rect 228954 446058 228986 446294
rect 229222 446058 229306 446294
rect 229542 446058 229574 446294
rect 228954 410614 229574 446058
rect 228954 410378 228986 410614
rect 229222 410378 229306 410614
rect 229542 410378 229574 410614
rect 228954 410294 229574 410378
rect 228954 410058 228986 410294
rect 229222 410058 229306 410294
rect 229542 410058 229574 410294
rect 228954 374614 229574 410058
rect 228954 374378 228986 374614
rect 229222 374378 229306 374614
rect 229542 374378 229574 374614
rect 228954 374294 229574 374378
rect 228954 374058 228986 374294
rect 229222 374058 229306 374294
rect 229542 374058 229574 374294
rect 228954 338614 229574 374058
rect 228954 338378 228986 338614
rect 229222 338378 229306 338614
rect 229542 338378 229574 338614
rect 228954 338294 229574 338378
rect 228954 338058 228986 338294
rect 229222 338058 229306 338294
rect 229542 338058 229574 338294
rect 228954 302614 229574 338058
rect 228954 302378 228986 302614
rect 229222 302378 229306 302614
rect 229542 302378 229574 302614
rect 228954 302294 229574 302378
rect 228954 302058 228986 302294
rect 229222 302058 229306 302294
rect 229542 302058 229574 302294
rect 228954 266614 229574 302058
rect 228954 266378 228986 266614
rect 229222 266378 229306 266614
rect 229542 266378 229574 266614
rect 228954 266294 229574 266378
rect 228954 266058 228986 266294
rect 229222 266058 229306 266294
rect 229542 266058 229574 266294
rect 228954 230614 229574 266058
rect 228954 230378 228986 230614
rect 229222 230378 229306 230614
rect 229542 230378 229574 230614
rect 228954 230294 229574 230378
rect 228954 230058 228986 230294
rect 229222 230058 229306 230294
rect 229542 230058 229574 230294
rect 228954 194614 229574 230058
rect 228954 194378 228986 194614
rect 229222 194378 229306 194614
rect 229542 194378 229574 194614
rect 228954 194294 229574 194378
rect 228954 194058 228986 194294
rect 229222 194058 229306 194294
rect 229542 194058 229574 194294
rect 228954 158614 229574 194058
rect 228954 158378 228986 158614
rect 229222 158378 229306 158614
rect 229542 158378 229574 158614
rect 228954 158294 229574 158378
rect 228954 158058 228986 158294
rect 229222 158058 229306 158294
rect 229542 158058 229574 158294
rect 228954 122614 229574 158058
rect 228954 122378 228986 122614
rect 229222 122378 229306 122614
rect 229542 122378 229574 122614
rect 228954 122294 229574 122378
rect 228954 122058 228986 122294
rect 229222 122058 229306 122294
rect 229542 122058 229574 122294
rect 228954 86614 229574 122058
rect 228954 86378 228986 86614
rect 229222 86378 229306 86614
rect 229542 86378 229574 86614
rect 228954 86294 229574 86378
rect 228954 86058 228986 86294
rect 229222 86058 229306 86294
rect 229542 86058 229574 86294
rect 228954 50614 229574 86058
rect 228954 50378 228986 50614
rect 229222 50378 229306 50614
rect 229542 50378 229574 50614
rect 228954 50294 229574 50378
rect 228954 50058 228986 50294
rect 229222 50058 229306 50294
rect 229542 50058 229574 50294
rect 228954 14614 229574 50058
rect 228954 14378 228986 14614
rect 229222 14378 229306 14614
rect 229542 14378 229574 14614
rect 228954 14294 229574 14378
rect 228954 14058 228986 14294
rect 229222 14058 229306 14294
rect 229542 14058 229574 14294
rect 228954 -3226 229574 14058
rect 228954 -3462 228986 -3226
rect 229222 -3462 229306 -3226
rect 229542 -3462 229574 -3226
rect 228954 -3546 229574 -3462
rect 228954 -3782 228986 -3546
rect 229222 -3782 229306 -3546
rect 229542 -3782 229574 -3546
rect 228954 -7654 229574 -3782
rect 232674 708678 233294 711590
rect 232674 708442 232706 708678
rect 232942 708442 233026 708678
rect 233262 708442 233294 708678
rect 232674 708358 233294 708442
rect 232674 708122 232706 708358
rect 232942 708122 233026 708358
rect 233262 708122 233294 708358
rect 232674 666334 233294 708122
rect 232674 666098 232706 666334
rect 232942 666098 233026 666334
rect 233262 666098 233294 666334
rect 232674 666014 233294 666098
rect 232674 665778 232706 666014
rect 232942 665778 233026 666014
rect 233262 665778 233294 666014
rect 232674 630334 233294 665778
rect 232674 630098 232706 630334
rect 232942 630098 233026 630334
rect 233262 630098 233294 630334
rect 232674 630014 233294 630098
rect 232674 629778 232706 630014
rect 232942 629778 233026 630014
rect 233262 629778 233294 630014
rect 232674 594334 233294 629778
rect 232674 594098 232706 594334
rect 232942 594098 233026 594334
rect 233262 594098 233294 594334
rect 232674 594014 233294 594098
rect 232674 593778 232706 594014
rect 232942 593778 233026 594014
rect 233262 593778 233294 594014
rect 232674 558334 233294 593778
rect 232674 558098 232706 558334
rect 232942 558098 233026 558334
rect 233262 558098 233294 558334
rect 232674 558014 233294 558098
rect 232674 557778 232706 558014
rect 232942 557778 233026 558014
rect 233262 557778 233294 558014
rect 232674 522334 233294 557778
rect 232674 522098 232706 522334
rect 232942 522098 233026 522334
rect 233262 522098 233294 522334
rect 232674 522014 233294 522098
rect 232674 521778 232706 522014
rect 232942 521778 233026 522014
rect 233262 521778 233294 522014
rect 232674 486334 233294 521778
rect 232674 486098 232706 486334
rect 232942 486098 233026 486334
rect 233262 486098 233294 486334
rect 232674 486014 233294 486098
rect 232674 485778 232706 486014
rect 232942 485778 233026 486014
rect 233262 485778 233294 486014
rect 232674 450334 233294 485778
rect 232674 450098 232706 450334
rect 232942 450098 233026 450334
rect 233262 450098 233294 450334
rect 232674 450014 233294 450098
rect 232674 449778 232706 450014
rect 232942 449778 233026 450014
rect 233262 449778 233294 450014
rect 232674 414334 233294 449778
rect 232674 414098 232706 414334
rect 232942 414098 233026 414334
rect 233262 414098 233294 414334
rect 232674 414014 233294 414098
rect 232674 413778 232706 414014
rect 232942 413778 233026 414014
rect 233262 413778 233294 414014
rect 232674 378334 233294 413778
rect 232674 378098 232706 378334
rect 232942 378098 233026 378334
rect 233262 378098 233294 378334
rect 232674 378014 233294 378098
rect 232674 377778 232706 378014
rect 232942 377778 233026 378014
rect 233262 377778 233294 378014
rect 232674 342334 233294 377778
rect 232674 342098 232706 342334
rect 232942 342098 233026 342334
rect 233262 342098 233294 342334
rect 232674 342014 233294 342098
rect 232674 341778 232706 342014
rect 232942 341778 233026 342014
rect 233262 341778 233294 342014
rect 232674 306334 233294 341778
rect 232674 306098 232706 306334
rect 232942 306098 233026 306334
rect 233262 306098 233294 306334
rect 232674 306014 233294 306098
rect 232674 305778 232706 306014
rect 232942 305778 233026 306014
rect 233262 305778 233294 306014
rect 232674 270334 233294 305778
rect 232674 270098 232706 270334
rect 232942 270098 233026 270334
rect 233262 270098 233294 270334
rect 232674 270014 233294 270098
rect 232674 269778 232706 270014
rect 232942 269778 233026 270014
rect 233262 269778 233294 270014
rect 232674 234334 233294 269778
rect 232674 234098 232706 234334
rect 232942 234098 233026 234334
rect 233262 234098 233294 234334
rect 232674 234014 233294 234098
rect 232674 233778 232706 234014
rect 232942 233778 233026 234014
rect 233262 233778 233294 234014
rect 232674 198334 233294 233778
rect 232674 198098 232706 198334
rect 232942 198098 233026 198334
rect 233262 198098 233294 198334
rect 232674 198014 233294 198098
rect 232674 197778 232706 198014
rect 232942 197778 233026 198014
rect 233262 197778 233294 198014
rect 232674 162334 233294 197778
rect 232674 162098 232706 162334
rect 232942 162098 233026 162334
rect 233262 162098 233294 162334
rect 232674 162014 233294 162098
rect 232674 161778 232706 162014
rect 232942 161778 233026 162014
rect 233262 161778 233294 162014
rect 232674 126334 233294 161778
rect 232674 126098 232706 126334
rect 232942 126098 233026 126334
rect 233262 126098 233294 126334
rect 232674 126014 233294 126098
rect 232674 125778 232706 126014
rect 232942 125778 233026 126014
rect 233262 125778 233294 126014
rect 232674 90334 233294 125778
rect 232674 90098 232706 90334
rect 232942 90098 233026 90334
rect 233262 90098 233294 90334
rect 232674 90014 233294 90098
rect 232674 89778 232706 90014
rect 232942 89778 233026 90014
rect 233262 89778 233294 90014
rect 232674 54334 233294 89778
rect 232674 54098 232706 54334
rect 232942 54098 233026 54334
rect 233262 54098 233294 54334
rect 232674 54014 233294 54098
rect 232674 53778 232706 54014
rect 232942 53778 233026 54014
rect 233262 53778 233294 54014
rect 232674 18334 233294 53778
rect 232674 18098 232706 18334
rect 232942 18098 233026 18334
rect 233262 18098 233294 18334
rect 232674 18014 233294 18098
rect 232674 17778 232706 18014
rect 232942 17778 233026 18014
rect 233262 17778 233294 18014
rect 232674 -4186 233294 17778
rect 232674 -4422 232706 -4186
rect 232942 -4422 233026 -4186
rect 233262 -4422 233294 -4186
rect 232674 -4506 233294 -4422
rect 232674 -4742 232706 -4506
rect 232942 -4742 233026 -4506
rect 233262 -4742 233294 -4506
rect 232674 -7654 233294 -4742
rect 236394 709638 237014 711590
rect 236394 709402 236426 709638
rect 236662 709402 236746 709638
rect 236982 709402 237014 709638
rect 236394 709318 237014 709402
rect 236394 709082 236426 709318
rect 236662 709082 236746 709318
rect 236982 709082 237014 709318
rect 236394 670054 237014 709082
rect 236394 669818 236426 670054
rect 236662 669818 236746 670054
rect 236982 669818 237014 670054
rect 236394 669734 237014 669818
rect 236394 669498 236426 669734
rect 236662 669498 236746 669734
rect 236982 669498 237014 669734
rect 236394 634054 237014 669498
rect 236394 633818 236426 634054
rect 236662 633818 236746 634054
rect 236982 633818 237014 634054
rect 236394 633734 237014 633818
rect 236394 633498 236426 633734
rect 236662 633498 236746 633734
rect 236982 633498 237014 633734
rect 236394 598054 237014 633498
rect 236394 597818 236426 598054
rect 236662 597818 236746 598054
rect 236982 597818 237014 598054
rect 236394 597734 237014 597818
rect 236394 597498 236426 597734
rect 236662 597498 236746 597734
rect 236982 597498 237014 597734
rect 236394 562054 237014 597498
rect 236394 561818 236426 562054
rect 236662 561818 236746 562054
rect 236982 561818 237014 562054
rect 236394 561734 237014 561818
rect 236394 561498 236426 561734
rect 236662 561498 236746 561734
rect 236982 561498 237014 561734
rect 236394 526054 237014 561498
rect 236394 525818 236426 526054
rect 236662 525818 236746 526054
rect 236982 525818 237014 526054
rect 236394 525734 237014 525818
rect 236394 525498 236426 525734
rect 236662 525498 236746 525734
rect 236982 525498 237014 525734
rect 236394 490054 237014 525498
rect 236394 489818 236426 490054
rect 236662 489818 236746 490054
rect 236982 489818 237014 490054
rect 236394 489734 237014 489818
rect 236394 489498 236426 489734
rect 236662 489498 236746 489734
rect 236982 489498 237014 489734
rect 236394 454054 237014 489498
rect 236394 453818 236426 454054
rect 236662 453818 236746 454054
rect 236982 453818 237014 454054
rect 236394 453734 237014 453818
rect 236394 453498 236426 453734
rect 236662 453498 236746 453734
rect 236982 453498 237014 453734
rect 236394 418054 237014 453498
rect 236394 417818 236426 418054
rect 236662 417818 236746 418054
rect 236982 417818 237014 418054
rect 236394 417734 237014 417818
rect 236394 417498 236426 417734
rect 236662 417498 236746 417734
rect 236982 417498 237014 417734
rect 236394 382054 237014 417498
rect 236394 381818 236426 382054
rect 236662 381818 236746 382054
rect 236982 381818 237014 382054
rect 236394 381734 237014 381818
rect 236394 381498 236426 381734
rect 236662 381498 236746 381734
rect 236982 381498 237014 381734
rect 236394 346054 237014 381498
rect 236394 345818 236426 346054
rect 236662 345818 236746 346054
rect 236982 345818 237014 346054
rect 236394 345734 237014 345818
rect 236394 345498 236426 345734
rect 236662 345498 236746 345734
rect 236982 345498 237014 345734
rect 236394 310054 237014 345498
rect 236394 309818 236426 310054
rect 236662 309818 236746 310054
rect 236982 309818 237014 310054
rect 236394 309734 237014 309818
rect 236394 309498 236426 309734
rect 236662 309498 236746 309734
rect 236982 309498 237014 309734
rect 236394 274054 237014 309498
rect 236394 273818 236426 274054
rect 236662 273818 236746 274054
rect 236982 273818 237014 274054
rect 236394 273734 237014 273818
rect 236394 273498 236426 273734
rect 236662 273498 236746 273734
rect 236982 273498 237014 273734
rect 236394 238054 237014 273498
rect 236394 237818 236426 238054
rect 236662 237818 236746 238054
rect 236982 237818 237014 238054
rect 236394 237734 237014 237818
rect 236394 237498 236426 237734
rect 236662 237498 236746 237734
rect 236982 237498 237014 237734
rect 236394 202054 237014 237498
rect 236394 201818 236426 202054
rect 236662 201818 236746 202054
rect 236982 201818 237014 202054
rect 236394 201734 237014 201818
rect 236394 201498 236426 201734
rect 236662 201498 236746 201734
rect 236982 201498 237014 201734
rect 236394 166054 237014 201498
rect 236394 165818 236426 166054
rect 236662 165818 236746 166054
rect 236982 165818 237014 166054
rect 236394 165734 237014 165818
rect 236394 165498 236426 165734
rect 236662 165498 236746 165734
rect 236982 165498 237014 165734
rect 236394 130054 237014 165498
rect 236394 129818 236426 130054
rect 236662 129818 236746 130054
rect 236982 129818 237014 130054
rect 236394 129734 237014 129818
rect 236394 129498 236426 129734
rect 236662 129498 236746 129734
rect 236982 129498 237014 129734
rect 236394 94054 237014 129498
rect 236394 93818 236426 94054
rect 236662 93818 236746 94054
rect 236982 93818 237014 94054
rect 236394 93734 237014 93818
rect 236394 93498 236426 93734
rect 236662 93498 236746 93734
rect 236982 93498 237014 93734
rect 236394 58054 237014 93498
rect 236394 57818 236426 58054
rect 236662 57818 236746 58054
rect 236982 57818 237014 58054
rect 236394 57734 237014 57818
rect 236394 57498 236426 57734
rect 236662 57498 236746 57734
rect 236982 57498 237014 57734
rect 236394 22054 237014 57498
rect 236394 21818 236426 22054
rect 236662 21818 236746 22054
rect 236982 21818 237014 22054
rect 236394 21734 237014 21818
rect 236394 21498 236426 21734
rect 236662 21498 236746 21734
rect 236982 21498 237014 21734
rect 236394 -5146 237014 21498
rect 236394 -5382 236426 -5146
rect 236662 -5382 236746 -5146
rect 236982 -5382 237014 -5146
rect 236394 -5466 237014 -5382
rect 236394 -5702 236426 -5466
rect 236662 -5702 236746 -5466
rect 236982 -5702 237014 -5466
rect 236394 -7654 237014 -5702
rect 240114 710598 240734 711590
rect 240114 710362 240146 710598
rect 240382 710362 240466 710598
rect 240702 710362 240734 710598
rect 240114 710278 240734 710362
rect 240114 710042 240146 710278
rect 240382 710042 240466 710278
rect 240702 710042 240734 710278
rect 240114 673774 240734 710042
rect 240114 673538 240146 673774
rect 240382 673538 240466 673774
rect 240702 673538 240734 673774
rect 240114 673454 240734 673538
rect 240114 673218 240146 673454
rect 240382 673218 240466 673454
rect 240702 673218 240734 673454
rect 240114 637774 240734 673218
rect 240114 637538 240146 637774
rect 240382 637538 240466 637774
rect 240702 637538 240734 637774
rect 240114 637454 240734 637538
rect 240114 637218 240146 637454
rect 240382 637218 240466 637454
rect 240702 637218 240734 637454
rect 240114 601774 240734 637218
rect 240114 601538 240146 601774
rect 240382 601538 240466 601774
rect 240702 601538 240734 601774
rect 240114 601454 240734 601538
rect 240114 601218 240146 601454
rect 240382 601218 240466 601454
rect 240702 601218 240734 601454
rect 240114 565774 240734 601218
rect 240114 565538 240146 565774
rect 240382 565538 240466 565774
rect 240702 565538 240734 565774
rect 240114 565454 240734 565538
rect 240114 565218 240146 565454
rect 240382 565218 240466 565454
rect 240702 565218 240734 565454
rect 240114 529774 240734 565218
rect 240114 529538 240146 529774
rect 240382 529538 240466 529774
rect 240702 529538 240734 529774
rect 240114 529454 240734 529538
rect 240114 529218 240146 529454
rect 240382 529218 240466 529454
rect 240702 529218 240734 529454
rect 240114 493774 240734 529218
rect 240114 493538 240146 493774
rect 240382 493538 240466 493774
rect 240702 493538 240734 493774
rect 240114 493454 240734 493538
rect 240114 493218 240146 493454
rect 240382 493218 240466 493454
rect 240702 493218 240734 493454
rect 240114 457774 240734 493218
rect 240114 457538 240146 457774
rect 240382 457538 240466 457774
rect 240702 457538 240734 457774
rect 240114 457454 240734 457538
rect 240114 457218 240146 457454
rect 240382 457218 240466 457454
rect 240702 457218 240734 457454
rect 240114 421774 240734 457218
rect 240114 421538 240146 421774
rect 240382 421538 240466 421774
rect 240702 421538 240734 421774
rect 240114 421454 240734 421538
rect 240114 421218 240146 421454
rect 240382 421218 240466 421454
rect 240702 421218 240734 421454
rect 240114 385774 240734 421218
rect 240114 385538 240146 385774
rect 240382 385538 240466 385774
rect 240702 385538 240734 385774
rect 240114 385454 240734 385538
rect 240114 385218 240146 385454
rect 240382 385218 240466 385454
rect 240702 385218 240734 385454
rect 240114 349774 240734 385218
rect 240114 349538 240146 349774
rect 240382 349538 240466 349774
rect 240702 349538 240734 349774
rect 240114 349454 240734 349538
rect 240114 349218 240146 349454
rect 240382 349218 240466 349454
rect 240702 349218 240734 349454
rect 240114 313774 240734 349218
rect 240114 313538 240146 313774
rect 240382 313538 240466 313774
rect 240702 313538 240734 313774
rect 240114 313454 240734 313538
rect 240114 313218 240146 313454
rect 240382 313218 240466 313454
rect 240702 313218 240734 313454
rect 240114 277774 240734 313218
rect 240114 277538 240146 277774
rect 240382 277538 240466 277774
rect 240702 277538 240734 277774
rect 240114 277454 240734 277538
rect 240114 277218 240146 277454
rect 240382 277218 240466 277454
rect 240702 277218 240734 277454
rect 240114 241774 240734 277218
rect 240114 241538 240146 241774
rect 240382 241538 240466 241774
rect 240702 241538 240734 241774
rect 240114 241454 240734 241538
rect 240114 241218 240146 241454
rect 240382 241218 240466 241454
rect 240702 241218 240734 241454
rect 240114 205774 240734 241218
rect 240114 205538 240146 205774
rect 240382 205538 240466 205774
rect 240702 205538 240734 205774
rect 240114 205454 240734 205538
rect 240114 205218 240146 205454
rect 240382 205218 240466 205454
rect 240702 205218 240734 205454
rect 240114 169774 240734 205218
rect 240114 169538 240146 169774
rect 240382 169538 240466 169774
rect 240702 169538 240734 169774
rect 240114 169454 240734 169538
rect 240114 169218 240146 169454
rect 240382 169218 240466 169454
rect 240702 169218 240734 169454
rect 240114 133774 240734 169218
rect 240114 133538 240146 133774
rect 240382 133538 240466 133774
rect 240702 133538 240734 133774
rect 240114 133454 240734 133538
rect 240114 133218 240146 133454
rect 240382 133218 240466 133454
rect 240702 133218 240734 133454
rect 240114 97774 240734 133218
rect 240114 97538 240146 97774
rect 240382 97538 240466 97774
rect 240702 97538 240734 97774
rect 240114 97454 240734 97538
rect 240114 97218 240146 97454
rect 240382 97218 240466 97454
rect 240702 97218 240734 97454
rect 240114 61774 240734 97218
rect 240114 61538 240146 61774
rect 240382 61538 240466 61774
rect 240702 61538 240734 61774
rect 240114 61454 240734 61538
rect 240114 61218 240146 61454
rect 240382 61218 240466 61454
rect 240702 61218 240734 61454
rect 240114 25774 240734 61218
rect 240114 25538 240146 25774
rect 240382 25538 240466 25774
rect 240702 25538 240734 25774
rect 240114 25454 240734 25538
rect 240114 25218 240146 25454
rect 240382 25218 240466 25454
rect 240702 25218 240734 25454
rect 240114 -6106 240734 25218
rect 240114 -6342 240146 -6106
rect 240382 -6342 240466 -6106
rect 240702 -6342 240734 -6106
rect 240114 -6426 240734 -6342
rect 240114 -6662 240146 -6426
rect 240382 -6662 240466 -6426
rect 240702 -6662 240734 -6426
rect 240114 -7654 240734 -6662
rect 243834 711558 244454 711590
rect 243834 711322 243866 711558
rect 244102 711322 244186 711558
rect 244422 711322 244454 711558
rect 243834 711238 244454 711322
rect 243834 711002 243866 711238
rect 244102 711002 244186 711238
rect 244422 711002 244454 711238
rect 243834 677494 244454 711002
rect 243834 677258 243866 677494
rect 244102 677258 244186 677494
rect 244422 677258 244454 677494
rect 243834 677174 244454 677258
rect 243834 676938 243866 677174
rect 244102 676938 244186 677174
rect 244422 676938 244454 677174
rect 243834 641494 244454 676938
rect 253794 704838 254414 711590
rect 253794 704602 253826 704838
rect 254062 704602 254146 704838
rect 254382 704602 254414 704838
rect 253794 704518 254414 704602
rect 253794 704282 253826 704518
rect 254062 704282 254146 704518
rect 254382 704282 254414 704518
rect 253794 687454 254414 704282
rect 253794 687218 253826 687454
rect 254062 687218 254146 687454
rect 254382 687218 254414 687454
rect 253794 687134 254414 687218
rect 253794 686898 253826 687134
rect 254062 686898 254146 687134
rect 254382 686898 254414 687134
rect 251771 670716 251837 670717
rect 251771 670652 251772 670716
rect 251836 670652 251837 670716
rect 251771 670651 251837 670652
rect 243834 641258 243866 641494
rect 244102 641258 244186 641494
rect 244422 641258 244454 641494
rect 243834 641174 244454 641258
rect 243834 640938 243866 641174
rect 244102 640938 244186 641174
rect 244422 640938 244454 641174
rect 243834 605494 244454 640938
rect 243834 605258 243866 605494
rect 244102 605258 244186 605494
rect 244422 605258 244454 605494
rect 243834 605174 244454 605258
rect 243834 604938 243866 605174
rect 244102 604938 244186 605174
rect 244422 604938 244454 605174
rect 243834 569494 244454 604938
rect 243834 569258 243866 569494
rect 244102 569258 244186 569494
rect 244422 569258 244454 569494
rect 243834 569174 244454 569258
rect 243834 568938 243866 569174
rect 244102 568938 244186 569174
rect 244422 568938 244454 569174
rect 243834 533494 244454 568938
rect 243834 533258 243866 533494
rect 244102 533258 244186 533494
rect 244422 533258 244454 533494
rect 243834 533174 244454 533258
rect 243834 532938 243866 533174
rect 244102 532938 244186 533174
rect 244422 532938 244454 533174
rect 243834 497494 244454 532938
rect 243834 497258 243866 497494
rect 244102 497258 244186 497494
rect 244422 497258 244454 497494
rect 243834 497174 244454 497258
rect 243834 496938 243866 497174
rect 244102 496938 244186 497174
rect 244422 496938 244454 497174
rect 243834 461494 244454 496938
rect 243834 461258 243866 461494
rect 244102 461258 244186 461494
rect 244422 461258 244454 461494
rect 243834 461174 244454 461258
rect 243834 460938 243866 461174
rect 244102 460938 244186 461174
rect 244422 460938 244454 461174
rect 243834 425494 244454 460938
rect 243834 425258 243866 425494
rect 244102 425258 244186 425494
rect 244422 425258 244454 425494
rect 243834 425174 244454 425258
rect 243834 424938 243866 425174
rect 244102 424938 244186 425174
rect 244422 424938 244454 425174
rect 243834 389494 244454 424938
rect 243834 389258 243866 389494
rect 244102 389258 244186 389494
rect 244422 389258 244454 389494
rect 243834 389174 244454 389258
rect 243834 388938 243866 389174
rect 244102 388938 244186 389174
rect 244422 388938 244454 389174
rect 243834 353494 244454 388938
rect 243834 353258 243866 353494
rect 244102 353258 244186 353494
rect 244422 353258 244454 353494
rect 243834 353174 244454 353258
rect 243834 352938 243866 353174
rect 244102 352938 244186 353174
rect 244422 352938 244454 353174
rect 243834 317494 244454 352938
rect 243834 317258 243866 317494
rect 244102 317258 244186 317494
rect 244422 317258 244454 317494
rect 243834 317174 244454 317258
rect 243834 316938 243866 317174
rect 244102 316938 244186 317174
rect 244422 316938 244454 317174
rect 243834 281494 244454 316938
rect 243834 281258 243866 281494
rect 244102 281258 244186 281494
rect 244422 281258 244454 281494
rect 243834 281174 244454 281258
rect 243834 280938 243866 281174
rect 244102 280938 244186 281174
rect 244422 280938 244454 281174
rect 243834 245494 244454 280938
rect 243834 245258 243866 245494
rect 244102 245258 244186 245494
rect 244422 245258 244454 245494
rect 243834 245174 244454 245258
rect 243834 244938 243866 245174
rect 244102 244938 244186 245174
rect 244422 244938 244454 245174
rect 243834 209494 244454 244938
rect 243834 209258 243866 209494
rect 244102 209258 244186 209494
rect 244422 209258 244454 209494
rect 243834 209174 244454 209258
rect 243834 208938 243866 209174
rect 244102 208938 244186 209174
rect 244422 208938 244454 209174
rect 243834 173494 244454 208938
rect 243834 173258 243866 173494
rect 244102 173258 244186 173494
rect 244422 173258 244454 173494
rect 243834 173174 244454 173258
rect 243834 172938 243866 173174
rect 244102 172938 244186 173174
rect 244422 172938 244454 173174
rect 243834 137494 244454 172938
rect 243834 137258 243866 137494
rect 244102 137258 244186 137494
rect 244422 137258 244454 137494
rect 243834 137174 244454 137258
rect 243834 136938 243866 137174
rect 244102 136938 244186 137174
rect 244422 136938 244454 137174
rect 243834 101494 244454 136938
rect 243834 101258 243866 101494
rect 244102 101258 244186 101494
rect 244422 101258 244454 101494
rect 243834 101174 244454 101258
rect 243834 100938 243866 101174
rect 244102 100938 244186 101174
rect 244422 100938 244454 101174
rect 243834 65494 244454 100938
rect 243834 65258 243866 65494
rect 244102 65258 244186 65494
rect 244422 65258 244454 65494
rect 243834 65174 244454 65258
rect 243834 64938 243866 65174
rect 244102 64938 244186 65174
rect 244422 64938 244454 65174
rect 243834 29494 244454 64938
rect 251774 52733 251834 670651
rect 253794 651454 254414 686898
rect 253794 651218 253826 651454
rect 254062 651218 254146 651454
rect 254382 651218 254414 651454
rect 253794 651134 254414 651218
rect 253794 650898 253826 651134
rect 254062 650898 254146 651134
rect 254382 650898 254414 651134
rect 253794 615454 254414 650898
rect 257514 705798 258134 711590
rect 257514 705562 257546 705798
rect 257782 705562 257866 705798
rect 258102 705562 258134 705798
rect 257514 705478 258134 705562
rect 257514 705242 257546 705478
rect 257782 705242 257866 705478
rect 258102 705242 258134 705478
rect 257514 691174 258134 705242
rect 257514 690938 257546 691174
rect 257782 690938 257866 691174
rect 258102 690938 258134 691174
rect 257514 690854 258134 690938
rect 257514 690618 257546 690854
rect 257782 690618 257866 690854
rect 258102 690618 258134 690854
rect 257514 655174 258134 690618
rect 257514 654938 257546 655174
rect 257782 654938 257866 655174
rect 258102 654938 258134 655174
rect 257514 654854 258134 654938
rect 257514 654618 257546 654854
rect 257782 654618 257866 654854
rect 258102 654618 258134 654854
rect 257514 649212 258134 654618
rect 261234 706758 261854 711590
rect 261234 706522 261266 706758
rect 261502 706522 261586 706758
rect 261822 706522 261854 706758
rect 261234 706438 261854 706522
rect 261234 706202 261266 706438
rect 261502 706202 261586 706438
rect 261822 706202 261854 706438
rect 261234 694894 261854 706202
rect 261234 694658 261266 694894
rect 261502 694658 261586 694894
rect 261822 694658 261854 694894
rect 261234 694574 261854 694658
rect 261234 694338 261266 694574
rect 261502 694338 261586 694574
rect 261822 694338 261854 694574
rect 261234 658894 261854 694338
rect 261234 658658 261266 658894
rect 261502 658658 261586 658894
rect 261822 658658 261854 658894
rect 261234 658574 261854 658658
rect 261234 658338 261266 658574
rect 261502 658338 261586 658574
rect 261822 658338 261854 658574
rect 261234 648313 261854 658338
rect 264954 707718 265574 711590
rect 264954 707482 264986 707718
rect 265222 707482 265306 707718
rect 265542 707482 265574 707718
rect 264954 707398 265574 707482
rect 264954 707162 264986 707398
rect 265222 707162 265306 707398
rect 265542 707162 265574 707398
rect 264954 698614 265574 707162
rect 264954 698378 264986 698614
rect 265222 698378 265306 698614
rect 265542 698378 265574 698614
rect 264954 698294 265574 698378
rect 264954 698058 264986 698294
rect 265222 698058 265306 698294
rect 265542 698058 265574 698294
rect 264954 662614 265574 698058
rect 264954 662378 264986 662614
rect 265222 662378 265306 662614
rect 265542 662378 265574 662614
rect 264954 662294 265574 662378
rect 264954 662058 264986 662294
rect 265222 662058 265306 662294
rect 265542 662058 265574 662294
rect 264954 648313 265574 662058
rect 268674 708678 269294 711590
rect 268674 708442 268706 708678
rect 268942 708442 269026 708678
rect 269262 708442 269294 708678
rect 268674 708358 269294 708442
rect 268674 708122 268706 708358
rect 268942 708122 269026 708358
rect 269262 708122 269294 708358
rect 268674 666334 269294 708122
rect 268674 666098 268706 666334
rect 268942 666098 269026 666334
rect 269262 666098 269294 666334
rect 268674 666014 269294 666098
rect 268674 665778 268706 666014
rect 268942 665778 269026 666014
rect 269262 665778 269294 666014
rect 268674 648313 269294 665778
rect 272394 709638 273014 711590
rect 272394 709402 272426 709638
rect 272662 709402 272746 709638
rect 272982 709402 273014 709638
rect 272394 709318 273014 709402
rect 272394 709082 272426 709318
rect 272662 709082 272746 709318
rect 272982 709082 273014 709318
rect 272394 670054 273014 709082
rect 272394 669818 272426 670054
rect 272662 669818 272746 670054
rect 272982 669818 273014 670054
rect 272394 669734 273014 669818
rect 272394 669498 272426 669734
rect 272662 669498 272746 669734
rect 272982 669498 273014 669734
rect 272394 648313 273014 669498
rect 276114 710598 276734 711590
rect 276114 710362 276146 710598
rect 276382 710362 276466 710598
rect 276702 710362 276734 710598
rect 276114 710278 276734 710362
rect 276114 710042 276146 710278
rect 276382 710042 276466 710278
rect 276702 710042 276734 710278
rect 276114 673774 276734 710042
rect 276114 673538 276146 673774
rect 276382 673538 276466 673774
rect 276702 673538 276734 673774
rect 276114 673454 276734 673538
rect 276114 673218 276146 673454
rect 276382 673218 276466 673454
rect 276702 673218 276734 673454
rect 276114 648313 276734 673218
rect 279834 711558 280454 711590
rect 279834 711322 279866 711558
rect 280102 711322 280186 711558
rect 280422 711322 280454 711558
rect 279834 711238 280454 711322
rect 279834 711002 279866 711238
rect 280102 711002 280186 711238
rect 280422 711002 280454 711238
rect 279834 677494 280454 711002
rect 279834 677258 279866 677494
rect 280102 677258 280186 677494
rect 280422 677258 280454 677494
rect 279834 677174 280454 677258
rect 279834 676938 279866 677174
rect 280102 676938 280186 677174
rect 280422 676938 280454 677174
rect 279834 648313 280454 676938
rect 289794 704838 290414 711590
rect 289794 704602 289826 704838
rect 290062 704602 290146 704838
rect 290382 704602 290414 704838
rect 289794 704518 290414 704602
rect 289794 704282 289826 704518
rect 290062 704282 290146 704518
rect 290382 704282 290414 704518
rect 289794 687454 290414 704282
rect 289794 687218 289826 687454
rect 290062 687218 290146 687454
rect 290382 687218 290414 687454
rect 289794 687134 290414 687218
rect 289794 686898 289826 687134
rect 290062 686898 290146 687134
rect 290382 686898 290414 687134
rect 289794 651454 290414 686898
rect 289794 651218 289826 651454
rect 290062 651218 290146 651454
rect 290382 651218 290414 651454
rect 289794 651134 290414 651218
rect 289794 650898 289826 651134
rect 290062 650898 290146 651134
rect 290382 650898 290414 651134
rect 289794 648313 290414 650898
rect 293514 705798 294134 711590
rect 293514 705562 293546 705798
rect 293782 705562 293866 705798
rect 294102 705562 294134 705798
rect 293514 705478 294134 705562
rect 293514 705242 293546 705478
rect 293782 705242 293866 705478
rect 294102 705242 294134 705478
rect 293514 691174 294134 705242
rect 293514 690938 293546 691174
rect 293782 690938 293866 691174
rect 294102 690938 294134 691174
rect 293514 690854 294134 690938
rect 293514 690618 293546 690854
rect 293782 690618 293866 690854
rect 294102 690618 294134 690854
rect 293514 655174 294134 690618
rect 293514 654938 293546 655174
rect 293782 654938 293866 655174
rect 294102 654938 294134 655174
rect 293514 654854 294134 654938
rect 293514 654618 293546 654854
rect 293782 654618 293866 654854
rect 294102 654618 294134 654854
rect 293514 648313 294134 654618
rect 297234 706758 297854 711590
rect 297234 706522 297266 706758
rect 297502 706522 297586 706758
rect 297822 706522 297854 706758
rect 297234 706438 297854 706522
rect 297234 706202 297266 706438
rect 297502 706202 297586 706438
rect 297822 706202 297854 706438
rect 297234 694894 297854 706202
rect 297234 694658 297266 694894
rect 297502 694658 297586 694894
rect 297822 694658 297854 694894
rect 297234 694574 297854 694658
rect 297234 694338 297266 694574
rect 297502 694338 297586 694574
rect 297822 694338 297854 694574
rect 297234 658894 297854 694338
rect 297234 658658 297266 658894
rect 297502 658658 297586 658894
rect 297822 658658 297854 658894
rect 297234 658574 297854 658658
rect 297234 658338 297266 658574
rect 297502 658338 297586 658574
rect 297822 658338 297854 658574
rect 297234 648313 297854 658338
rect 300954 707718 301574 711590
rect 300954 707482 300986 707718
rect 301222 707482 301306 707718
rect 301542 707482 301574 707718
rect 300954 707398 301574 707482
rect 300954 707162 300986 707398
rect 301222 707162 301306 707398
rect 301542 707162 301574 707398
rect 300954 698614 301574 707162
rect 300954 698378 300986 698614
rect 301222 698378 301306 698614
rect 301542 698378 301574 698614
rect 300954 698294 301574 698378
rect 300954 698058 300986 698294
rect 301222 698058 301306 698294
rect 301542 698058 301574 698294
rect 300954 662614 301574 698058
rect 300954 662378 300986 662614
rect 301222 662378 301306 662614
rect 301542 662378 301574 662614
rect 300954 662294 301574 662378
rect 300954 662058 300986 662294
rect 301222 662058 301306 662294
rect 301542 662058 301574 662294
rect 300954 648313 301574 662058
rect 304674 708678 305294 711590
rect 304674 708442 304706 708678
rect 304942 708442 305026 708678
rect 305262 708442 305294 708678
rect 304674 708358 305294 708442
rect 304674 708122 304706 708358
rect 304942 708122 305026 708358
rect 305262 708122 305294 708358
rect 304674 666334 305294 708122
rect 304674 666098 304706 666334
rect 304942 666098 305026 666334
rect 305262 666098 305294 666334
rect 304674 666014 305294 666098
rect 304674 665778 304706 666014
rect 304942 665778 305026 666014
rect 305262 665778 305294 666014
rect 304674 648313 305294 665778
rect 308394 709638 309014 711590
rect 308394 709402 308426 709638
rect 308662 709402 308746 709638
rect 308982 709402 309014 709638
rect 308394 709318 309014 709402
rect 308394 709082 308426 709318
rect 308662 709082 308746 709318
rect 308982 709082 309014 709318
rect 308394 670054 309014 709082
rect 308394 669818 308426 670054
rect 308662 669818 308746 670054
rect 308982 669818 309014 670054
rect 308394 669734 309014 669818
rect 308394 669498 308426 669734
rect 308662 669498 308746 669734
rect 308982 669498 309014 669734
rect 308394 648313 309014 669498
rect 312114 710598 312734 711590
rect 312114 710362 312146 710598
rect 312382 710362 312466 710598
rect 312702 710362 312734 710598
rect 312114 710278 312734 710362
rect 312114 710042 312146 710278
rect 312382 710042 312466 710278
rect 312702 710042 312734 710278
rect 312114 673774 312734 710042
rect 312114 673538 312146 673774
rect 312382 673538 312466 673774
rect 312702 673538 312734 673774
rect 312114 673454 312734 673538
rect 312114 673218 312146 673454
rect 312382 673218 312466 673454
rect 312702 673218 312734 673454
rect 312114 648313 312734 673218
rect 315834 711558 316454 711590
rect 315834 711322 315866 711558
rect 316102 711322 316186 711558
rect 316422 711322 316454 711558
rect 315834 711238 316454 711322
rect 315834 711002 315866 711238
rect 316102 711002 316186 711238
rect 316422 711002 316454 711238
rect 315834 677494 316454 711002
rect 315834 677258 315866 677494
rect 316102 677258 316186 677494
rect 316422 677258 316454 677494
rect 315834 677174 316454 677258
rect 315834 676938 315866 677174
rect 316102 676938 316186 677174
rect 316422 676938 316454 677174
rect 315834 648313 316454 676938
rect 325794 704838 326414 711590
rect 325794 704602 325826 704838
rect 326062 704602 326146 704838
rect 326382 704602 326414 704838
rect 325794 704518 326414 704602
rect 325794 704282 325826 704518
rect 326062 704282 326146 704518
rect 326382 704282 326414 704518
rect 325794 687454 326414 704282
rect 325794 687218 325826 687454
rect 326062 687218 326146 687454
rect 326382 687218 326414 687454
rect 325794 687134 326414 687218
rect 325794 686898 325826 687134
rect 326062 686898 326146 687134
rect 326382 686898 326414 687134
rect 325794 651454 326414 686898
rect 325794 651218 325826 651454
rect 326062 651218 326146 651454
rect 326382 651218 326414 651454
rect 325794 651134 326414 651218
rect 325794 650898 325826 651134
rect 326062 650898 326146 651134
rect 326382 650898 326414 651134
rect 325794 648313 326414 650898
rect 329514 705798 330134 711590
rect 329514 705562 329546 705798
rect 329782 705562 329866 705798
rect 330102 705562 330134 705798
rect 329514 705478 330134 705562
rect 329514 705242 329546 705478
rect 329782 705242 329866 705478
rect 330102 705242 330134 705478
rect 329514 691174 330134 705242
rect 329514 690938 329546 691174
rect 329782 690938 329866 691174
rect 330102 690938 330134 691174
rect 329514 690854 330134 690938
rect 329514 690618 329546 690854
rect 329782 690618 329866 690854
rect 330102 690618 330134 690854
rect 329514 655174 330134 690618
rect 329514 654938 329546 655174
rect 329782 654938 329866 655174
rect 330102 654938 330134 655174
rect 329514 654854 330134 654938
rect 329514 654618 329546 654854
rect 329782 654618 329866 654854
rect 330102 654618 330134 654854
rect 329514 648313 330134 654618
rect 333234 706758 333854 711590
rect 333234 706522 333266 706758
rect 333502 706522 333586 706758
rect 333822 706522 333854 706758
rect 333234 706438 333854 706522
rect 333234 706202 333266 706438
rect 333502 706202 333586 706438
rect 333822 706202 333854 706438
rect 333234 694894 333854 706202
rect 333234 694658 333266 694894
rect 333502 694658 333586 694894
rect 333822 694658 333854 694894
rect 333234 694574 333854 694658
rect 333234 694338 333266 694574
rect 333502 694338 333586 694574
rect 333822 694338 333854 694574
rect 333234 658894 333854 694338
rect 333234 658658 333266 658894
rect 333502 658658 333586 658894
rect 333822 658658 333854 658894
rect 333234 658574 333854 658658
rect 333234 658338 333266 658574
rect 333502 658338 333586 658574
rect 333822 658338 333854 658574
rect 333234 648313 333854 658338
rect 336954 707718 337574 711590
rect 336954 707482 336986 707718
rect 337222 707482 337306 707718
rect 337542 707482 337574 707718
rect 336954 707398 337574 707482
rect 336954 707162 336986 707398
rect 337222 707162 337306 707398
rect 337542 707162 337574 707398
rect 336954 698614 337574 707162
rect 336954 698378 336986 698614
rect 337222 698378 337306 698614
rect 337542 698378 337574 698614
rect 336954 698294 337574 698378
rect 336954 698058 336986 698294
rect 337222 698058 337306 698294
rect 337542 698058 337574 698294
rect 336954 662614 337574 698058
rect 336954 662378 336986 662614
rect 337222 662378 337306 662614
rect 337542 662378 337574 662614
rect 336954 662294 337574 662378
rect 336954 662058 336986 662294
rect 337222 662058 337306 662294
rect 337542 662058 337574 662294
rect 336954 648313 337574 662058
rect 340674 708678 341294 711590
rect 340674 708442 340706 708678
rect 340942 708442 341026 708678
rect 341262 708442 341294 708678
rect 340674 708358 341294 708442
rect 340674 708122 340706 708358
rect 340942 708122 341026 708358
rect 341262 708122 341294 708358
rect 340674 666334 341294 708122
rect 340674 666098 340706 666334
rect 340942 666098 341026 666334
rect 341262 666098 341294 666334
rect 340674 666014 341294 666098
rect 340674 665778 340706 666014
rect 340942 665778 341026 666014
rect 341262 665778 341294 666014
rect 340674 648313 341294 665778
rect 344394 709638 345014 711590
rect 344394 709402 344426 709638
rect 344662 709402 344746 709638
rect 344982 709402 345014 709638
rect 344394 709318 345014 709402
rect 344394 709082 344426 709318
rect 344662 709082 344746 709318
rect 344982 709082 345014 709318
rect 344394 670054 345014 709082
rect 344394 669818 344426 670054
rect 344662 669818 344746 670054
rect 344982 669818 345014 670054
rect 344394 669734 345014 669818
rect 344394 669498 344426 669734
rect 344662 669498 344746 669734
rect 344982 669498 345014 669734
rect 344394 648313 345014 669498
rect 348114 710598 348734 711590
rect 348114 710362 348146 710598
rect 348382 710362 348466 710598
rect 348702 710362 348734 710598
rect 348114 710278 348734 710362
rect 348114 710042 348146 710278
rect 348382 710042 348466 710278
rect 348702 710042 348734 710278
rect 348114 673774 348734 710042
rect 348114 673538 348146 673774
rect 348382 673538 348466 673774
rect 348702 673538 348734 673774
rect 348114 673454 348734 673538
rect 348114 673218 348146 673454
rect 348382 673218 348466 673454
rect 348702 673218 348734 673454
rect 348114 648313 348734 673218
rect 351834 711558 352454 711590
rect 351834 711322 351866 711558
rect 352102 711322 352186 711558
rect 352422 711322 352454 711558
rect 351834 711238 352454 711322
rect 351834 711002 351866 711238
rect 352102 711002 352186 711238
rect 352422 711002 352454 711238
rect 351834 677494 352454 711002
rect 351834 677258 351866 677494
rect 352102 677258 352186 677494
rect 352422 677258 352454 677494
rect 351834 677174 352454 677258
rect 351834 676938 351866 677174
rect 352102 676938 352186 677174
rect 352422 676938 352454 677174
rect 351834 648313 352454 676938
rect 361794 704838 362414 711590
rect 361794 704602 361826 704838
rect 362062 704602 362146 704838
rect 362382 704602 362414 704838
rect 361794 704518 362414 704602
rect 361794 704282 361826 704518
rect 362062 704282 362146 704518
rect 362382 704282 362414 704518
rect 361794 687454 362414 704282
rect 361794 687218 361826 687454
rect 362062 687218 362146 687454
rect 362382 687218 362414 687454
rect 361794 687134 362414 687218
rect 361794 686898 361826 687134
rect 362062 686898 362146 687134
rect 362382 686898 362414 687134
rect 361794 651454 362414 686898
rect 361794 651218 361826 651454
rect 362062 651218 362146 651454
rect 362382 651218 362414 651454
rect 361794 651134 362414 651218
rect 361794 650898 361826 651134
rect 362062 650898 362146 651134
rect 362382 650898 362414 651134
rect 361794 648313 362414 650898
rect 365514 705798 366134 711590
rect 365514 705562 365546 705798
rect 365782 705562 365866 705798
rect 366102 705562 366134 705798
rect 365514 705478 366134 705562
rect 365514 705242 365546 705478
rect 365782 705242 365866 705478
rect 366102 705242 366134 705478
rect 365514 691174 366134 705242
rect 365514 690938 365546 691174
rect 365782 690938 365866 691174
rect 366102 690938 366134 691174
rect 365514 690854 366134 690938
rect 365514 690618 365546 690854
rect 365782 690618 365866 690854
rect 366102 690618 366134 690854
rect 365514 655174 366134 690618
rect 365514 654938 365546 655174
rect 365782 654938 365866 655174
rect 366102 654938 366134 655174
rect 365514 654854 366134 654938
rect 365514 654618 365546 654854
rect 365782 654618 365866 654854
rect 366102 654618 366134 654854
rect 365514 649212 366134 654618
rect 369234 706758 369854 711590
rect 369234 706522 369266 706758
rect 369502 706522 369586 706758
rect 369822 706522 369854 706758
rect 369234 706438 369854 706522
rect 369234 706202 369266 706438
rect 369502 706202 369586 706438
rect 369822 706202 369854 706438
rect 369234 694894 369854 706202
rect 369234 694658 369266 694894
rect 369502 694658 369586 694894
rect 369822 694658 369854 694894
rect 369234 694574 369854 694658
rect 369234 694338 369266 694574
rect 369502 694338 369586 694574
rect 369822 694338 369854 694574
rect 369234 658894 369854 694338
rect 369234 658658 369266 658894
rect 369502 658658 369586 658894
rect 369822 658658 369854 658894
rect 369234 658574 369854 658658
rect 369234 658338 369266 658574
rect 369502 658338 369586 658574
rect 369822 658338 369854 658574
rect 369234 648313 369854 658338
rect 372954 707718 373574 711590
rect 372954 707482 372986 707718
rect 373222 707482 373306 707718
rect 373542 707482 373574 707718
rect 372954 707398 373574 707482
rect 372954 707162 372986 707398
rect 373222 707162 373306 707398
rect 373542 707162 373574 707398
rect 372954 698614 373574 707162
rect 372954 698378 372986 698614
rect 373222 698378 373306 698614
rect 373542 698378 373574 698614
rect 372954 698294 373574 698378
rect 372954 698058 372986 698294
rect 373222 698058 373306 698294
rect 373542 698058 373574 698294
rect 372954 662614 373574 698058
rect 372954 662378 372986 662614
rect 373222 662378 373306 662614
rect 373542 662378 373574 662614
rect 372954 662294 373574 662378
rect 372954 662058 372986 662294
rect 373222 662058 373306 662294
rect 373542 662058 373574 662294
rect 372954 648313 373574 662058
rect 376674 708678 377294 711590
rect 376674 708442 376706 708678
rect 376942 708442 377026 708678
rect 377262 708442 377294 708678
rect 376674 708358 377294 708442
rect 376674 708122 376706 708358
rect 376942 708122 377026 708358
rect 377262 708122 377294 708358
rect 376674 666334 377294 708122
rect 376674 666098 376706 666334
rect 376942 666098 377026 666334
rect 377262 666098 377294 666334
rect 376674 666014 377294 666098
rect 376674 665778 376706 666014
rect 376942 665778 377026 666014
rect 377262 665778 377294 666014
rect 376674 648313 377294 665778
rect 380394 709638 381014 711590
rect 380394 709402 380426 709638
rect 380662 709402 380746 709638
rect 380982 709402 381014 709638
rect 380394 709318 381014 709402
rect 380394 709082 380426 709318
rect 380662 709082 380746 709318
rect 380982 709082 381014 709318
rect 380394 670054 381014 709082
rect 380394 669818 380426 670054
rect 380662 669818 380746 670054
rect 380982 669818 381014 670054
rect 380394 669734 381014 669818
rect 380394 669498 380426 669734
rect 380662 669498 380746 669734
rect 380982 669498 381014 669734
rect 380394 649212 381014 669498
rect 384114 710598 384734 711590
rect 384114 710362 384146 710598
rect 384382 710362 384466 710598
rect 384702 710362 384734 710598
rect 384114 710278 384734 710362
rect 384114 710042 384146 710278
rect 384382 710042 384466 710278
rect 384702 710042 384734 710278
rect 384114 673774 384734 710042
rect 384114 673538 384146 673774
rect 384382 673538 384466 673774
rect 384702 673538 384734 673774
rect 384114 673454 384734 673538
rect 384114 673218 384146 673454
rect 384382 673218 384466 673454
rect 384702 673218 384734 673454
rect 384114 648313 384734 673218
rect 387834 711558 388454 711590
rect 387834 711322 387866 711558
rect 388102 711322 388186 711558
rect 388422 711322 388454 711558
rect 387834 711238 388454 711322
rect 387834 711002 387866 711238
rect 388102 711002 388186 711238
rect 388422 711002 388454 711238
rect 387834 677494 388454 711002
rect 387834 677258 387866 677494
rect 388102 677258 388186 677494
rect 388422 677258 388454 677494
rect 387834 677174 388454 677258
rect 387834 676938 387866 677174
rect 388102 676938 388186 677174
rect 388422 676938 388454 677174
rect 387834 648313 388454 676938
rect 397794 704838 398414 711590
rect 397794 704602 397826 704838
rect 398062 704602 398146 704838
rect 398382 704602 398414 704838
rect 397794 704518 398414 704602
rect 397794 704282 397826 704518
rect 398062 704282 398146 704518
rect 398382 704282 398414 704518
rect 397794 687454 398414 704282
rect 397794 687218 397826 687454
rect 398062 687218 398146 687454
rect 398382 687218 398414 687454
rect 397794 687134 398414 687218
rect 397794 686898 397826 687134
rect 398062 686898 398146 687134
rect 398382 686898 398414 687134
rect 397794 651454 398414 686898
rect 397794 651218 397826 651454
rect 398062 651218 398146 651454
rect 398382 651218 398414 651454
rect 397794 651134 398414 651218
rect 397794 650898 397826 651134
rect 398062 650898 398146 651134
rect 398382 650898 398414 651134
rect 397794 648313 398414 650898
rect 401514 705798 402134 711590
rect 401514 705562 401546 705798
rect 401782 705562 401866 705798
rect 402102 705562 402134 705798
rect 401514 705478 402134 705562
rect 401514 705242 401546 705478
rect 401782 705242 401866 705478
rect 402102 705242 402134 705478
rect 401514 691174 402134 705242
rect 401514 690938 401546 691174
rect 401782 690938 401866 691174
rect 402102 690938 402134 691174
rect 401514 690854 402134 690938
rect 401514 690618 401546 690854
rect 401782 690618 401866 690854
rect 402102 690618 402134 690854
rect 401514 655174 402134 690618
rect 401514 654938 401546 655174
rect 401782 654938 401866 655174
rect 402102 654938 402134 655174
rect 401514 654854 402134 654938
rect 401514 654618 401546 654854
rect 401782 654618 401866 654854
rect 402102 654618 402134 654854
rect 401514 648313 402134 654618
rect 405234 706758 405854 711590
rect 405234 706522 405266 706758
rect 405502 706522 405586 706758
rect 405822 706522 405854 706758
rect 405234 706438 405854 706522
rect 405234 706202 405266 706438
rect 405502 706202 405586 706438
rect 405822 706202 405854 706438
rect 405234 694894 405854 706202
rect 405234 694658 405266 694894
rect 405502 694658 405586 694894
rect 405822 694658 405854 694894
rect 405234 694574 405854 694658
rect 405234 694338 405266 694574
rect 405502 694338 405586 694574
rect 405822 694338 405854 694574
rect 405234 658894 405854 694338
rect 405234 658658 405266 658894
rect 405502 658658 405586 658894
rect 405822 658658 405854 658894
rect 405234 658574 405854 658658
rect 405234 658338 405266 658574
rect 405502 658338 405586 658574
rect 405822 658338 405854 658574
rect 405234 648313 405854 658338
rect 408954 707718 409574 711590
rect 408954 707482 408986 707718
rect 409222 707482 409306 707718
rect 409542 707482 409574 707718
rect 408954 707398 409574 707482
rect 408954 707162 408986 707398
rect 409222 707162 409306 707398
rect 409542 707162 409574 707398
rect 408954 698614 409574 707162
rect 408954 698378 408986 698614
rect 409222 698378 409306 698614
rect 409542 698378 409574 698614
rect 408954 698294 409574 698378
rect 408954 698058 408986 698294
rect 409222 698058 409306 698294
rect 409542 698058 409574 698294
rect 408954 662614 409574 698058
rect 408954 662378 408986 662614
rect 409222 662378 409306 662614
rect 409542 662378 409574 662614
rect 408954 662294 409574 662378
rect 408954 662058 408986 662294
rect 409222 662058 409306 662294
rect 409542 662058 409574 662294
rect 408954 648313 409574 662058
rect 412674 708678 413294 711590
rect 412674 708442 412706 708678
rect 412942 708442 413026 708678
rect 413262 708442 413294 708678
rect 412674 708358 413294 708442
rect 412674 708122 412706 708358
rect 412942 708122 413026 708358
rect 413262 708122 413294 708358
rect 412674 666334 413294 708122
rect 412674 666098 412706 666334
rect 412942 666098 413026 666334
rect 413262 666098 413294 666334
rect 412674 666014 413294 666098
rect 412674 665778 412706 666014
rect 412942 665778 413026 666014
rect 413262 665778 413294 666014
rect 412674 648313 413294 665778
rect 416394 709638 417014 711590
rect 416394 709402 416426 709638
rect 416662 709402 416746 709638
rect 416982 709402 417014 709638
rect 416394 709318 417014 709402
rect 416394 709082 416426 709318
rect 416662 709082 416746 709318
rect 416982 709082 417014 709318
rect 416394 670054 417014 709082
rect 416394 669818 416426 670054
rect 416662 669818 416746 670054
rect 416982 669818 417014 670054
rect 416394 669734 417014 669818
rect 416394 669498 416426 669734
rect 416662 669498 416746 669734
rect 416982 669498 417014 669734
rect 416394 648313 417014 669498
rect 420114 710598 420734 711590
rect 420114 710362 420146 710598
rect 420382 710362 420466 710598
rect 420702 710362 420734 710598
rect 420114 710278 420734 710362
rect 420114 710042 420146 710278
rect 420382 710042 420466 710278
rect 420702 710042 420734 710278
rect 420114 673774 420734 710042
rect 420114 673538 420146 673774
rect 420382 673538 420466 673774
rect 420702 673538 420734 673774
rect 420114 673454 420734 673538
rect 420114 673218 420146 673454
rect 420382 673218 420466 673454
rect 420702 673218 420734 673454
rect 420114 648313 420734 673218
rect 423834 711558 424454 711590
rect 423834 711322 423866 711558
rect 424102 711322 424186 711558
rect 424422 711322 424454 711558
rect 423834 711238 424454 711322
rect 423834 711002 423866 711238
rect 424102 711002 424186 711238
rect 424422 711002 424454 711238
rect 423834 677494 424454 711002
rect 423834 677258 423866 677494
rect 424102 677258 424186 677494
rect 424422 677258 424454 677494
rect 423834 677174 424454 677258
rect 423834 676938 423866 677174
rect 424102 676938 424186 677174
rect 424422 676938 424454 677174
rect 423834 648313 424454 676938
rect 433794 704838 434414 711590
rect 433794 704602 433826 704838
rect 434062 704602 434146 704838
rect 434382 704602 434414 704838
rect 433794 704518 434414 704602
rect 433794 704282 433826 704518
rect 434062 704282 434146 704518
rect 434382 704282 434414 704518
rect 433794 687454 434414 704282
rect 433794 687218 433826 687454
rect 434062 687218 434146 687454
rect 434382 687218 434414 687454
rect 433794 687134 434414 687218
rect 433794 686898 433826 687134
rect 434062 686898 434146 687134
rect 434382 686898 434414 687134
rect 433794 651454 434414 686898
rect 433794 651218 433826 651454
rect 434062 651218 434146 651454
rect 434382 651218 434414 651454
rect 433794 651134 434414 651218
rect 433794 650898 433826 651134
rect 434062 650898 434146 651134
rect 434382 650898 434414 651134
rect 433794 648313 434414 650898
rect 437514 705798 438134 711590
rect 437514 705562 437546 705798
rect 437782 705562 437866 705798
rect 438102 705562 438134 705798
rect 437514 705478 438134 705562
rect 437514 705242 437546 705478
rect 437782 705242 437866 705478
rect 438102 705242 438134 705478
rect 437514 691174 438134 705242
rect 437514 690938 437546 691174
rect 437782 690938 437866 691174
rect 438102 690938 438134 691174
rect 437514 690854 438134 690938
rect 437514 690618 437546 690854
rect 437782 690618 437866 690854
rect 438102 690618 438134 690854
rect 437514 655174 438134 690618
rect 437514 654938 437546 655174
rect 437782 654938 437866 655174
rect 438102 654938 438134 655174
rect 437514 654854 438134 654938
rect 437514 654618 437546 654854
rect 437782 654618 437866 654854
rect 438102 654618 438134 654854
rect 437514 648313 438134 654618
rect 441234 706758 441854 711590
rect 441234 706522 441266 706758
rect 441502 706522 441586 706758
rect 441822 706522 441854 706758
rect 441234 706438 441854 706522
rect 441234 706202 441266 706438
rect 441502 706202 441586 706438
rect 441822 706202 441854 706438
rect 441234 694894 441854 706202
rect 441234 694658 441266 694894
rect 441502 694658 441586 694894
rect 441822 694658 441854 694894
rect 441234 694574 441854 694658
rect 441234 694338 441266 694574
rect 441502 694338 441586 694574
rect 441822 694338 441854 694574
rect 441234 658894 441854 694338
rect 441234 658658 441266 658894
rect 441502 658658 441586 658894
rect 441822 658658 441854 658894
rect 441234 658574 441854 658658
rect 441234 658338 441266 658574
rect 441502 658338 441586 658574
rect 441822 658338 441854 658574
rect 441234 648313 441854 658338
rect 444954 707718 445574 711590
rect 444954 707482 444986 707718
rect 445222 707482 445306 707718
rect 445542 707482 445574 707718
rect 444954 707398 445574 707482
rect 444954 707162 444986 707398
rect 445222 707162 445306 707398
rect 445542 707162 445574 707398
rect 444954 698614 445574 707162
rect 444954 698378 444986 698614
rect 445222 698378 445306 698614
rect 445542 698378 445574 698614
rect 444954 698294 445574 698378
rect 444954 698058 444986 698294
rect 445222 698058 445306 698294
rect 445542 698058 445574 698294
rect 444954 662614 445574 698058
rect 444954 662378 444986 662614
rect 445222 662378 445306 662614
rect 445542 662378 445574 662614
rect 444954 662294 445574 662378
rect 444954 662058 444986 662294
rect 445222 662058 445306 662294
rect 445542 662058 445574 662294
rect 444954 648313 445574 662058
rect 448674 708678 449294 711590
rect 448674 708442 448706 708678
rect 448942 708442 449026 708678
rect 449262 708442 449294 708678
rect 448674 708358 449294 708442
rect 448674 708122 448706 708358
rect 448942 708122 449026 708358
rect 449262 708122 449294 708358
rect 448674 666334 449294 708122
rect 448674 666098 448706 666334
rect 448942 666098 449026 666334
rect 449262 666098 449294 666334
rect 448674 666014 449294 666098
rect 448674 665778 448706 666014
rect 448942 665778 449026 666014
rect 449262 665778 449294 666014
rect 448674 648313 449294 665778
rect 452394 709638 453014 711590
rect 452394 709402 452426 709638
rect 452662 709402 452746 709638
rect 452982 709402 453014 709638
rect 452394 709318 453014 709402
rect 452394 709082 452426 709318
rect 452662 709082 452746 709318
rect 452982 709082 453014 709318
rect 452394 670054 453014 709082
rect 452394 669818 452426 670054
rect 452662 669818 452746 670054
rect 452982 669818 453014 670054
rect 452394 669734 453014 669818
rect 452394 669498 452426 669734
rect 452662 669498 452746 669734
rect 452982 669498 453014 669734
rect 452394 648313 453014 669498
rect 456114 710598 456734 711590
rect 456114 710362 456146 710598
rect 456382 710362 456466 710598
rect 456702 710362 456734 710598
rect 456114 710278 456734 710362
rect 456114 710042 456146 710278
rect 456382 710042 456466 710278
rect 456702 710042 456734 710278
rect 456114 673774 456734 710042
rect 456114 673538 456146 673774
rect 456382 673538 456466 673774
rect 456702 673538 456734 673774
rect 456114 673454 456734 673538
rect 456114 673218 456146 673454
rect 456382 673218 456466 673454
rect 456702 673218 456734 673454
rect 456114 648313 456734 673218
rect 459834 711558 460454 711590
rect 459834 711322 459866 711558
rect 460102 711322 460186 711558
rect 460422 711322 460454 711558
rect 459834 711238 460454 711322
rect 459834 711002 459866 711238
rect 460102 711002 460186 711238
rect 460422 711002 460454 711238
rect 459834 677494 460454 711002
rect 459834 677258 459866 677494
rect 460102 677258 460186 677494
rect 460422 677258 460454 677494
rect 459834 677174 460454 677258
rect 459834 676938 459866 677174
rect 460102 676938 460186 677174
rect 460422 676938 460454 677174
rect 459834 648313 460454 676938
rect 469794 704838 470414 711590
rect 469794 704602 469826 704838
rect 470062 704602 470146 704838
rect 470382 704602 470414 704838
rect 469794 704518 470414 704602
rect 469794 704282 469826 704518
rect 470062 704282 470146 704518
rect 470382 704282 470414 704518
rect 469794 687454 470414 704282
rect 469794 687218 469826 687454
rect 470062 687218 470146 687454
rect 470382 687218 470414 687454
rect 469794 687134 470414 687218
rect 469794 686898 469826 687134
rect 470062 686898 470146 687134
rect 470382 686898 470414 687134
rect 469794 651454 470414 686898
rect 469794 651218 469826 651454
rect 470062 651218 470146 651454
rect 470382 651218 470414 651454
rect 469794 651134 470414 651218
rect 469794 650898 469826 651134
rect 470062 650898 470146 651134
rect 470382 650898 470414 651134
rect 469794 648313 470414 650898
rect 473514 705798 474134 711590
rect 473514 705562 473546 705798
rect 473782 705562 473866 705798
rect 474102 705562 474134 705798
rect 473514 705478 474134 705562
rect 473514 705242 473546 705478
rect 473782 705242 473866 705478
rect 474102 705242 474134 705478
rect 473514 691174 474134 705242
rect 473514 690938 473546 691174
rect 473782 690938 473866 691174
rect 474102 690938 474134 691174
rect 473514 690854 474134 690938
rect 473514 690618 473546 690854
rect 473782 690618 473866 690854
rect 474102 690618 474134 690854
rect 473514 655174 474134 690618
rect 473514 654938 473546 655174
rect 473782 654938 473866 655174
rect 474102 654938 474134 655174
rect 473514 654854 474134 654938
rect 473514 654618 473546 654854
rect 473782 654618 473866 654854
rect 474102 654618 474134 654854
rect 473514 648313 474134 654618
rect 477234 706758 477854 711590
rect 477234 706522 477266 706758
rect 477502 706522 477586 706758
rect 477822 706522 477854 706758
rect 477234 706438 477854 706522
rect 477234 706202 477266 706438
rect 477502 706202 477586 706438
rect 477822 706202 477854 706438
rect 477234 694894 477854 706202
rect 477234 694658 477266 694894
rect 477502 694658 477586 694894
rect 477822 694658 477854 694894
rect 477234 694574 477854 694658
rect 477234 694338 477266 694574
rect 477502 694338 477586 694574
rect 477822 694338 477854 694574
rect 477234 658894 477854 694338
rect 477234 658658 477266 658894
rect 477502 658658 477586 658894
rect 477822 658658 477854 658894
rect 477234 658574 477854 658658
rect 477234 658338 477266 658574
rect 477502 658338 477586 658574
rect 477822 658338 477854 658574
rect 477234 648313 477854 658338
rect 480954 707718 481574 711590
rect 480954 707482 480986 707718
rect 481222 707482 481306 707718
rect 481542 707482 481574 707718
rect 480954 707398 481574 707482
rect 480954 707162 480986 707398
rect 481222 707162 481306 707398
rect 481542 707162 481574 707398
rect 480954 698614 481574 707162
rect 480954 698378 480986 698614
rect 481222 698378 481306 698614
rect 481542 698378 481574 698614
rect 480954 698294 481574 698378
rect 480954 698058 480986 698294
rect 481222 698058 481306 698294
rect 481542 698058 481574 698294
rect 480954 662614 481574 698058
rect 480954 662378 480986 662614
rect 481222 662378 481306 662614
rect 481542 662378 481574 662614
rect 480954 662294 481574 662378
rect 480954 662058 480986 662294
rect 481222 662058 481306 662294
rect 481542 662058 481574 662294
rect 480954 648313 481574 662058
rect 484674 708678 485294 711590
rect 484674 708442 484706 708678
rect 484942 708442 485026 708678
rect 485262 708442 485294 708678
rect 484674 708358 485294 708442
rect 484674 708122 484706 708358
rect 484942 708122 485026 708358
rect 485262 708122 485294 708358
rect 484674 666334 485294 708122
rect 484674 666098 484706 666334
rect 484942 666098 485026 666334
rect 485262 666098 485294 666334
rect 484674 666014 485294 666098
rect 484674 665778 484706 666014
rect 484942 665778 485026 666014
rect 485262 665778 485294 666014
rect 484674 648313 485294 665778
rect 488394 709638 489014 711590
rect 488394 709402 488426 709638
rect 488662 709402 488746 709638
rect 488982 709402 489014 709638
rect 488394 709318 489014 709402
rect 488394 709082 488426 709318
rect 488662 709082 488746 709318
rect 488982 709082 489014 709318
rect 488394 670054 489014 709082
rect 488394 669818 488426 670054
rect 488662 669818 488746 670054
rect 488982 669818 489014 670054
rect 488394 669734 489014 669818
rect 488394 669498 488426 669734
rect 488662 669498 488746 669734
rect 488982 669498 489014 669734
rect 488394 649212 489014 669498
rect 492114 710598 492734 711590
rect 492114 710362 492146 710598
rect 492382 710362 492466 710598
rect 492702 710362 492734 710598
rect 492114 710278 492734 710362
rect 492114 710042 492146 710278
rect 492382 710042 492466 710278
rect 492702 710042 492734 710278
rect 492114 673774 492734 710042
rect 492114 673538 492146 673774
rect 492382 673538 492466 673774
rect 492702 673538 492734 673774
rect 492114 673454 492734 673538
rect 492114 673218 492146 673454
rect 492382 673218 492466 673454
rect 492702 673218 492734 673454
rect 492114 648313 492734 673218
rect 495834 711558 496454 711590
rect 495834 711322 495866 711558
rect 496102 711322 496186 711558
rect 496422 711322 496454 711558
rect 495834 711238 496454 711322
rect 495834 711002 495866 711238
rect 496102 711002 496186 711238
rect 496422 711002 496454 711238
rect 495834 677494 496454 711002
rect 495834 677258 495866 677494
rect 496102 677258 496186 677494
rect 496422 677258 496454 677494
rect 495834 677174 496454 677258
rect 495834 676938 495866 677174
rect 496102 676938 496186 677174
rect 496422 676938 496454 677174
rect 495834 648313 496454 676938
rect 505794 704838 506414 711590
rect 505794 704602 505826 704838
rect 506062 704602 506146 704838
rect 506382 704602 506414 704838
rect 505794 704518 506414 704602
rect 505794 704282 505826 704518
rect 506062 704282 506146 704518
rect 506382 704282 506414 704518
rect 505794 687454 506414 704282
rect 505794 687218 505826 687454
rect 506062 687218 506146 687454
rect 506382 687218 506414 687454
rect 505794 687134 506414 687218
rect 505794 686898 505826 687134
rect 506062 686898 506146 687134
rect 506382 686898 506414 687134
rect 505794 651454 506414 686898
rect 505794 651218 505826 651454
rect 506062 651218 506146 651454
rect 506382 651218 506414 651454
rect 505794 651134 506414 651218
rect 505794 650898 505826 651134
rect 506062 650898 506146 651134
rect 506382 650898 506414 651134
rect 505794 648313 506414 650898
rect 509514 705798 510134 711590
rect 509514 705562 509546 705798
rect 509782 705562 509866 705798
rect 510102 705562 510134 705798
rect 509514 705478 510134 705562
rect 509514 705242 509546 705478
rect 509782 705242 509866 705478
rect 510102 705242 510134 705478
rect 509514 691174 510134 705242
rect 509514 690938 509546 691174
rect 509782 690938 509866 691174
rect 510102 690938 510134 691174
rect 509514 690854 510134 690938
rect 509514 690618 509546 690854
rect 509782 690618 509866 690854
rect 510102 690618 510134 690854
rect 509514 655174 510134 690618
rect 509514 654938 509546 655174
rect 509782 654938 509866 655174
rect 510102 654938 510134 655174
rect 509514 654854 510134 654938
rect 509514 654618 509546 654854
rect 509782 654618 509866 654854
rect 510102 654618 510134 654854
rect 509514 648313 510134 654618
rect 513234 706758 513854 711590
rect 513234 706522 513266 706758
rect 513502 706522 513586 706758
rect 513822 706522 513854 706758
rect 513234 706438 513854 706522
rect 513234 706202 513266 706438
rect 513502 706202 513586 706438
rect 513822 706202 513854 706438
rect 513234 694894 513854 706202
rect 513234 694658 513266 694894
rect 513502 694658 513586 694894
rect 513822 694658 513854 694894
rect 513234 694574 513854 694658
rect 513234 694338 513266 694574
rect 513502 694338 513586 694574
rect 513822 694338 513854 694574
rect 513234 658894 513854 694338
rect 513234 658658 513266 658894
rect 513502 658658 513586 658894
rect 513822 658658 513854 658894
rect 513234 658574 513854 658658
rect 513234 658338 513266 658574
rect 513502 658338 513586 658574
rect 513822 658338 513854 658574
rect 513234 648313 513854 658338
rect 516954 707718 517574 711590
rect 516954 707482 516986 707718
rect 517222 707482 517306 707718
rect 517542 707482 517574 707718
rect 516954 707398 517574 707482
rect 516954 707162 516986 707398
rect 517222 707162 517306 707398
rect 517542 707162 517574 707398
rect 516954 698614 517574 707162
rect 516954 698378 516986 698614
rect 517222 698378 517306 698614
rect 517542 698378 517574 698614
rect 516954 698294 517574 698378
rect 516954 698058 516986 698294
rect 517222 698058 517306 698294
rect 517542 698058 517574 698294
rect 516954 662614 517574 698058
rect 516954 662378 516986 662614
rect 517222 662378 517306 662614
rect 517542 662378 517574 662614
rect 516954 662294 517574 662378
rect 516954 662058 516986 662294
rect 517222 662058 517306 662294
rect 517542 662058 517574 662294
rect 516954 648313 517574 662058
rect 520674 708678 521294 711590
rect 520674 708442 520706 708678
rect 520942 708442 521026 708678
rect 521262 708442 521294 708678
rect 520674 708358 521294 708442
rect 520674 708122 520706 708358
rect 520942 708122 521026 708358
rect 521262 708122 521294 708358
rect 520674 666334 521294 708122
rect 520674 666098 520706 666334
rect 520942 666098 521026 666334
rect 521262 666098 521294 666334
rect 520674 666014 521294 666098
rect 520674 665778 520706 666014
rect 520942 665778 521026 666014
rect 521262 665778 521294 666014
rect 520674 648313 521294 665778
rect 524394 709638 525014 711590
rect 524394 709402 524426 709638
rect 524662 709402 524746 709638
rect 524982 709402 525014 709638
rect 524394 709318 525014 709402
rect 524394 709082 524426 709318
rect 524662 709082 524746 709318
rect 524982 709082 525014 709318
rect 524394 670054 525014 709082
rect 524394 669818 524426 670054
rect 524662 669818 524746 670054
rect 524982 669818 525014 670054
rect 524394 669734 525014 669818
rect 524394 669498 524426 669734
rect 524662 669498 524746 669734
rect 524982 669498 525014 669734
rect 524394 648313 525014 669498
rect 528114 710598 528734 711590
rect 528114 710362 528146 710598
rect 528382 710362 528466 710598
rect 528702 710362 528734 710598
rect 528114 710278 528734 710362
rect 528114 710042 528146 710278
rect 528382 710042 528466 710278
rect 528702 710042 528734 710278
rect 528114 673774 528734 710042
rect 528114 673538 528146 673774
rect 528382 673538 528466 673774
rect 528702 673538 528734 673774
rect 528114 673454 528734 673538
rect 528114 673218 528146 673454
rect 528382 673218 528466 673454
rect 528702 673218 528734 673454
rect 528114 648313 528734 673218
rect 531834 711558 532454 711590
rect 531834 711322 531866 711558
rect 532102 711322 532186 711558
rect 532422 711322 532454 711558
rect 531834 711238 532454 711322
rect 531834 711002 531866 711238
rect 532102 711002 532186 711238
rect 532422 711002 532454 711238
rect 531834 677494 532454 711002
rect 531834 677258 531866 677494
rect 532102 677258 532186 677494
rect 532422 677258 532454 677494
rect 531834 677174 532454 677258
rect 531834 676938 531866 677174
rect 532102 676938 532186 677174
rect 532422 676938 532454 677174
rect 531834 648313 532454 676938
rect 541794 704838 542414 711590
rect 541794 704602 541826 704838
rect 542062 704602 542146 704838
rect 542382 704602 542414 704838
rect 541794 704518 542414 704602
rect 541794 704282 541826 704518
rect 542062 704282 542146 704518
rect 542382 704282 542414 704518
rect 541794 687454 542414 704282
rect 541794 687218 541826 687454
rect 542062 687218 542146 687454
rect 542382 687218 542414 687454
rect 541794 687134 542414 687218
rect 541794 686898 541826 687134
rect 542062 686898 542146 687134
rect 542382 686898 542414 687134
rect 541794 651454 542414 686898
rect 541794 651218 541826 651454
rect 542062 651218 542146 651454
rect 542382 651218 542414 651454
rect 541794 651134 542414 651218
rect 541794 650898 541826 651134
rect 542062 650898 542146 651134
rect 542382 650898 542414 651134
rect 273168 619174 273488 619206
rect 273168 618938 273210 619174
rect 273446 618938 273488 619174
rect 273168 618854 273488 618938
rect 273168 618618 273210 618854
rect 273446 618618 273488 618854
rect 273168 618586 273488 618618
rect 303888 619174 304208 619206
rect 303888 618938 303930 619174
rect 304166 618938 304208 619174
rect 303888 618854 304208 618938
rect 303888 618618 303930 618854
rect 304166 618618 304208 618854
rect 303888 618586 304208 618618
rect 334608 619174 334928 619206
rect 334608 618938 334650 619174
rect 334886 618938 334928 619174
rect 334608 618854 334928 618938
rect 334608 618618 334650 618854
rect 334886 618618 334928 618854
rect 334608 618586 334928 618618
rect 365328 619174 365648 619206
rect 365328 618938 365370 619174
rect 365606 618938 365648 619174
rect 365328 618854 365648 618938
rect 365328 618618 365370 618854
rect 365606 618618 365648 618854
rect 365328 618586 365648 618618
rect 396048 619174 396368 619206
rect 396048 618938 396090 619174
rect 396326 618938 396368 619174
rect 396048 618854 396368 618938
rect 396048 618618 396090 618854
rect 396326 618618 396368 618854
rect 396048 618586 396368 618618
rect 426768 619174 427088 619206
rect 426768 618938 426810 619174
rect 427046 618938 427088 619174
rect 426768 618854 427088 618938
rect 426768 618618 426810 618854
rect 427046 618618 427088 618854
rect 426768 618586 427088 618618
rect 457488 619174 457808 619206
rect 457488 618938 457530 619174
rect 457766 618938 457808 619174
rect 457488 618854 457808 618938
rect 457488 618618 457530 618854
rect 457766 618618 457808 618854
rect 457488 618586 457808 618618
rect 488208 619174 488528 619206
rect 488208 618938 488250 619174
rect 488486 618938 488528 619174
rect 488208 618854 488528 618938
rect 488208 618618 488250 618854
rect 488486 618618 488528 618854
rect 488208 618586 488528 618618
rect 518928 619174 519248 619206
rect 518928 618938 518970 619174
rect 519206 618938 519248 619174
rect 518928 618854 519248 618938
rect 518928 618618 518970 618854
rect 519206 618618 519248 618854
rect 518928 618586 519248 618618
rect 253794 615218 253826 615454
rect 254062 615218 254146 615454
rect 254382 615218 254414 615454
rect 253794 615134 254414 615218
rect 253794 614898 253826 615134
rect 254062 614898 254146 615134
rect 254382 614898 254414 615134
rect 253794 579454 254414 614898
rect 257808 615454 258128 615486
rect 257808 615218 257850 615454
rect 258086 615218 258128 615454
rect 257808 615134 258128 615218
rect 257808 614898 257850 615134
rect 258086 614898 258128 615134
rect 257808 614866 258128 614898
rect 288528 615454 288848 615486
rect 288528 615218 288570 615454
rect 288806 615218 288848 615454
rect 288528 615134 288848 615218
rect 288528 614898 288570 615134
rect 288806 614898 288848 615134
rect 288528 614866 288848 614898
rect 319248 615454 319568 615486
rect 319248 615218 319290 615454
rect 319526 615218 319568 615454
rect 319248 615134 319568 615218
rect 319248 614898 319290 615134
rect 319526 614898 319568 615134
rect 319248 614866 319568 614898
rect 349968 615454 350288 615486
rect 349968 615218 350010 615454
rect 350246 615218 350288 615454
rect 349968 615134 350288 615218
rect 349968 614898 350010 615134
rect 350246 614898 350288 615134
rect 349968 614866 350288 614898
rect 380688 615454 381008 615486
rect 380688 615218 380730 615454
rect 380966 615218 381008 615454
rect 380688 615134 381008 615218
rect 380688 614898 380730 615134
rect 380966 614898 381008 615134
rect 380688 614866 381008 614898
rect 411408 615454 411728 615486
rect 411408 615218 411450 615454
rect 411686 615218 411728 615454
rect 411408 615134 411728 615218
rect 411408 614898 411450 615134
rect 411686 614898 411728 615134
rect 411408 614866 411728 614898
rect 442128 615454 442448 615486
rect 442128 615218 442170 615454
rect 442406 615218 442448 615454
rect 442128 615134 442448 615218
rect 442128 614898 442170 615134
rect 442406 614898 442448 615134
rect 442128 614866 442448 614898
rect 472848 615454 473168 615486
rect 472848 615218 472890 615454
rect 473126 615218 473168 615454
rect 472848 615134 473168 615218
rect 472848 614898 472890 615134
rect 473126 614898 473168 615134
rect 472848 614866 473168 614898
rect 503568 615454 503888 615486
rect 503568 615218 503610 615454
rect 503846 615218 503888 615454
rect 503568 615134 503888 615218
rect 503568 614898 503610 615134
rect 503846 614898 503888 615134
rect 503568 614866 503888 614898
rect 534288 615454 534608 615486
rect 534288 615218 534330 615454
rect 534566 615218 534608 615454
rect 534288 615134 534608 615218
rect 534288 614898 534330 615134
rect 534566 614898 534608 615134
rect 534288 614866 534608 614898
rect 541794 615454 542414 650898
rect 541794 615218 541826 615454
rect 542062 615218 542146 615454
rect 542382 615218 542414 615454
rect 541794 615134 542414 615218
rect 541794 614898 541826 615134
rect 542062 614898 542146 615134
rect 542382 614898 542414 615134
rect 273168 583174 273488 583206
rect 273168 582938 273210 583174
rect 273446 582938 273488 583174
rect 273168 582854 273488 582938
rect 273168 582618 273210 582854
rect 273446 582618 273488 582854
rect 273168 582586 273488 582618
rect 303888 583174 304208 583206
rect 303888 582938 303930 583174
rect 304166 582938 304208 583174
rect 303888 582854 304208 582938
rect 303888 582618 303930 582854
rect 304166 582618 304208 582854
rect 303888 582586 304208 582618
rect 334608 583174 334928 583206
rect 334608 582938 334650 583174
rect 334886 582938 334928 583174
rect 334608 582854 334928 582938
rect 334608 582618 334650 582854
rect 334886 582618 334928 582854
rect 334608 582586 334928 582618
rect 365328 583174 365648 583206
rect 365328 582938 365370 583174
rect 365606 582938 365648 583174
rect 365328 582854 365648 582938
rect 365328 582618 365370 582854
rect 365606 582618 365648 582854
rect 365328 582586 365648 582618
rect 396048 583174 396368 583206
rect 396048 582938 396090 583174
rect 396326 582938 396368 583174
rect 396048 582854 396368 582938
rect 396048 582618 396090 582854
rect 396326 582618 396368 582854
rect 396048 582586 396368 582618
rect 426768 583174 427088 583206
rect 426768 582938 426810 583174
rect 427046 582938 427088 583174
rect 426768 582854 427088 582938
rect 426768 582618 426810 582854
rect 427046 582618 427088 582854
rect 426768 582586 427088 582618
rect 457488 583174 457808 583206
rect 457488 582938 457530 583174
rect 457766 582938 457808 583174
rect 457488 582854 457808 582938
rect 457488 582618 457530 582854
rect 457766 582618 457808 582854
rect 457488 582586 457808 582618
rect 488208 583174 488528 583206
rect 488208 582938 488250 583174
rect 488486 582938 488528 583174
rect 488208 582854 488528 582938
rect 488208 582618 488250 582854
rect 488486 582618 488528 582854
rect 488208 582586 488528 582618
rect 518928 583174 519248 583206
rect 518928 582938 518970 583174
rect 519206 582938 519248 583174
rect 518928 582854 519248 582938
rect 518928 582618 518970 582854
rect 519206 582618 519248 582854
rect 518928 582586 519248 582618
rect 253794 579218 253826 579454
rect 254062 579218 254146 579454
rect 254382 579218 254414 579454
rect 253794 579134 254414 579218
rect 253794 578898 253826 579134
rect 254062 578898 254146 579134
rect 254382 578898 254414 579134
rect 253794 543454 254414 578898
rect 257808 579454 258128 579486
rect 257808 579218 257850 579454
rect 258086 579218 258128 579454
rect 257808 579134 258128 579218
rect 257808 578898 257850 579134
rect 258086 578898 258128 579134
rect 257808 578866 258128 578898
rect 288528 579454 288848 579486
rect 288528 579218 288570 579454
rect 288806 579218 288848 579454
rect 288528 579134 288848 579218
rect 288528 578898 288570 579134
rect 288806 578898 288848 579134
rect 288528 578866 288848 578898
rect 319248 579454 319568 579486
rect 319248 579218 319290 579454
rect 319526 579218 319568 579454
rect 319248 579134 319568 579218
rect 319248 578898 319290 579134
rect 319526 578898 319568 579134
rect 319248 578866 319568 578898
rect 349968 579454 350288 579486
rect 349968 579218 350010 579454
rect 350246 579218 350288 579454
rect 349968 579134 350288 579218
rect 349968 578898 350010 579134
rect 350246 578898 350288 579134
rect 349968 578866 350288 578898
rect 380688 579454 381008 579486
rect 380688 579218 380730 579454
rect 380966 579218 381008 579454
rect 380688 579134 381008 579218
rect 380688 578898 380730 579134
rect 380966 578898 381008 579134
rect 380688 578866 381008 578898
rect 411408 579454 411728 579486
rect 411408 579218 411450 579454
rect 411686 579218 411728 579454
rect 411408 579134 411728 579218
rect 411408 578898 411450 579134
rect 411686 578898 411728 579134
rect 411408 578866 411728 578898
rect 442128 579454 442448 579486
rect 442128 579218 442170 579454
rect 442406 579218 442448 579454
rect 442128 579134 442448 579218
rect 442128 578898 442170 579134
rect 442406 578898 442448 579134
rect 442128 578866 442448 578898
rect 472848 579454 473168 579486
rect 472848 579218 472890 579454
rect 473126 579218 473168 579454
rect 472848 579134 473168 579218
rect 472848 578898 472890 579134
rect 473126 578898 473168 579134
rect 472848 578866 473168 578898
rect 503568 579454 503888 579486
rect 503568 579218 503610 579454
rect 503846 579218 503888 579454
rect 503568 579134 503888 579218
rect 503568 578898 503610 579134
rect 503846 578898 503888 579134
rect 503568 578866 503888 578898
rect 534288 579454 534608 579486
rect 534288 579218 534330 579454
rect 534566 579218 534608 579454
rect 534288 579134 534608 579218
rect 534288 578898 534330 579134
rect 534566 578898 534608 579134
rect 534288 578866 534608 578898
rect 541794 579454 542414 614898
rect 541794 579218 541826 579454
rect 542062 579218 542146 579454
rect 542382 579218 542414 579454
rect 541794 579134 542414 579218
rect 541794 578898 541826 579134
rect 542062 578898 542146 579134
rect 542382 578898 542414 579134
rect 273168 547174 273488 547206
rect 273168 546938 273210 547174
rect 273446 546938 273488 547174
rect 273168 546854 273488 546938
rect 273168 546618 273210 546854
rect 273446 546618 273488 546854
rect 273168 546586 273488 546618
rect 303888 547174 304208 547206
rect 303888 546938 303930 547174
rect 304166 546938 304208 547174
rect 303888 546854 304208 546938
rect 303888 546618 303930 546854
rect 304166 546618 304208 546854
rect 303888 546586 304208 546618
rect 334608 547174 334928 547206
rect 334608 546938 334650 547174
rect 334886 546938 334928 547174
rect 334608 546854 334928 546938
rect 334608 546618 334650 546854
rect 334886 546618 334928 546854
rect 334608 546586 334928 546618
rect 365328 547174 365648 547206
rect 365328 546938 365370 547174
rect 365606 546938 365648 547174
rect 365328 546854 365648 546938
rect 365328 546618 365370 546854
rect 365606 546618 365648 546854
rect 365328 546586 365648 546618
rect 396048 547174 396368 547206
rect 396048 546938 396090 547174
rect 396326 546938 396368 547174
rect 396048 546854 396368 546938
rect 396048 546618 396090 546854
rect 396326 546618 396368 546854
rect 396048 546586 396368 546618
rect 426768 547174 427088 547206
rect 426768 546938 426810 547174
rect 427046 546938 427088 547174
rect 426768 546854 427088 546938
rect 426768 546618 426810 546854
rect 427046 546618 427088 546854
rect 426768 546586 427088 546618
rect 457488 547174 457808 547206
rect 457488 546938 457530 547174
rect 457766 546938 457808 547174
rect 457488 546854 457808 546938
rect 457488 546618 457530 546854
rect 457766 546618 457808 546854
rect 457488 546586 457808 546618
rect 488208 547174 488528 547206
rect 488208 546938 488250 547174
rect 488486 546938 488528 547174
rect 488208 546854 488528 546938
rect 488208 546618 488250 546854
rect 488486 546618 488528 546854
rect 488208 546586 488528 546618
rect 518928 547174 519248 547206
rect 518928 546938 518970 547174
rect 519206 546938 519248 547174
rect 518928 546854 519248 546938
rect 518928 546618 518970 546854
rect 519206 546618 519248 546854
rect 518928 546586 519248 546618
rect 253794 543218 253826 543454
rect 254062 543218 254146 543454
rect 254382 543218 254414 543454
rect 253794 543134 254414 543218
rect 253794 542898 253826 543134
rect 254062 542898 254146 543134
rect 254382 542898 254414 543134
rect 253794 507454 254414 542898
rect 257808 543454 258128 543486
rect 257808 543218 257850 543454
rect 258086 543218 258128 543454
rect 257808 543134 258128 543218
rect 257808 542898 257850 543134
rect 258086 542898 258128 543134
rect 257808 542866 258128 542898
rect 288528 543454 288848 543486
rect 288528 543218 288570 543454
rect 288806 543218 288848 543454
rect 288528 543134 288848 543218
rect 288528 542898 288570 543134
rect 288806 542898 288848 543134
rect 288528 542866 288848 542898
rect 319248 543454 319568 543486
rect 319248 543218 319290 543454
rect 319526 543218 319568 543454
rect 319248 543134 319568 543218
rect 319248 542898 319290 543134
rect 319526 542898 319568 543134
rect 319248 542866 319568 542898
rect 349968 543454 350288 543486
rect 349968 543218 350010 543454
rect 350246 543218 350288 543454
rect 349968 543134 350288 543218
rect 349968 542898 350010 543134
rect 350246 542898 350288 543134
rect 349968 542866 350288 542898
rect 380688 543454 381008 543486
rect 380688 543218 380730 543454
rect 380966 543218 381008 543454
rect 380688 543134 381008 543218
rect 380688 542898 380730 543134
rect 380966 542898 381008 543134
rect 380688 542866 381008 542898
rect 411408 543454 411728 543486
rect 411408 543218 411450 543454
rect 411686 543218 411728 543454
rect 411408 543134 411728 543218
rect 411408 542898 411450 543134
rect 411686 542898 411728 543134
rect 411408 542866 411728 542898
rect 442128 543454 442448 543486
rect 442128 543218 442170 543454
rect 442406 543218 442448 543454
rect 442128 543134 442448 543218
rect 442128 542898 442170 543134
rect 442406 542898 442448 543134
rect 442128 542866 442448 542898
rect 472848 543454 473168 543486
rect 472848 543218 472890 543454
rect 473126 543218 473168 543454
rect 472848 543134 473168 543218
rect 472848 542898 472890 543134
rect 473126 542898 473168 543134
rect 472848 542866 473168 542898
rect 503568 543454 503888 543486
rect 503568 543218 503610 543454
rect 503846 543218 503888 543454
rect 503568 543134 503888 543218
rect 503568 542898 503610 543134
rect 503846 542898 503888 543134
rect 503568 542866 503888 542898
rect 534288 543454 534608 543486
rect 534288 543218 534330 543454
rect 534566 543218 534608 543454
rect 534288 543134 534608 543218
rect 534288 542898 534330 543134
rect 534566 542898 534608 543134
rect 534288 542866 534608 542898
rect 541794 543454 542414 578898
rect 541794 543218 541826 543454
rect 542062 543218 542146 543454
rect 542382 543218 542414 543454
rect 541794 543134 542414 543218
rect 541794 542898 541826 543134
rect 542062 542898 542146 543134
rect 542382 542898 542414 543134
rect 253794 507218 253826 507454
rect 254062 507218 254146 507454
rect 254382 507218 254414 507454
rect 253794 507134 254414 507218
rect 253794 506898 253826 507134
rect 254062 506898 254146 507134
rect 254382 506898 254414 507134
rect 253794 471454 254414 506898
rect 276114 529774 276734 530431
rect 276114 529538 276146 529774
rect 276382 529538 276466 529774
rect 276702 529538 276734 529774
rect 276114 529454 276734 529538
rect 276114 529218 276146 529454
rect 276382 529218 276466 529454
rect 276702 529218 276734 529454
rect 276114 498713 276734 529218
rect 312114 529774 312734 530431
rect 312114 529538 312146 529774
rect 312382 529538 312466 529774
rect 312702 529538 312734 529774
rect 312114 529454 312734 529538
rect 312114 529218 312146 529454
rect 312382 529218 312466 529454
rect 312702 529218 312734 529454
rect 312114 498713 312734 529218
rect 348114 529774 348734 530431
rect 348114 529538 348146 529774
rect 348382 529538 348466 529774
rect 348702 529538 348734 529774
rect 348114 529454 348734 529538
rect 348114 529218 348146 529454
rect 348382 529218 348466 529454
rect 348702 529218 348734 529454
rect 348114 498713 348734 529218
rect 384114 529774 384734 530431
rect 384114 529538 384146 529774
rect 384382 529538 384466 529774
rect 384702 529538 384734 529774
rect 384114 529454 384734 529538
rect 384114 529218 384146 529454
rect 384382 529218 384466 529454
rect 384702 529218 384734 529454
rect 384114 498713 384734 529218
rect 420114 529774 420734 530431
rect 420114 529538 420146 529774
rect 420382 529538 420466 529774
rect 420702 529538 420734 529774
rect 420114 529454 420734 529538
rect 420114 529218 420146 529454
rect 420382 529218 420466 529454
rect 420702 529218 420734 529454
rect 420114 498713 420734 529218
rect 456114 529774 456734 530431
rect 456114 529538 456146 529774
rect 456382 529538 456466 529774
rect 456702 529538 456734 529774
rect 456114 529454 456734 529538
rect 456114 529218 456146 529454
rect 456382 529218 456466 529454
rect 456702 529218 456734 529454
rect 456114 498713 456734 529218
rect 492114 529774 492734 530431
rect 492114 529538 492146 529774
rect 492382 529538 492466 529774
rect 492702 529538 492734 529774
rect 492114 529454 492734 529538
rect 492114 529218 492146 529454
rect 492382 529218 492466 529454
rect 492702 529218 492734 529454
rect 492114 498713 492734 529218
rect 528114 529774 528734 530431
rect 528114 529538 528146 529774
rect 528382 529538 528466 529774
rect 528702 529538 528734 529774
rect 528114 529454 528734 529538
rect 528114 529218 528146 529454
rect 528382 529218 528466 529454
rect 528702 529218 528734 529454
rect 528114 498713 528734 529218
rect 541794 507454 542414 542898
rect 541794 507218 541826 507454
rect 542062 507218 542146 507454
rect 542382 507218 542414 507454
rect 541794 507134 542414 507218
rect 541794 506898 541826 507134
rect 542062 506898 542146 507134
rect 542382 506898 542414 507134
rect 273168 475174 273488 475206
rect 273168 474938 273210 475174
rect 273446 474938 273488 475174
rect 273168 474854 273488 474938
rect 273168 474618 273210 474854
rect 273446 474618 273488 474854
rect 273168 474586 273488 474618
rect 303888 475174 304208 475206
rect 303888 474938 303930 475174
rect 304166 474938 304208 475174
rect 303888 474854 304208 474938
rect 303888 474618 303930 474854
rect 304166 474618 304208 474854
rect 303888 474586 304208 474618
rect 334608 475174 334928 475206
rect 334608 474938 334650 475174
rect 334886 474938 334928 475174
rect 334608 474854 334928 474938
rect 334608 474618 334650 474854
rect 334886 474618 334928 474854
rect 334608 474586 334928 474618
rect 365328 475174 365648 475206
rect 365328 474938 365370 475174
rect 365606 474938 365648 475174
rect 365328 474854 365648 474938
rect 365328 474618 365370 474854
rect 365606 474618 365648 474854
rect 365328 474586 365648 474618
rect 396048 475174 396368 475206
rect 396048 474938 396090 475174
rect 396326 474938 396368 475174
rect 396048 474854 396368 474938
rect 396048 474618 396090 474854
rect 396326 474618 396368 474854
rect 396048 474586 396368 474618
rect 426768 475174 427088 475206
rect 426768 474938 426810 475174
rect 427046 474938 427088 475174
rect 426768 474854 427088 474938
rect 426768 474618 426810 474854
rect 427046 474618 427088 474854
rect 426768 474586 427088 474618
rect 457488 475174 457808 475206
rect 457488 474938 457530 475174
rect 457766 474938 457808 475174
rect 457488 474854 457808 474938
rect 457488 474618 457530 474854
rect 457766 474618 457808 474854
rect 457488 474586 457808 474618
rect 488208 475174 488528 475206
rect 488208 474938 488250 475174
rect 488486 474938 488528 475174
rect 488208 474854 488528 474938
rect 488208 474618 488250 474854
rect 488486 474618 488528 474854
rect 488208 474586 488528 474618
rect 518928 475174 519248 475206
rect 518928 474938 518970 475174
rect 519206 474938 519248 475174
rect 518928 474854 519248 474938
rect 518928 474618 518970 474854
rect 519206 474618 519248 474854
rect 518928 474586 519248 474618
rect 253794 471218 253826 471454
rect 254062 471218 254146 471454
rect 254382 471218 254414 471454
rect 253794 471134 254414 471218
rect 253794 470898 253826 471134
rect 254062 470898 254146 471134
rect 254382 470898 254414 471134
rect 253794 435454 254414 470898
rect 257808 471454 258128 471486
rect 257808 471218 257850 471454
rect 258086 471218 258128 471454
rect 257808 471134 258128 471218
rect 257808 470898 257850 471134
rect 258086 470898 258128 471134
rect 257808 470866 258128 470898
rect 288528 471454 288848 471486
rect 288528 471218 288570 471454
rect 288806 471218 288848 471454
rect 288528 471134 288848 471218
rect 288528 470898 288570 471134
rect 288806 470898 288848 471134
rect 288528 470866 288848 470898
rect 319248 471454 319568 471486
rect 319248 471218 319290 471454
rect 319526 471218 319568 471454
rect 319248 471134 319568 471218
rect 319248 470898 319290 471134
rect 319526 470898 319568 471134
rect 319248 470866 319568 470898
rect 349968 471454 350288 471486
rect 349968 471218 350010 471454
rect 350246 471218 350288 471454
rect 349968 471134 350288 471218
rect 349968 470898 350010 471134
rect 350246 470898 350288 471134
rect 349968 470866 350288 470898
rect 380688 471454 381008 471486
rect 380688 471218 380730 471454
rect 380966 471218 381008 471454
rect 380688 471134 381008 471218
rect 380688 470898 380730 471134
rect 380966 470898 381008 471134
rect 380688 470866 381008 470898
rect 411408 471454 411728 471486
rect 411408 471218 411450 471454
rect 411686 471218 411728 471454
rect 411408 471134 411728 471218
rect 411408 470898 411450 471134
rect 411686 470898 411728 471134
rect 411408 470866 411728 470898
rect 442128 471454 442448 471486
rect 442128 471218 442170 471454
rect 442406 471218 442448 471454
rect 442128 471134 442448 471218
rect 442128 470898 442170 471134
rect 442406 470898 442448 471134
rect 442128 470866 442448 470898
rect 472848 471454 473168 471486
rect 472848 471218 472890 471454
rect 473126 471218 473168 471454
rect 472848 471134 473168 471218
rect 472848 470898 472890 471134
rect 473126 470898 473168 471134
rect 472848 470866 473168 470898
rect 503568 471454 503888 471486
rect 503568 471218 503610 471454
rect 503846 471218 503888 471454
rect 503568 471134 503888 471218
rect 503568 470898 503610 471134
rect 503846 470898 503888 471134
rect 503568 470866 503888 470898
rect 534288 471454 534608 471486
rect 534288 471218 534330 471454
rect 534566 471218 534608 471454
rect 534288 471134 534608 471218
rect 534288 470898 534330 471134
rect 534566 470898 534608 471134
rect 534288 470866 534608 470898
rect 541794 471454 542414 506898
rect 541794 471218 541826 471454
rect 542062 471218 542146 471454
rect 542382 471218 542414 471454
rect 541794 471134 542414 471218
rect 541794 470898 541826 471134
rect 542062 470898 542146 471134
rect 542382 470898 542414 471134
rect 273168 439174 273488 439206
rect 273168 438938 273210 439174
rect 273446 438938 273488 439174
rect 273168 438854 273488 438938
rect 273168 438618 273210 438854
rect 273446 438618 273488 438854
rect 273168 438586 273488 438618
rect 303888 439174 304208 439206
rect 303888 438938 303930 439174
rect 304166 438938 304208 439174
rect 303888 438854 304208 438938
rect 303888 438618 303930 438854
rect 304166 438618 304208 438854
rect 303888 438586 304208 438618
rect 334608 439174 334928 439206
rect 334608 438938 334650 439174
rect 334886 438938 334928 439174
rect 334608 438854 334928 438938
rect 334608 438618 334650 438854
rect 334886 438618 334928 438854
rect 334608 438586 334928 438618
rect 365328 439174 365648 439206
rect 365328 438938 365370 439174
rect 365606 438938 365648 439174
rect 365328 438854 365648 438938
rect 365328 438618 365370 438854
rect 365606 438618 365648 438854
rect 365328 438586 365648 438618
rect 396048 439174 396368 439206
rect 396048 438938 396090 439174
rect 396326 438938 396368 439174
rect 396048 438854 396368 438938
rect 396048 438618 396090 438854
rect 396326 438618 396368 438854
rect 396048 438586 396368 438618
rect 426768 439174 427088 439206
rect 426768 438938 426810 439174
rect 427046 438938 427088 439174
rect 426768 438854 427088 438938
rect 426768 438618 426810 438854
rect 427046 438618 427088 438854
rect 426768 438586 427088 438618
rect 457488 439174 457808 439206
rect 457488 438938 457530 439174
rect 457766 438938 457808 439174
rect 457488 438854 457808 438938
rect 457488 438618 457530 438854
rect 457766 438618 457808 438854
rect 457488 438586 457808 438618
rect 488208 439174 488528 439206
rect 488208 438938 488250 439174
rect 488486 438938 488528 439174
rect 488208 438854 488528 438938
rect 488208 438618 488250 438854
rect 488486 438618 488528 438854
rect 488208 438586 488528 438618
rect 518928 439174 519248 439206
rect 518928 438938 518970 439174
rect 519206 438938 519248 439174
rect 518928 438854 519248 438938
rect 518928 438618 518970 438854
rect 519206 438618 519248 438854
rect 518928 438586 519248 438618
rect 253794 435218 253826 435454
rect 254062 435218 254146 435454
rect 254382 435218 254414 435454
rect 253794 435134 254414 435218
rect 253794 434898 253826 435134
rect 254062 434898 254146 435134
rect 254382 434898 254414 435134
rect 253794 399454 254414 434898
rect 257808 435454 258128 435486
rect 257808 435218 257850 435454
rect 258086 435218 258128 435454
rect 257808 435134 258128 435218
rect 257808 434898 257850 435134
rect 258086 434898 258128 435134
rect 257808 434866 258128 434898
rect 288528 435454 288848 435486
rect 288528 435218 288570 435454
rect 288806 435218 288848 435454
rect 288528 435134 288848 435218
rect 288528 434898 288570 435134
rect 288806 434898 288848 435134
rect 288528 434866 288848 434898
rect 319248 435454 319568 435486
rect 319248 435218 319290 435454
rect 319526 435218 319568 435454
rect 319248 435134 319568 435218
rect 319248 434898 319290 435134
rect 319526 434898 319568 435134
rect 319248 434866 319568 434898
rect 349968 435454 350288 435486
rect 349968 435218 350010 435454
rect 350246 435218 350288 435454
rect 349968 435134 350288 435218
rect 349968 434898 350010 435134
rect 350246 434898 350288 435134
rect 349968 434866 350288 434898
rect 380688 435454 381008 435486
rect 380688 435218 380730 435454
rect 380966 435218 381008 435454
rect 380688 435134 381008 435218
rect 380688 434898 380730 435134
rect 380966 434898 381008 435134
rect 380688 434866 381008 434898
rect 411408 435454 411728 435486
rect 411408 435218 411450 435454
rect 411686 435218 411728 435454
rect 411408 435134 411728 435218
rect 411408 434898 411450 435134
rect 411686 434898 411728 435134
rect 411408 434866 411728 434898
rect 442128 435454 442448 435486
rect 442128 435218 442170 435454
rect 442406 435218 442448 435454
rect 442128 435134 442448 435218
rect 442128 434898 442170 435134
rect 442406 434898 442448 435134
rect 442128 434866 442448 434898
rect 472848 435454 473168 435486
rect 472848 435218 472890 435454
rect 473126 435218 473168 435454
rect 472848 435134 473168 435218
rect 472848 434898 472890 435134
rect 473126 434898 473168 435134
rect 472848 434866 473168 434898
rect 503568 435454 503888 435486
rect 503568 435218 503610 435454
rect 503846 435218 503888 435454
rect 503568 435134 503888 435218
rect 503568 434898 503610 435134
rect 503846 434898 503888 435134
rect 503568 434866 503888 434898
rect 534288 435454 534608 435486
rect 534288 435218 534330 435454
rect 534566 435218 534608 435454
rect 534288 435134 534608 435218
rect 534288 434898 534330 435134
rect 534566 434898 534608 435134
rect 534288 434866 534608 434898
rect 541794 435454 542414 470898
rect 541794 435218 541826 435454
rect 542062 435218 542146 435454
rect 542382 435218 542414 435454
rect 541794 435134 542414 435218
rect 541794 434898 541826 435134
rect 542062 434898 542146 435134
rect 542382 434898 542414 435134
rect 273168 403174 273488 403206
rect 273168 402938 273210 403174
rect 273446 402938 273488 403174
rect 273168 402854 273488 402938
rect 273168 402618 273210 402854
rect 273446 402618 273488 402854
rect 273168 402586 273488 402618
rect 303888 403174 304208 403206
rect 303888 402938 303930 403174
rect 304166 402938 304208 403174
rect 303888 402854 304208 402938
rect 303888 402618 303930 402854
rect 304166 402618 304208 402854
rect 303888 402586 304208 402618
rect 334608 403174 334928 403206
rect 334608 402938 334650 403174
rect 334886 402938 334928 403174
rect 334608 402854 334928 402938
rect 334608 402618 334650 402854
rect 334886 402618 334928 402854
rect 334608 402586 334928 402618
rect 365328 403174 365648 403206
rect 365328 402938 365370 403174
rect 365606 402938 365648 403174
rect 365328 402854 365648 402938
rect 365328 402618 365370 402854
rect 365606 402618 365648 402854
rect 365328 402586 365648 402618
rect 396048 403174 396368 403206
rect 396048 402938 396090 403174
rect 396326 402938 396368 403174
rect 396048 402854 396368 402938
rect 396048 402618 396090 402854
rect 396326 402618 396368 402854
rect 396048 402586 396368 402618
rect 426768 403174 427088 403206
rect 426768 402938 426810 403174
rect 427046 402938 427088 403174
rect 426768 402854 427088 402938
rect 426768 402618 426810 402854
rect 427046 402618 427088 402854
rect 426768 402586 427088 402618
rect 457488 403174 457808 403206
rect 457488 402938 457530 403174
rect 457766 402938 457808 403174
rect 457488 402854 457808 402938
rect 457488 402618 457530 402854
rect 457766 402618 457808 402854
rect 457488 402586 457808 402618
rect 488208 403174 488528 403206
rect 488208 402938 488250 403174
rect 488486 402938 488528 403174
rect 488208 402854 488528 402938
rect 488208 402618 488250 402854
rect 488486 402618 488528 402854
rect 488208 402586 488528 402618
rect 518928 403174 519248 403206
rect 518928 402938 518970 403174
rect 519206 402938 519248 403174
rect 518928 402854 519248 402938
rect 518928 402618 518970 402854
rect 519206 402618 519248 402854
rect 518928 402586 519248 402618
rect 253794 399218 253826 399454
rect 254062 399218 254146 399454
rect 254382 399218 254414 399454
rect 253794 399134 254414 399218
rect 253794 398898 253826 399134
rect 254062 398898 254146 399134
rect 254382 398898 254414 399134
rect 253794 363454 254414 398898
rect 257808 399454 258128 399486
rect 257808 399218 257850 399454
rect 258086 399218 258128 399454
rect 257808 399134 258128 399218
rect 257808 398898 257850 399134
rect 258086 398898 258128 399134
rect 257808 398866 258128 398898
rect 288528 399454 288848 399486
rect 288528 399218 288570 399454
rect 288806 399218 288848 399454
rect 288528 399134 288848 399218
rect 288528 398898 288570 399134
rect 288806 398898 288848 399134
rect 288528 398866 288848 398898
rect 319248 399454 319568 399486
rect 319248 399218 319290 399454
rect 319526 399218 319568 399454
rect 319248 399134 319568 399218
rect 319248 398898 319290 399134
rect 319526 398898 319568 399134
rect 319248 398866 319568 398898
rect 349968 399454 350288 399486
rect 349968 399218 350010 399454
rect 350246 399218 350288 399454
rect 349968 399134 350288 399218
rect 349968 398898 350010 399134
rect 350246 398898 350288 399134
rect 349968 398866 350288 398898
rect 380688 399454 381008 399486
rect 380688 399218 380730 399454
rect 380966 399218 381008 399454
rect 380688 399134 381008 399218
rect 380688 398898 380730 399134
rect 380966 398898 381008 399134
rect 380688 398866 381008 398898
rect 411408 399454 411728 399486
rect 411408 399218 411450 399454
rect 411686 399218 411728 399454
rect 411408 399134 411728 399218
rect 411408 398898 411450 399134
rect 411686 398898 411728 399134
rect 411408 398866 411728 398898
rect 442128 399454 442448 399486
rect 442128 399218 442170 399454
rect 442406 399218 442448 399454
rect 442128 399134 442448 399218
rect 442128 398898 442170 399134
rect 442406 398898 442448 399134
rect 442128 398866 442448 398898
rect 472848 399454 473168 399486
rect 472848 399218 472890 399454
rect 473126 399218 473168 399454
rect 472848 399134 473168 399218
rect 472848 398898 472890 399134
rect 473126 398898 473168 399134
rect 472848 398866 473168 398898
rect 503568 399454 503888 399486
rect 503568 399218 503610 399454
rect 503846 399218 503888 399454
rect 503568 399134 503888 399218
rect 503568 398898 503610 399134
rect 503846 398898 503888 399134
rect 503568 398866 503888 398898
rect 534288 399454 534608 399486
rect 534288 399218 534330 399454
rect 534566 399218 534608 399454
rect 534288 399134 534608 399218
rect 534288 398898 534330 399134
rect 534566 398898 534608 399134
rect 534288 398866 534608 398898
rect 541794 399454 542414 434898
rect 541794 399218 541826 399454
rect 542062 399218 542146 399454
rect 542382 399218 542414 399454
rect 541794 399134 542414 399218
rect 541794 398898 541826 399134
rect 542062 398898 542146 399134
rect 542382 398898 542414 399134
rect 253794 363218 253826 363454
rect 254062 363218 254146 363454
rect 254382 363218 254414 363454
rect 253794 363134 254414 363218
rect 253794 362898 253826 363134
rect 254062 362898 254146 363134
rect 254382 362898 254414 363134
rect 253794 327454 254414 362898
rect 253794 327218 253826 327454
rect 254062 327218 254146 327454
rect 254382 327218 254414 327454
rect 253794 327134 254414 327218
rect 253794 326898 253826 327134
rect 254062 326898 254146 327134
rect 254382 326898 254414 327134
rect 253794 291454 254414 326898
rect 253794 291218 253826 291454
rect 254062 291218 254146 291454
rect 254382 291218 254414 291454
rect 253794 291134 254414 291218
rect 253794 290898 253826 291134
rect 254062 290898 254146 291134
rect 254382 290898 254414 291134
rect 253794 255454 254414 290898
rect 253794 255218 253826 255454
rect 254062 255218 254146 255454
rect 254382 255218 254414 255454
rect 253794 255134 254414 255218
rect 253794 254898 253826 255134
rect 254062 254898 254146 255134
rect 254382 254898 254414 255134
rect 253794 219454 254414 254898
rect 253794 219218 253826 219454
rect 254062 219218 254146 219454
rect 254382 219218 254414 219454
rect 253794 219134 254414 219218
rect 253794 218898 253826 219134
rect 254062 218898 254146 219134
rect 254382 218898 254414 219134
rect 253794 183454 254414 218898
rect 253794 183218 253826 183454
rect 254062 183218 254146 183454
rect 254382 183218 254414 183454
rect 253794 183134 254414 183218
rect 253794 182898 253826 183134
rect 254062 182898 254146 183134
rect 254382 182898 254414 183134
rect 253794 147454 254414 182898
rect 253794 147218 253826 147454
rect 254062 147218 254146 147454
rect 254382 147218 254414 147454
rect 253794 147134 254414 147218
rect 253794 146898 253826 147134
rect 254062 146898 254146 147134
rect 254382 146898 254414 147134
rect 253794 111454 254414 146898
rect 253794 111218 253826 111454
rect 254062 111218 254146 111454
rect 254382 111218 254414 111454
rect 253794 111134 254414 111218
rect 253794 110898 253826 111134
rect 254062 110898 254146 111134
rect 254382 110898 254414 111134
rect 253794 75454 254414 110898
rect 253794 75218 253826 75454
rect 254062 75218 254146 75454
rect 254382 75218 254414 75454
rect 253794 75134 254414 75218
rect 253794 74898 253826 75134
rect 254062 74898 254146 75134
rect 254382 74898 254414 75134
rect 251771 52732 251837 52733
rect 251771 52668 251772 52732
rect 251836 52668 251837 52732
rect 251771 52667 251837 52668
rect 243834 29258 243866 29494
rect 244102 29258 244186 29494
rect 244422 29258 244454 29494
rect 243834 29174 244454 29258
rect 243834 28938 243866 29174
rect 244102 28938 244186 29174
rect 244422 28938 244454 29174
rect 243834 -7066 244454 28938
rect 243834 -7302 243866 -7066
rect 244102 -7302 244186 -7066
rect 244422 -7302 244454 -7066
rect 243834 -7386 244454 -7302
rect 243834 -7622 243866 -7386
rect 244102 -7622 244186 -7386
rect 244422 -7622 244454 -7386
rect 243834 -7654 244454 -7622
rect 253794 39454 254414 74898
rect 253794 39218 253826 39454
rect 254062 39218 254146 39454
rect 254382 39218 254414 39454
rect 253794 39134 254414 39218
rect 253794 38898 253826 39134
rect 254062 38898 254146 39134
rect 254382 38898 254414 39134
rect 253794 3454 254414 38898
rect 253794 3218 253826 3454
rect 254062 3218 254146 3454
rect 254382 3218 254414 3454
rect 253794 3134 254414 3218
rect 253794 2898 253826 3134
rect 254062 2898 254146 3134
rect 254382 2898 254414 3134
rect 253794 -346 254414 2898
rect 253794 -582 253826 -346
rect 254062 -582 254146 -346
rect 254382 -582 254414 -346
rect 253794 -666 254414 -582
rect 253794 -902 253826 -666
rect 254062 -902 254146 -666
rect 254382 -902 254414 -666
rect 253794 -7654 254414 -902
rect 257514 367174 258134 380068
rect 257514 366938 257546 367174
rect 257782 366938 257866 367174
rect 258102 366938 258134 367174
rect 257514 366854 258134 366938
rect 257514 366618 257546 366854
rect 257782 366618 257866 366854
rect 258102 366618 258134 366854
rect 257514 331174 258134 366618
rect 257514 330938 257546 331174
rect 257782 330938 257866 331174
rect 258102 330938 258134 331174
rect 257514 330854 258134 330938
rect 257514 330618 257546 330854
rect 257782 330618 257866 330854
rect 258102 330618 258134 330854
rect 257514 295174 258134 330618
rect 261234 370894 261854 380831
rect 261234 370658 261266 370894
rect 261502 370658 261586 370894
rect 261822 370658 261854 370894
rect 261234 370574 261854 370658
rect 261234 370338 261266 370574
rect 261502 370338 261586 370574
rect 261822 370338 261854 370574
rect 261234 334894 261854 370338
rect 261234 334658 261266 334894
rect 261502 334658 261586 334894
rect 261822 334658 261854 334894
rect 261234 334574 261854 334658
rect 261234 334338 261266 334574
rect 261502 334338 261586 334574
rect 261822 334338 261854 334574
rect 261234 320417 261854 334338
rect 264954 374614 265574 380831
rect 264954 374378 264986 374614
rect 265222 374378 265306 374614
rect 265542 374378 265574 374614
rect 264954 374294 265574 374378
rect 264954 374058 264986 374294
rect 265222 374058 265306 374294
rect 265542 374058 265574 374294
rect 264954 338614 265574 374058
rect 264954 338378 264986 338614
rect 265222 338378 265306 338614
rect 265542 338378 265574 338614
rect 264954 338294 265574 338378
rect 264954 338058 264986 338294
rect 265222 338058 265306 338294
rect 265542 338058 265574 338294
rect 264954 320417 265574 338058
rect 268674 378334 269294 380831
rect 268674 378098 268706 378334
rect 268942 378098 269026 378334
rect 269262 378098 269294 378334
rect 268674 378014 269294 378098
rect 268674 377778 268706 378014
rect 268942 377778 269026 378014
rect 269262 377778 269294 378014
rect 268674 342334 269294 377778
rect 268674 342098 268706 342334
rect 268942 342098 269026 342334
rect 269262 342098 269294 342334
rect 268674 342014 269294 342098
rect 268674 341778 268706 342014
rect 268942 341778 269026 342014
rect 269262 341778 269294 342014
rect 268674 320417 269294 341778
rect 289794 363454 290414 380831
rect 289794 363218 289826 363454
rect 290062 363218 290146 363454
rect 290382 363218 290414 363454
rect 289794 363134 290414 363218
rect 289794 362898 289826 363134
rect 290062 362898 290146 363134
rect 290382 362898 290414 363134
rect 289794 327454 290414 362898
rect 289794 327218 289826 327454
rect 290062 327218 290146 327454
rect 290382 327218 290414 327454
rect 289794 327134 290414 327218
rect 289794 326898 289826 327134
rect 290062 326898 290146 327134
rect 290382 326898 290414 327134
rect 289794 320417 290414 326898
rect 293514 367174 294134 380831
rect 293514 366938 293546 367174
rect 293782 366938 293866 367174
rect 294102 366938 294134 367174
rect 293514 366854 294134 366938
rect 293514 366618 293546 366854
rect 293782 366618 293866 366854
rect 294102 366618 294134 366854
rect 293514 331174 294134 366618
rect 293514 330938 293546 331174
rect 293782 330938 293866 331174
rect 294102 330938 294134 331174
rect 293514 330854 294134 330938
rect 293514 330618 293546 330854
rect 293782 330618 293866 330854
rect 294102 330618 294134 330854
rect 293514 320417 294134 330618
rect 297234 370894 297854 380831
rect 297234 370658 297266 370894
rect 297502 370658 297586 370894
rect 297822 370658 297854 370894
rect 297234 370574 297854 370658
rect 297234 370338 297266 370574
rect 297502 370338 297586 370574
rect 297822 370338 297854 370574
rect 297234 334894 297854 370338
rect 297234 334658 297266 334894
rect 297502 334658 297586 334894
rect 297822 334658 297854 334894
rect 297234 334574 297854 334658
rect 297234 334338 297266 334574
rect 297502 334338 297586 334574
rect 297822 334338 297854 334574
rect 297234 320417 297854 334338
rect 300954 374614 301574 380831
rect 300954 374378 300986 374614
rect 301222 374378 301306 374614
rect 301542 374378 301574 374614
rect 300954 374294 301574 374378
rect 300954 374058 300986 374294
rect 301222 374058 301306 374294
rect 301542 374058 301574 374294
rect 300954 338614 301574 374058
rect 300954 338378 300986 338614
rect 301222 338378 301306 338614
rect 301542 338378 301574 338614
rect 300954 338294 301574 338378
rect 300954 338058 300986 338294
rect 301222 338058 301306 338294
rect 301542 338058 301574 338294
rect 300954 320417 301574 338058
rect 304674 378334 305294 380831
rect 304674 378098 304706 378334
rect 304942 378098 305026 378334
rect 305262 378098 305294 378334
rect 304674 378014 305294 378098
rect 304674 377778 304706 378014
rect 304942 377778 305026 378014
rect 305262 377778 305294 378014
rect 304674 342334 305294 377778
rect 304674 342098 304706 342334
rect 304942 342098 305026 342334
rect 305262 342098 305294 342334
rect 304674 342014 305294 342098
rect 304674 341778 304706 342014
rect 304942 341778 305026 342014
rect 305262 341778 305294 342014
rect 304674 320417 305294 341778
rect 325794 363454 326414 380831
rect 325794 363218 325826 363454
rect 326062 363218 326146 363454
rect 326382 363218 326414 363454
rect 325794 363134 326414 363218
rect 325794 362898 325826 363134
rect 326062 362898 326146 363134
rect 326382 362898 326414 363134
rect 325794 327454 326414 362898
rect 325794 327218 325826 327454
rect 326062 327218 326146 327454
rect 326382 327218 326414 327454
rect 325794 327134 326414 327218
rect 325794 326898 325826 327134
rect 326062 326898 326146 327134
rect 326382 326898 326414 327134
rect 325794 320417 326414 326898
rect 329514 367174 330134 380831
rect 329514 366938 329546 367174
rect 329782 366938 329866 367174
rect 330102 366938 330134 367174
rect 329514 366854 330134 366938
rect 329514 366618 329546 366854
rect 329782 366618 329866 366854
rect 330102 366618 330134 366854
rect 329514 331174 330134 366618
rect 329514 330938 329546 331174
rect 329782 330938 329866 331174
rect 330102 330938 330134 331174
rect 329514 330854 330134 330938
rect 329514 330618 329546 330854
rect 329782 330618 329866 330854
rect 330102 330618 330134 330854
rect 329514 320417 330134 330618
rect 333234 370894 333854 380831
rect 333234 370658 333266 370894
rect 333502 370658 333586 370894
rect 333822 370658 333854 370894
rect 333234 370574 333854 370658
rect 333234 370338 333266 370574
rect 333502 370338 333586 370574
rect 333822 370338 333854 370574
rect 333234 334894 333854 370338
rect 333234 334658 333266 334894
rect 333502 334658 333586 334894
rect 333822 334658 333854 334894
rect 333234 334574 333854 334658
rect 333234 334338 333266 334574
rect 333502 334338 333586 334574
rect 333822 334338 333854 334574
rect 333234 320417 333854 334338
rect 336954 374614 337574 380831
rect 336954 374378 336986 374614
rect 337222 374378 337306 374614
rect 337542 374378 337574 374614
rect 336954 374294 337574 374378
rect 336954 374058 336986 374294
rect 337222 374058 337306 374294
rect 337542 374058 337574 374294
rect 336954 338614 337574 374058
rect 336954 338378 336986 338614
rect 337222 338378 337306 338614
rect 337542 338378 337574 338614
rect 336954 338294 337574 338378
rect 336954 338058 336986 338294
rect 337222 338058 337306 338294
rect 337542 338058 337574 338294
rect 336954 320417 337574 338058
rect 340674 378334 341294 380831
rect 340674 378098 340706 378334
rect 340942 378098 341026 378334
rect 341262 378098 341294 378334
rect 340674 378014 341294 378098
rect 340674 377778 340706 378014
rect 340942 377778 341026 378014
rect 341262 377778 341294 378014
rect 340674 342334 341294 377778
rect 340674 342098 340706 342334
rect 340942 342098 341026 342334
rect 341262 342098 341294 342334
rect 340674 342014 341294 342098
rect 340674 341778 340706 342014
rect 340942 341778 341026 342014
rect 341262 341778 341294 342014
rect 340674 320417 341294 341778
rect 361794 363454 362414 380831
rect 361794 363218 361826 363454
rect 362062 363218 362146 363454
rect 362382 363218 362414 363454
rect 361794 363134 362414 363218
rect 361794 362898 361826 363134
rect 362062 362898 362146 363134
rect 362382 362898 362414 363134
rect 361794 327454 362414 362898
rect 361794 327218 361826 327454
rect 362062 327218 362146 327454
rect 362382 327218 362414 327454
rect 361794 327134 362414 327218
rect 361794 326898 361826 327134
rect 362062 326898 362146 327134
rect 362382 326898 362414 327134
rect 361794 320417 362414 326898
rect 365514 367174 366134 380068
rect 365514 366938 365546 367174
rect 365782 366938 365866 367174
rect 366102 366938 366134 367174
rect 365514 366854 366134 366938
rect 365514 366618 365546 366854
rect 365782 366618 365866 366854
rect 366102 366618 366134 366854
rect 365514 331174 366134 366618
rect 365514 330938 365546 331174
rect 365782 330938 365866 331174
rect 366102 330938 366134 331174
rect 365514 330854 366134 330938
rect 365514 330618 365546 330854
rect 365782 330618 365866 330854
rect 366102 330618 366134 330854
rect 365514 320417 366134 330618
rect 369234 370894 369854 380831
rect 369234 370658 369266 370894
rect 369502 370658 369586 370894
rect 369822 370658 369854 370894
rect 369234 370574 369854 370658
rect 369234 370338 369266 370574
rect 369502 370338 369586 370574
rect 369822 370338 369854 370574
rect 369234 334894 369854 370338
rect 369234 334658 369266 334894
rect 369502 334658 369586 334894
rect 369822 334658 369854 334894
rect 369234 334574 369854 334658
rect 369234 334338 369266 334574
rect 369502 334338 369586 334574
rect 369822 334338 369854 334574
rect 369234 320417 369854 334338
rect 372954 374614 373574 380831
rect 372954 374378 372986 374614
rect 373222 374378 373306 374614
rect 373542 374378 373574 374614
rect 372954 374294 373574 374378
rect 372954 374058 372986 374294
rect 373222 374058 373306 374294
rect 373542 374058 373574 374294
rect 372954 338614 373574 374058
rect 372954 338378 372986 338614
rect 373222 338378 373306 338614
rect 373542 338378 373574 338614
rect 372954 338294 373574 338378
rect 372954 338058 372986 338294
rect 373222 338058 373306 338294
rect 373542 338058 373574 338294
rect 372954 320417 373574 338058
rect 376674 378334 377294 380831
rect 376674 378098 376706 378334
rect 376942 378098 377026 378334
rect 377262 378098 377294 378334
rect 376674 378014 377294 378098
rect 376674 377778 376706 378014
rect 376942 377778 377026 378014
rect 377262 377778 377294 378014
rect 376674 342334 377294 377778
rect 376674 342098 376706 342334
rect 376942 342098 377026 342334
rect 377262 342098 377294 342334
rect 376674 342014 377294 342098
rect 376674 341778 376706 342014
rect 376942 341778 377026 342014
rect 377262 341778 377294 342014
rect 376674 320417 377294 341778
rect 397794 363454 398414 380831
rect 397794 363218 397826 363454
rect 398062 363218 398146 363454
rect 398382 363218 398414 363454
rect 397794 363134 398414 363218
rect 397794 362898 397826 363134
rect 398062 362898 398146 363134
rect 398382 362898 398414 363134
rect 397794 327454 398414 362898
rect 397794 327218 397826 327454
rect 398062 327218 398146 327454
rect 398382 327218 398414 327454
rect 397794 327134 398414 327218
rect 397794 326898 397826 327134
rect 398062 326898 398146 327134
rect 398382 326898 398414 327134
rect 397794 320417 398414 326898
rect 401514 367174 402134 380831
rect 401514 366938 401546 367174
rect 401782 366938 401866 367174
rect 402102 366938 402134 367174
rect 401514 366854 402134 366938
rect 401514 366618 401546 366854
rect 401782 366618 401866 366854
rect 402102 366618 402134 366854
rect 401514 331174 402134 366618
rect 401514 330938 401546 331174
rect 401782 330938 401866 331174
rect 402102 330938 402134 331174
rect 401514 330854 402134 330938
rect 401514 330618 401546 330854
rect 401782 330618 401866 330854
rect 402102 330618 402134 330854
rect 401514 320417 402134 330618
rect 405234 370894 405854 380831
rect 405234 370658 405266 370894
rect 405502 370658 405586 370894
rect 405822 370658 405854 370894
rect 405234 370574 405854 370658
rect 405234 370338 405266 370574
rect 405502 370338 405586 370574
rect 405822 370338 405854 370574
rect 405234 334894 405854 370338
rect 405234 334658 405266 334894
rect 405502 334658 405586 334894
rect 405822 334658 405854 334894
rect 405234 334574 405854 334658
rect 405234 334338 405266 334574
rect 405502 334338 405586 334574
rect 405822 334338 405854 334574
rect 405234 320417 405854 334338
rect 408954 374614 409574 380831
rect 408954 374378 408986 374614
rect 409222 374378 409306 374614
rect 409542 374378 409574 374614
rect 408954 374294 409574 374378
rect 408954 374058 408986 374294
rect 409222 374058 409306 374294
rect 409542 374058 409574 374294
rect 408954 338614 409574 374058
rect 408954 338378 408986 338614
rect 409222 338378 409306 338614
rect 409542 338378 409574 338614
rect 408954 338294 409574 338378
rect 408954 338058 408986 338294
rect 409222 338058 409306 338294
rect 409542 338058 409574 338294
rect 408954 320417 409574 338058
rect 412674 378334 413294 380831
rect 412674 378098 412706 378334
rect 412942 378098 413026 378334
rect 413262 378098 413294 378334
rect 412674 378014 413294 378098
rect 412674 377778 412706 378014
rect 412942 377778 413026 378014
rect 413262 377778 413294 378014
rect 412674 342334 413294 377778
rect 412674 342098 412706 342334
rect 412942 342098 413026 342334
rect 413262 342098 413294 342334
rect 412674 342014 413294 342098
rect 412674 341778 412706 342014
rect 412942 341778 413026 342014
rect 413262 341778 413294 342014
rect 412674 320417 413294 341778
rect 433794 363454 434414 380831
rect 433794 363218 433826 363454
rect 434062 363218 434146 363454
rect 434382 363218 434414 363454
rect 433794 363134 434414 363218
rect 433794 362898 433826 363134
rect 434062 362898 434146 363134
rect 434382 362898 434414 363134
rect 433794 327454 434414 362898
rect 433794 327218 433826 327454
rect 434062 327218 434146 327454
rect 434382 327218 434414 327454
rect 433794 327134 434414 327218
rect 433794 326898 433826 327134
rect 434062 326898 434146 327134
rect 434382 326898 434414 327134
rect 433794 320417 434414 326898
rect 437514 367174 438134 380831
rect 437514 366938 437546 367174
rect 437782 366938 437866 367174
rect 438102 366938 438134 367174
rect 437514 366854 438134 366938
rect 437514 366618 437546 366854
rect 437782 366618 437866 366854
rect 438102 366618 438134 366854
rect 437514 331174 438134 366618
rect 437514 330938 437546 331174
rect 437782 330938 437866 331174
rect 438102 330938 438134 331174
rect 437514 330854 438134 330938
rect 437514 330618 437546 330854
rect 437782 330618 437866 330854
rect 438102 330618 438134 330854
rect 437514 320417 438134 330618
rect 441234 370894 441854 380831
rect 441234 370658 441266 370894
rect 441502 370658 441586 370894
rect 441822 370658 441854 370894
rect 441234 370574 441854 370658
rect 441234 370338 441266 370574
rect 441502 370338 441586 370574
rect 441822 370338 441854 370574
rect 441234 334894 441854 370338
rect 441234 334658 441266 334894
rect 441502 334658 441586 334894
rect 441822 334658 441854 334894
rect 441234 334574 441854 334658
rect 441234 334338 441266 334574
rect 441502 334338 441586 334574
rect 441822 334338 441854 334574
rect 441234 320417 441854 334338
rect 444954 374614 445574 380831
rect 444954 374378 444986 374614
rect 445222 374378 445306 374614
rect 445542 374378 445574 374614
rect 444954 374294 445574 374378
rect 444954 374058 444986 374294
rect 445222 374058 445306 374294
rect 445542 374058 445574 374294
rect 444954 338614 445574 374058
rect 444954 338378 444986 338614
rect 445222 338378 445306 338614
rect 445542 338378 445574 338614
rect 444954 338294 445574 338378
rect 444954 338058 444986 338294
rect 445222 338058 445306 338294
rect 445542 338058 445574 338294
rect 444954 320417 445574 338058
rect 448674 378334 449294 380831
rect 448674 378098 448706 378334
rect 448942 378098 449026 378334
rect 449262 378098 449294 378334
rect 448674 378014 449294 378098
rect 448674 377778 448706 378014
rect 448942 377778 449026 378014
rect 449262 377778 449294 378014
rect 448674 342334 449294 377778
rect 448674 342098 448706 342334
rect 448942 342098 449026 342334
rect 449262 342098 449294 342334
rect 448674 342014 449294 342098
rect 448674 341778 448706 342014
rect 448942 341778 449026 342014
rect 449262 341778 449294 342014
rect 448674 320417 449294 341778
rect 469794 363454 470414 380831
rect 469794 363218 469826 363454
rect 470062 363218 470146 363454
rect 470382 363218 470414 363454
rect 469794 363134 470414 363218
rect 469794 362898 469826 363134
rect 470062 362898 470146 363134
rect 470382 362898 470414 363134
rect 469794 327454 470414 362898
rect 469794 327218 469826 327454
rect 470062 327218 470146 327454
rect 470382 327218 470414 327454
rect 469794 327134 470414 327218
rect 469794 326898 469826 327134
rect 470062 326898 470146 327134
rect 470382 326898 470414 327134
rect 469794 320417 470414 326898
rect 473514 367174 474134 380831
rect 473514 366938 473546 367174
rect 473782 366938 473866 367174
rect 474102 366938 474134 367174
rect 473514 366854 474134 366938
rect 473514 366618 473546 366854
rect 473782 366618 473866 366854
rect 474102 366618 474134 366854
rect 473514 331174 474134 366618
rect 473514 330938 473546 331174
rect 473782 330938 473866 331174
rect 474102 330938 474134 331174
rect 473514 330854 474134 330938
rect 473514 330618 473546 330854
rect 473782 330618 473866 330854
rect 474102 330618 474134 330854
rect 473514 320417 474134 330618
rect 477234 370894 477854 380831
rect 477234 370658 477266 370894
rect 477502 370658 477586 370894
rect 477822 370658 477854 370894
rect 477234 370574 477854 370658
rect 477234 370338 477266 370574
rect 477502 370338 477586 370574
rect 477822 370338 477854 370574
rect 477234 334894 477854 370338
rect 477234 334658 477266 334894
rect 477502 334658 477586 334894
rect 477822 334658 477854 334894
rect 477234 334574 477854 334658
rect 477234 334338 477266 334574
rect 477502 334338 477586 334574
rect 477822 334338 477854 334574
rect 477234 320417 477854 334338
rect 480954 374614 481574 380831
rect 480954 374378 480986 374614
rect 481222 374378 481306 374614
rect 481542 374378 481574 374614
rect 480954 374294 481574 374378
rect 480954 374058 480986 374294
rect 481222 374058 481306 374294
rect 481542 374058 481574 374294
rect 480954 338614 481574 374058
rect 480954 338378 480986 338614
rect 481222 338378 481306 338614
rect 481542 338378 481574 338614
rect 480954 338294 481574 338378
rect 480954 338058 480986 338294
rect 481222 338058 481306 338294
rect 481542 338058 481574 338294
rect 480954 320417 481574 338058
rect 484674 378334 485294 380831
rect 484674 378098 484706 378334
rect 484942 378098 485026 378334
rect 485262 378098 485294 378334
rect 484674 378014 485294 378098
rect 484674 377778 484706 378014
rect 484942 377778 485026 378014
rect 485262 377778 485294 378014
rect 484674 342334 485294 377778
rect 484674 342098 484706 342334
rect 484942 342098 485026 342334
rect 485262 342098 485294 342334
rect 484674 342014 485294 342098
rect 484674 341778 484706 342014
rect 484942 341778 485026 342014
rect 485262 341778 485294 342014
rect 484674 320417 485294 341778
rect 505794 363454 506414 380831
rect 505794 363218 505826 363454
rect 506062 363218 506146 363454
rect 506382 363218 506414 363454
rect 505794 363134 506414 363218
rect 505794 362898 505826 363134
rect 506062 362898 506146 363134
rect 506382 362898 506414 363134
rect 505794 327454 506414 362898
rect 505794 327218 505826 327454
rect 506062 327218 506146 327454
rect 506382 327218 506414 327454
rect 505794 327134 506414 327218
rect 505794 326898 505826 327134
rect 506062 326898 506146 327134
rect 506382 326898 506414 327134
rect 505794 320417 506414 326898
rect 509514 367174 510134 380831
rect 509514 366938 509546 367174
rect 509782 366938 509866 367174
rect 510102 366938 510134 367174
rect 509514 366854 510134 366938
rect 509514 366618 509546 366854
rect 509782 366618 509866 366854
rect 510102 366618 510134 366854
rect 509514 331174 510134 366618
rect 509514 330938 509546 331174
rect 509782 330938 509866 331174
rect 510102 330938 510134 331174
rect 509514 330854 510134 330938
rect 509514 330618 509546 330854
rect 509782 330618 509866 330854
rect 510102 330618 510134 330854
rect 509514 320417 510134 330618
rect 513234 370894 513854 380831
rect 513234 370658 513266 370894
rect 513502 370658 513586 370894
rect 513822 370658 513854 370894
rect 513234 370574 513854 370658
rect 513234 370338 513266 370574
rect 513502 370338 513586 370574
rect 513822 370338 513854 370574
rect 513234 334894 513854 370338
rect 513234 334658 513266 334894
rect 513502 334658 513586 334894
rect 513822 334658 513854 334894
rect 513234 334574 513854 334658
rect 513234 334338 513266 334574
rect 513502 334338 513586 334574
rect 513822 334338 513854 334574
rect 513234 320417 513854 334338
rect 516954 374614 517574 380831
rect 516954 374378 516986 374614
rect 517222 374378 517306 374614
rect 517542 374378 517574 374614
rect 516954 374294 517574 374378
rect 516954 374058 516986 374294
rect 517222 374058 517306 374294
rect 517542 374058 517574 374294
rect 516954 338614 517574 374058
rect 516954 338378 516986 338614
rect 517222 338378 517306 338614
rect 517542 338378 517574 338614
rect 516954 338294 517574 338378
rect 516954 338058 516986 338294
rect 517222 338058 517306 338294
rect 517542 338058 517574 338294
rect 516954 320417 517574 338058
rect 520674 378334 521294 380831
rect 520674 378098 520706 378334
rect 520942 378098 521026 378334
rect 521262 378098 521294 378334
rect 520674 378014 521294 378098
rect 520674 377778 520706 378014
rect 520942 377778 521026 378014
rect 521262 377778 521294 378014
rect 520674 342334 521294 377778
rect 520674 342098 520706 342334
rect 520942 342098 521026 342334
rect 521262 342098 521294 342334
rect 520674 342014 521294 342098
rect 520674 341778 520706 342014
rect 520942 341778 521026 342014
rect 521262 341778 521294 342014
rect 520674 320417 521294 341778
rect 541794 363454 542414 398898
rect 541794 363218 541826 363454
rect 542062 363218 542146 363454
rect 542382 363218 542414 363454
rect 541794 363134 542414 363218
rect 541794 362898 541826 363134
rect 542062 362898 542146 363134
rect 542382 362898 542414 363134
rect 541794 327454 542414 362898
rect 541794 327218 541826 327454
rect 542062 327218 542146 327454
rect 542382 327218 542414 327454
rect 541794 327134 542414 327218
rect 541794 326898 541826 327134
rect 542062 326898 542146 327134
rect 542382 326898 542414 327134
rect 541794 320417 542414 326898
rect 545514 705798 546134 711590
rect 545514 705562 545546 705798
rect 545782 705562 545866 705798
rect 546102 705562 546134 705798
rect 545514 705478 546134 705562
rect 545514 705242 545546 705478
rect 545782 705242 545866 705478
rect 546102 705242 546134 705478
rect 545514 691174 546134 705242
rect 545514 690938 545546 691174
rect 545782 690938 545866 691174
rect 546102 690938 546134 691174
rect 545514 690854 546134 690938
rect 545514 690618 545546 690854
rect 545782 690618 545866 690854
rect 546102 690618 546134 690854
rect 545514 655174 546134 690618
rect 545514 654938 545546 655174
rect 545782 654938 545866 655174
rect 546102 654938 546134 655174
rect 545514 654854 546134 654938
rect 545514 654618 545546 654854
rect 545782 654618 545866 654854
rect 546102 654618 546134 654854
rect 545514 619174 546134 654618
rect 549234 706758 549854 711590
rect 549234 706522 549266 706758
rect 549502 706522 549586 706758
rect 549822 706522 549854 706758
rect 549234 706438 549854 706522
rect 549234 706202 549266 706438
rect 549502 706202 549586 706438
rect 549822 706202 549854 706438
rect 549234 694894 549854 706202
rect 549234 694658 549266 694894
rect 549502 694658 549586 694894
rect 549822 694658 549854 694894
rect 549234 694574 549854 694658
rect 549234 694338 549266 694574
rect 549502 694338 549586 694574
rect 549822 694338 549854 694574
rect 549234 658894 549854 694338
rect 549234 658658 549266 658894
rect 549502 658658 549586 658894
rect 549822 658658 549854 658894
rect 549234 658574 549854 658658
rect 549234 658338 549266 658574
rect 549502 658338 549586 658574
rect 549822 658338 549854 658574
rect 549234 649212 549854 658338
rect 552954 707718 553574 711590
rect 552954 707482 552986 707718
rect 553222 707482 553306 707718
rect 553542 707482 553574 707718
rect 552954 707398 553574 707482
rect 552954 707162 552986 707398
rect 553222 707162 553306 707398
rect 553542 707162 553574 707398
rect 552954 698614 553574 707162
rect 552954 698378 552986 698614
rect 553222 698378 553306 698614
rect 553542 698378 553574 698614
rect 552954 698294 553574 698378
rect 552954 698058 552986 698294
rect 553222 698058 553306 698294
rect 553542 698058 553574 698294
rect 552954 662614 553574 698058
rect 552954 662378 552986 662614
rect 553222 662378 553306 662614
rect 553542 662378 553574 662614
rect 552954 662294 553574 662378
rect 552954 662058 552986 662294
rect 553222 662058 553306 662294
rect 553542 662058 553574 662294
rect 552954 626614 553574 662058
rect 552954 626378 552986 626614
rect 553222 626378 553306 626614
rect 553542 626378 553574 626614
rect 552954 626294 553574 626378
rect 552954 626058 552986 626294
rect 553222 626058 553306 626294
rect 553542 626058 553574 626294
rect 545514 618938 545546 619174
rect 545782 618938 545866 619174
rect 546102 618938 546134 619174
rect 545514 618854 546134 618938
rect 545514 618618 545546 618854
rect 545782 618618 545866 618854
rect 546102 618618 546134 618854
rect 545514 583174 546134 618618
rect 549648 619174 549968 619206
rect 549648 618938 549690 619174
rect 549926 618938 549968 619174
rect 549648 618854 549968 618938
rect 549648 618618 549690 618854
rect 549926 618618 549968 618854
rect 549648 618586 549968 618618
rect 552954 590614 553574 626058
rect 552954 590378 552986 590614
rect 553222 590378 553306 590614
rect 553542 590378 553574 590614
rect 552954 590294 553574 590378
rect 552954 590058 552986 590294
rect 553222 590058 553306 590294
rect 553542 590058 553574 590294
rect 545514 582938 545546 583174
rect 545782 582938 545866 583174
rect 546102 582938 546134 583174
rect 545514 582854 546134 582938
rect 545514 582618 545546 582854
rect 545782 582618 545866 582854
rect 546102 582618 546134 582854
rect 545514 547174 546134 582618
rect 549648 583174 549968 583206
rect 549648 582938 549690 583174
rect 549926 582938 549968 583174
rect 549648 582854 549968 582938
rect 549648 582618 549690 582854
rect 549926 582618 549968 582854
rect 549648 582586 549968 582618
rect 552954 554614 553574 590058
rect 552954 554378 552986 554614
rect 553222 554378 553306 554614
rect 553542 554378 553574 554614
rect 552954 554294 553574 554378
rect 552954 554058 552986 554294
rect 553222 554058 553306 554294
rect 553542 554058 553574 554294
rect 545514 546938 545546 547174
rect 545782 546938 545866 547174
rect 546102 546938 546134 547174
rect 545514 546854 546134 546938
rect 545514 546618 545546 546854
rect 545782 546618 545866 546854
rect 546102 546618 546134 546854
rect 545514 511174 546134 546618
rect 549648 547174 549968 547206
rect 549648 546938 549690 547174
rect 549926 546938 549968 547174
rect 549648 546854 549968 546938
rect 549648 546618 549690 546854
rect 549926 546618 549968 546854
rect 549648 546586 549968 546618
rect 545514 510938 545546 511174
rect 545782 510938 545866 511174
rect 546102 510938 546134 511174
rect 545514 510854 546134 510938
rect 545514 510618 545546 510854
rect 545782 510618 545866 510854
rect 546102 510618 546134 510854
rect 545514 475174 546134 510618
rect 552954 518614 553574 554058
rect 552954 518378 552986 518614
rect 553222 518378 553306 518614
rect 553542 518378 553574 518614
rect 552954 518294 553574 518378
rect 552954 518058 552986 518294
rect 553222 518058 553306 518294
rect 553542 518058 553574 518294
rect 552954 482614 553574 518058
rect 552954 482378 552986 482614
rect 553222 482378 553306 482614
rect 553542 482378 553574 482614
rect 552954 482294 553574 482378
rect 552954 482058 552986 482294
rect 553222 482058 553306 482294
rect 553542 482058 553574 482294
rect 545514 474938 545546 475174
rect 545782 474938 545866 475174
rect 546102 474938 546134 475174
rect 545514 474854 546134 474938
rect 545514 474618 545546 474854
rect 545782 474618 545866 474854
rect 546102 474618 546134 474854
rect 545514 439174 546134 474618
rect 549648 475174 549968 475206
rect 549648 474938 549690 475174
rect 549926 474938 549968 475174
rect 549648 474854 549968 474938
rect 549648 474618 549690 474854
rect 549926 474618 549968 474854
rect 549648 474586 549968 474618
rect 552954 446614 553574 482058
rect 552954 446378 552986 446614
rect 553222 446378 553306 446614
rect 553542 446378 553574 446614
rect 552954 446294 553574 446378
rect 552954 446058 552986 446294
rect 553222 446058 553306 446294
rect 553542 446058 553574 446294
rect 545514 438938 545546 439174
rect 545782 438938 545866 439174
rect 546102 438938 546134 439174
rect 545514 438854 546134 438938
rect 545514 438618 545546 438854
rect 545782 438618 545866 438854
rect 546102 438618 546134 438854
rect 545514 403174 546134 438618
rect 549648 439174 549968 439206
rect 549648 438938 549690 439174
rect 549926 438938 549968 439174
rect 549648 438854 549968 438938
rect 549648 438618 549690 438854
rect 549926 438618 549968 438854
rect 549648 438586 549968 438618
rect 552954 410614 553574 446058
rect 552954 410378 552986 410614
rect 553222 410378 553306 410614
rect 553542 410378 553574 410614
rect 552954 410294 553574 410378
rect 552954 410058 552986 410294
rect 553222 410058 553306 410294
rect 553542 410058 553574 410294
rect 545514 402938 545546 403174
rect 545782 402938 545866 403174
rect 546102 402938 546134 403174
rect 545514 402854 546134 402938
rect 545514 402618 545546 402854
rect 545782 402618 545866 402854
rect 546102 402618 546134 402854
rect 545514 367174 546134 402618
rect 549648 403174 549968 403206
rect 549648 402938 549690 403174
rect 549926 402938 549968 403174
rect 549648 402854 549968 402938
rect 549648 402618 549690 402854
rect 549926 402618 549968 402854
rect 549648 402586 549968 402618
rect 545514 366938 545546 367174
rect 545782 366938 545866 367174
rect 546102 366938 546134 367174
rect 545514 366854 546134 366938
rect 545514 366618 545546 366854
rect 545782 366618 545866 366854
rect 546102 366618 546134 366854
rect 545514 331174 546134 366618
rect 545514 330938 545546 331174
rect 545782 330938 545866 331174
rect 546102 330938 546134 331174
rect 545514 330854 546134 330938
rect 545514 330618 545546 330854
rect 545782 330618 545866 330854
rect 546102 330618 546134 330854
rect 545514 320417 546134 330618
rect 549234 370894 549854 380068
rect 549234 370658 549266 370894
rect 549502 370658 549586 370894
rect 549822 370658 549854 370894
rect 549234 370574 549854 370658
rect 549234 370338 549266 370574
rect 549502 370338 549586 370574
rect 549822 370338 549854 370574
rect 549234 334894 549854 370338
rect 549234 334658 549266 334894
rect 549502 334658 549586 334894
rect 549822 334658 549854 334894
rect 549234 334574 549854 334658
rect 549234 334338 549266 334574
rect 549502 334338 549586 334574
rect 549822 334338 549854 334574
rect 549234 320417 549854 334338
rect 552954 374614 553574 410058
rect 552954 374378 552986 374614
rect 553222 374378 553306 374614
rect 553542 374378 553574 374614
rect 552954 374294 553574 374378
rect 552954 374058 552986 374294
rect 553222 374058 553306 374294
rect 553542 374058 553574 374294
rect 552954 338614 553574 374058
rect 552954 338378 552986 338614
rect 553222 338378 553306 338614
rect 553542 338378 553574 338614
rect 552954 338294 553574 338378
rect 552954 338058 552986 338294
rect 553222 338058 553306 338294
rect 553542 338058 553574 338294
rect 552954 302614 553574 338058
rect 552954 302378 552986 302614
rect 553222 302378 553306 302614
rect 553542 302378 553574 302614
rect 552954 302294 553574 302378
rect 552954 302058 552986 302294
rect 553222 302058 553306 302294
rect 553542 302058 553574 302294
rect 257514 294938 257546 295174
rect 257782 294938 257866 295174
rect 258102 294938 258134 295174
rect 257514 294854 258134 294938
rect 257514 294618 257546 294854
rect 257782 294618 257866 294854
rect 258102 294618 258134 294854
rect 257514 259174 258134 294618
rect 279568 295174 279888 295206
rect 279568 294938 279610 295174
rect 279846 294938 279888 295174
rect 279568 294854 279888 294938
rect 279568 294618 279610 294854
rect 279846 294618 279888 294854
rect 279568 294586 279888 294618
rect 310288 295174 310608 295206
rect 310288 294938 310330 295174
rect 310566 294938 310608 295174
rect 310288 294854 310608 294938
rect 310288 294618 310330 294854
rect 310566 294618 310608 294854
rect 310288 294586 310608 294618
rect 341008 295174 341328 295206
rect 341008 294938 341050 295174
rect 341286 294938 341328 295174
rect 341008 294854 341328 294938
rect 341008 294618 341050 294854
rect 341286 294618 341328 294854
rect 341008 294586 341328 294618
rect 371728 295174 372048 295206
rect 371728 294938 371770 295174
rect 372006 294938 372048 295174
rect 371728 294854 372048 294938
rect 371728 294618 371770 294854
rect 372006 294618 372048 294854
rect 371728 294586 372048 294618
rect 402448 295174 402768 295206
rect 402448 294938 402490 295174
rect 402726 294938 402768 295174
rect 402448 294854 402768 294938
rect 402448 294618 402490 294854
rect 402726 294618 402768 294854
rect 402448 294586 402768 294618
rect 433168 295174 433488 295206
rect 433168 294938 433210 295174
rect 433446 294938 433488 295174
rect 433168 294854 433488 294938
rect 433168 294618 433210 294854
rect 433446 294618 433488 294854
rect 433168 294586 433488 294618
rect 463888 295174 464208 295206
rect 463888 294938 463930 295174
rect 464166 294938 464208 295174
rect 463888 294854 464208 294938
rect 463888 294618 463930 294854
rect 464166 294618 464208 294854
rect 463888 294586 464208 294618
rect 494608 295174 494928 295206
rect 494608 294938 494650 295174
rect 494886 294938 494928 295174
rect 494608 294854 494928 294938
rect 494608 294618 494650 294854
rect 494886 294618 494928 294854
rect 494608 294586 494928 294618
rect 525328 295174 525648 295206
rect 525328 294938 525370 295174
rect 525606 294938 525648 295174
rect 525328 294854 525648 294938
rect 525328 294618 525370 294854
rect 525606 294618 525648 294854
rect 525328 294586 525648 294618
rect 264208 291454 264528 291486
rect 264208 291218 264250 291454
rect 264486 291218 264528 291454
rect 264208 291134 264528 291218
rect 264208 290898 264250 291134
rect 264486 290898 264528 291134
rect 264208 290866 264528 290898
rect 294928 291454 295248 291486
rect 294928 291218 294970 291454
rect 295206 291218 295248 291454
rect 294928 291134 295248 291218
rect 294928 290898 294970 291134
rect 295206 290898 295248 291134
rect 294928 290866 295248 290898
rect 325648 291454 325968 291486
rect 325648 291218 325690 291454
rect 325926 291218 325968 291454
rect 325648 291134 325968 291218
rect 325648 290898 325690 291134
rect 325926 290898 325968 291134
rect 325648 290866 325968 290898
rect 356368 291454 356688 291486
rect 356368 291218 356410 291454
rect 356646 291218 356688 291454
rect 356368 291134 356688 291218
rect 356368 290898 356410 291134
rect 356646 290898 356688 291134
rect 356368 290866 356688 290898
rect 387088 291454 387408 291486
rect 387088 291218 387130 291454
rect 387366 291218 387408 291454
rect 387088 291134 387408 291218
rect 387088 290898 387130 291134
rect 387366 290898 387408 291134
rect 387088 290866 387408 290898
rect 417808 291454 418128 291486
rect 417808 291218 417850 291454
rect 418086 291218 418128 291454
rect 417808 291134 418128 291218
rect 417808 290898 417850 291134
rect 418086 290898 418128 291134
rect 417808 290866 418128 290898
rect 448528 291454 448848 291486
rect 448528 291218 448570 291454
rect 448806 291218 448848 291454
rect 448528 291134 448848 291218
rect 448528 290898 448570 291134
rect 448806 290898 448848 291134
rect 448528 290866 448848 290898
rect 479248 291454 479568 291486
rect 479248 291218 479290 291454
rect 479526 291218 479568 291454
rect 479248 291134 479568 291218
rect 479248 290898 479290 291134
rect 479526 290898 479568 291134
rect 479248 290866 479568 290898
rect 509968 291454 510288 291486
rect 509968 291218 510010 291454
rect 510246 291218 510288 291454
rect 509968 291134 510288 291218
rect 509968 290898 510010 291134
rect 510246 290898 510288 291134
rect 509968 290866 510288 290898
rect 540688 291454 541008 291486
rect 540688 291218 540730 291454
rect 540966 291218 541008 291454
rect 540688 291134 541008 291218
rect 540688 290898 540730 291134
rect 540966 290898 541008 291134
rect 540688 290866 541008 290898
rect 552954 266614 553574 302058
rect 552954 266378 552986 266614
rect 553222 266378 553306 266614
rect 553542 266378 553574 266614
rect 552954 266294 553574 266378
rect 552954 266058 552986 266294
rect 553222 266058 553306 266294
rect 553542 266058 553574 266294
rect 257514 258938 257546 259174
rect 257782 258938 257866 259174
rect 258102 258938 258134 259174
rect 257514 258854 258134 258938
rect 257514 258618 257546 258854
rect 257782 258618 257866 258854
rect 258102 258618 258134 258854
rect 257514 223174 258134 258618
rect 279568 259174 279888 259206
rect 279568 258938 279610 259174
rect 279846 258938 279888 259174
rect 279568 258854 279888 258938
rect 279568 258618 279610 258854
rect 279846 258618 279888 258854
rect 279568 258586 279888 258618
rect 310288 259174 310608 259206
rect 310288 258938 310330 259174
rect 310566 258938 310608 259174
rect 310288 258854 310608 258938
rect 310288 258618 310330 258854
rect 310566 258618 310608 258854
rect 310288 258586 310608 258618
rect 341008 259174 341328 259206
rect 341008 258938 341050 259174
rect 341286 258938 341328 259174
rect 341008 258854 341328 258938
rect 341008 258618 341050 258854
rect 341286 258618 341328 258854
rect 341008 258586 341328 258618
rect 371728 259174 372048 259206
rect 371728 258938 371770 259174
rect 372006 258938 372048 259174
rect 371728 258854 372048 258938
rect 371728 258618 371770 258854
rect 372006 258618 372048 258854
rect 371728 258586 372048 258618
rect 402448 259174 402768 259206
rect 402448 258938 402490 259174
rect 402726 258938 402768 259174
rect 402448 258854 402768 258938
rect 402448 258618 402490 258854
rect 402726 258618 402768 258854
rect 402448 258586 402768 258618
rect 433168 259174 433488 259206
rect 433168 258938 433210 259174
rect 433446 258938 433488 259174
rect 433168 258854 433488 258938
rect 433168 258618 433210 258854
rect 433446 258618 433488 258854
rect 433168 258586 433488 258618
rect 463888 259174 464208 259206
rect 463888 258938 463930 259174
rect 464166 258938 464208 259174
rect 463888 258854 464208 258938
rect 463888 258618 463930 258854
rect 464166 258618 464208 258854
rect 463888 258586 464208 258618
rect 494608 259174 494928 259206
rect 494608 258938 494650 259174
rect 494886 258938 494928 259174
rect 494608 258854 494928 258938
rect 494608 258618 494650 258854
rect 494886 258618 494928 258854
rect 494608 258586 494928 258618
rect 525328 259174 525648 259206
rect 525328 258938 525370 259174
rect 525606 258938 525648 259174
rect 525328 258854 525648 258938
rect 525328 258618 525370 258854
rect 525606 258618 525648 258854
rect 525328 258586 525648 258618
rect 264208 255454 264528 255486
rect 264208 255218 264250 255454
rect 264486 255218 264528 255454
rect 264208 255134 264528 255218
rect 264208 254898 264250 255134
rect 264486 254898 264528 255134
rect 264208 254866 264528 254898
rect 294928 255454 295248 255486
rect 294928 255218 294970 255454
rect 295206 255218 295248 255454
rect 294928 255134 295248 255218
rect 294928 254898 294970 255134
rect 295206 254898 295248 255134
rect 294928 254866 295248 254898
rect 325648 255454 325968 255486
rect 325648 255218 325690 255454
rect 325926 255218 325968 255454
rect 325648 255134 325968 255218
rect 325648 254898 325690 255134
rect 325926 254898 325968 255134
rect 325648 254866 325968 254898
rect 356368 255454 356688 255486
rect 356368 255218 356410 255454
rect 356646 255218 356688 255454
rect 356368 255134 356688 255218
rect 356368 254898 356410 255134
rect 356646 254898 356688 255134
rect 356368 254866 356688 254898
rect 387088 255454 387408 255486
rect 387088 255218 387130 255454
rect 387366 255218 387408 255454
rect 387088 255134 387408 255218
rect 387088 254898 387130 255134
rect 387366 254898 387408 255134
rect 387088 254866 387408 254898
rect 417808 255454 418128 255486
rect 417808 255218 417850 255454
rect 418086 255218 418128 255454
rect 417808 255134 418128 255218
rect 417808 254898 417850 255134
rect 418086 254898 418128 255134
rect 417808 254866 418128 254898
rect 448528 255454 448848 255486
rect 448528 255218 448570 255454
rect 448806 255218 448848 255454
rect 448528 255134 448848 255218
rect 448528 254898 448570 255134
rect 448806 254898 448848 255134
rect 448528 254866 448848 254898
rect 479248 255454 479568 255486
rect 479248 255218 479290 255454
rect 479526 255218 479568 255454
rect 479248 255134 479568 255218
rect 479248 254898 479290 255134
rect 479526 254898 479568 255134
rect 479248 254866 479568 254898
rect 509968 255454 510288 255486
rect 509968 255218 510010 255454
rect 510246 255218 510288 255454
rect 509968 255134 510288 255218
rect 509968 254898 510010 255134
rect 510246 254898 510288 255134
rect 509968 254866 510288 254898
rect 540688 255454 541008 255486
rect 540688 255218 540730 255454
rect 540966 255218 541008 255454
rect 540688 255134 541008 255218
rect 540688 254898 540730 255134
rect 540966 254898 541008 255134
rect 540688 254866 541008 254898
rect 552954 230614 553574 266058
rect 552954 230378 552986 230614
rect 553222 230378 553306 230614
rect 553542 230378 553574 230614
rect 552954 230294 553574 230378
rect 552954 230058 552986 230294
rect 553222 230058 553306 230294
rect 553542 230058 553574 230294
rect 257514 222938 257546 223174
rect 257782 222938 257866 223174
rect 258102 222938 258134 223174
rect 257514 222854 258134 222938
rect 257514 222618 257546 222854
rect 257782 222618 257866 222854
rect 258102 222618 258134 222854
rect 257514 187174 258134 222618
rect 279568 223174 279888 223206
rect 279568 222938 279610 223174
rect 279846 222938 279888 223174
rect 279568 222854 279888 222938
rect 279568 222618 279610 222854
rect 279846 222618 279888 222854
rect 279568 222586 279888 222618
rect 310288 223174 310608 223206
rect 310288 222938 310330 223174
rect 310566 222938 310608 223174
rect 310288 222854 310608 222938
rect 310288 222618 310330 222854
rect 310566 222618 310608 222854
rect 310288 222586 310608 222618
rect 341008 223174 341328 223206
rect 341008 222938 341050 223174
rect 341286 222938 341328 223174
rect 341008 222854 341328 222938
rect 341008 222618 341050 222854
rect 341286 222618 341328 222854
rect 341008 222586 341328 222618
rect 371728 223174 372048 223206
rect 371728 222938 371770 223174
rect 372006 222938 372048 223174
rect 371728 222854 372048 222938
rect 371728 222618 371770 222854
rect 372006 222618 372048 222854
rect 371728 222586 372048 222618
rect 402448 223174 402768 223206
rect 402448 222938 402490 223174
rect 402726 222938 402768 223174
rect 402448 222854 402768 222938
rect 402448 222618 402490 222854
rect 402726 222618 402768 222854
rect 402448 222586 402768 222618
rect 433168 223174 433488 223206
rect 433168 222938 433210 223174
rect 433446 222938 433488 223174
rect 433168 222854 433488 222938
rect 433168 222618 433210 222854
rect 433446 222618 433488 222854
rect 433168 222586 433488 222618
rect 463888 223174 464208 223206
rect 463888 222938 463930 223174
rect 464166 222938 464208 223174
rect 463888 222854 464208 222938
rect 463888 222618 463930 222854
rect 464166 222618 464208 222854
rect 463888 222586 464208 222618
rect 494608 223174 494928 223206
rect 494608 222938 494650 223174
rect 494886 222938 494928 223174
rect 494608 222854 494928 222938
rect 494608 222618 494650 222854
rect 494886 222618 494928 222854
rect 494608 222586 494928 222618
rect 525328 223174 525648 223206
rect 525328 222938 525370 223174
rect 525606 222938 525648 223174
rect 525328 222854 525648 222938
rect 525328 222618 525370 222854
rect 525606 222618 525648 222854
rect 525328 222586 525648 222618
rect 264208 219454 264528 219486
rect 264208 219218 264250 219454
rect 264486 219218 264528 219454
rect 264208 219134 264528 219218
rect 264208 218898 264250 219134
rect 264486 218898 264528 219134
rect 264208 218866 264528 218898
rect 294928 219454 295248 219486
rect 294928 219218 294970 219454
rect 295206 219218 295248 219454
rect 294928 219134 295248 219218
rect 294928 218898 294970 219134
rect 295206 218898 295248 219134
rect 294928 218866 295248 218898
rect 325648 219454 325968 219486
rect 325648 219218 325690 219454
rect 325926 219218 325968 219454
rect 325648 219134 325968 219218
rect 325648 218898 325690 219134
rect 325926 218898 325968 219134
rect 325648 218866 325968 218898
rect 356368 219454 356688 219486
rect 356368 219218 356410 219454
rect 356646 219218 356688 219454
rect 356368 219134 356688 219218
rect 356368 218898 356410 219134
rect 356646 218898 356688 219134
rect 356368 218866 356688 218898
rect 387088 219454 387408 219486
rect 387088 219218 387130 219454
rect 387366 219218 387408 219454
rect 387088 219134 387408 219218
rect 387088 218898 387130 219134
rect 387366 218898 387408 219134
rect 387088 218866 387408 218898
rect 417808 219454 418128 219486
rect 417808 219218 417850 219454
rect 418086 219218 418128 219454
rect 417808 219134 418128 219218
rect 417808 218898 417850 219134
rect 418086 218898 418128 219134
rect 417808 218866 418128 218898
rect 448528 219454 448848 219486
rect 448528 219218 448570 219454
rect 448806 219218 448848 219454
rect 448528 219134 448848 219218
rect 448528 218898 448570 219134
rect 448806 218898 448848 219134
rect 448528 218866 448848 218898
rect 479248 219454 479568 219486
rect 479248 219218 479290 219454
rect 479526 219218 479568 219454
rect 479248 219134 479568 219218
rect 479248 218898 479290 219134
rect 479526 218898 479568 219134
rect 479248 218866 479568 218898
rect 509968 219454 510288 219486
rect 509968 219218 510010 219454
rect 510246 219218 510288 219454
rect 509968 219134 510288 219218
rect 509968 218898 510010 219134
rect 510246 218898 510288 219134
rect 509968 218866 510288 218898
rect 540688 219454 541008 219486
rect 540688 219218 540730 219454
rect 540966 219218 541008 219454
rect 540688 219134 541008 219218
rect 540688 218898 540730 219134
rect 540966 218898 541008 219134
rect 540688 218866 541008 218898
rect 552954 194614 553574 230058
rect 552954 194378 552986 194614
rect 553222 194378 553306 194614
rect 553542 194378 553574 194614
rect 552954 194294 553574 194378
rect 552954 194058 552986 194294
rect 553222 194058 553306 194294
rect 553542 194058 553574 194294
rect 257514 186938 257546 187174
rect 257782 186938 257866 187174
rect 258102 186938 258134 187174
rect 257514 186854 258134 186938
rect 257514 186618 257546 186854
rect 257782 186618 257866 186854
rect 258102 186618 258134 186854
rect 257514 151174 258134 186618
rect 279568 187174 279888 187206
rect 279568 186938 279610 187174
rect 279846 186938 279888 187174
rect 279568 186854 279888 186938
rect 279568 186618 279610 186854
rect 279846 186618 279888 186854
rect 279568 186586 279888 186618
rect 310288 187174 310608 187206
rect 310288 186938 310330 187174
rect 310566 186938 310608 187174
rect 310288 186854 310608 186938
rect 310288 186618 310330 186854
rect 310566 186618 310608 186854
rect 310288 186586 310608 186618
rect 341008 187174 341328 187206
rect 341008 186938 341050 187174
rect 341286 186938 341328 187174
rect 341008 186854 341328 186938
rect 341008 186618 341050 186854
rect 341286 186618 341328 186854
rect 341008 186586 341328 186618
rect 371728 187174 372048 187206
rect 371728 186938 371770 187174
rect 372006 186938 372048 187174
rect 371728 186854 372048 186938
rect 371728 186618 371770 186854
rect 372006 186618 372048 186854
rect 371728 186586 372048 186618
rect 402448 187174 402768 187206
rect 402448 186938 402490 187174
rect 402726 186938 402768 187174
rect 402448 186854 402768 186938
rect 402448 186618 402490 186854
rect 402726 186618 402768 186854
rect 402448 186586 402768 186618
rect 433168 187174 433488 187206
rect 433168 186938 433210 187174
rect 433446 186938 433488 187174
rect 433168 186854 433488 186938
rect 433168 186618 433210 186854
rect 433446 186618 433488 186854
rect 433168 186586 433488 186618
rect 463888 187174 464208 187206
rect 463888 186938 463930 187174
rect 464166 186938 464208 187174
rect 463888 186854 464208 186938
rect 463888 186618 463930 186854
rect 464166 186618 464208 186854
rect 463888 186586 464208 186618
rect 494608 187174 494928 187206
rect 494608 186938 494650 187174
rect 494886 186938 494928 187174
rect 494608 186854 494928 186938
rect 494608 186618 494650 186854
rect 494886 186618 494928 186854
rect 494608 186586 494928 186618
rect 525328 187174 525648 187206
rect 525328 186938 525370 187174
rect 525606 186938 525648 187174
rect 525328 186854 525648 186938
rect 525328 186618 525370 186854
rect 525606 186618 525648 186854
rect 525328 186586 525648 186618
rect 264208 183454 264528 183486
rect 264208 183218 264250 183454
rect 264486 183218 264528 183454
rect 264208 183134 264528 183218
rect 264208 182898 264250 183134
rect 264486 182898 264528 183134
rect 264208 182866 264528 182898
rect 294928 183454 295248 183486
rect 294928 183218 294970 183454
rect 295206 183218 295248 183454
rect 294928 183134 295248 183218
rect 294928 182898 294970 183134
rect 295206 182898 295248 183134
rect 294928 182866 295248 182898
rect 325648 183454 325968 183486
rect 325648 183218 325690 183454
rect 325926 183218 325968 183454
rect 325648 183134 325968 183218
rect 325648 182898 325690 183134
rect 325926 182898 325968 183134
rect 325648 182866 325968 182898
rect 356368 183454 356688 183486
rect 356368 183218 356410 183454
rect 356646 183218 356688 183454
rect 356368 183134 356688 183218
rect 356368 182898 356410 183134
rect 356646 182898 356688 183134
rect 356368 182866 356688 182898
rect 387088 183454 387408 183486
rect 387088 183218 387130 183454
rect 387366 183218 387408 183454
rect 387088 183134 387408 183218
rect 387088 182898 387130 183134
rect 387366 182898 387408 183134
rect 387088 182866 387408 182898
rect 417808 183454 418128 183486
rect 417808 183218 417850 183454
rect 418086 183218 418128 183454
rect 417808 183134 418128 183218
rect 417808 182898 417850 183134
rect 418086 182898 418128 183134
rect 417808 182866 418128 182898
rect 448528 183454 448848 183486
rect 448528 183218 448570 183454
rect 448806 183218 448848 183454
rect 448528 183134 448848 183218
rect 448528 182898 448570 183134
rect 448806 182898 448848 183134
rect 448528 182866 448848 182898
rect 479248 183454 479568 183486
rect 479248 183218 479290 183454
rect 479526 183218 479568 183454
rect 479248 183134 479568 183218
rect 479248 182898 479290 183134
rect 479526 182898 479568 183134
rect 479248 182866 479568 182898
rect 509968 183454 510288 183486
rect 509968 183218 510010 183454
rect 510246 183218 510288 183454
rect 509968 183134 510288 183218
rect 509968 182898 510010 183134
rect 510246 182898 510288 183134
rect 509968 182866 510288 182898
rect 540688 183454 541008 183486
rect 540688 183218 540730 183454
rect 540966 183218 541008 183454
rect 540688 183134 541008 183218
rect 540688 182898 540730 183134
rect 540966 182898 541008 183134
rect 540688 182866 541008 182898
rect 552954 158614 553574 194058
rect 552954 158378 552986 158614
rect 553222 158378 553306 158614
rect 553542 158378 553574 158614
rect 552954 158294 553574 158378
rect 552954 158058 552986 158294
rect 553222 158058 553306 158294
rect 553542 158058 553574 158294
rect 257514 150938 257546 151174
rect 257782 150938 257866 151174
rect 258102 150938 258134 151174
rect 257514 150854 258134 150938
rect 257514 150618 257546 150854
rect 257782 150618 257866 150854
rect 258102 150618 258134 150854
rect 257514 115174 258134 150618
rect 279568 151174 279888 151206
rect 279568 150938 279610 151174
rect 279846 150938 279888 151174
rect 279568 150854 279888 150938
rect 279568 150618 279610 150854
rect 279846 150618 279888 150854
rect 279568 150586 279888 150618
rect 310288 151174 310608 151206
rect 310288 150938 310330 151174
rect 310566 150938 310608 151174
rect 310288 150854 310608 150938
rect 310288 150618 310330 150854
rect 310566 150618 310608 150854
rect 310288 150586 310608 150618
rect 341008 151174 341328 151206
rect 341008 150938 341050 151174
rect 341286 150938 341328 151174
rect 341008 150854 341328 150938
rect 341008 150618 341050 150854
rect 341286 150618 341328 150854
rect 341008 150586 341328 150618
rect 371728 151174 372048 151206
rect 371728 150938 371770 151174
rect 372006 150938 372048 151174
rect 371728 150854 372048 150938
rect 371728 150618 371770 150854
rect 372006 150618 372048 150854
rect 371728 150586 372048 150618
rect 402448 151174 402768 151206
rect 402448 150938 402490 151174
rect 402726 150938 402768 151174
rect 402448 150854 402768 150938
rect 402448 150618 402490 150854
rect 402726 150618 402768 150854
rect 402448 150586 402768 150618
rect 433168 151174 433488 151206
rect 433168 150938 433210 151174
rect 433446 150938 433488 151174
rect 433168 150854 433488 150938
rect 433168 150618 433210 150854
rect 433446 150618 433488 150854
rect 433168 150586 433488 150618
rect 463888 151174 464208 151206
rect 463888 150938 463930 151174
rect 464166 150938 464208 151174
rect 463888 150854 464208 150938
rect 463888 150618 463930 150854
rect 464166 150618 464208 150854
rect 463888 150586 464208 150618
rect 494608 151174 494928 151206
rect 494608 150938 494650 151174
rect 494886 150938 494928 151174
rect 494608 150854 494928 150938
rect 494608 150618 494650 150854
rect 494886 150618 494928 150854
rect 494608 150586 494928 150618
rect 525328 151174 525648 151206
rect 525328 150938 525370 151174
rect 525606 150938 525648 151174
rect 525328 150854 525648 150938
rect 525328 150618 525370 150854
rect 525606 150618 525648 150854
rect 525328 150586 525648 150618
rect 264208 147454 264528 147486
rect 264208 147218 264250 147454
rect 264486 147218 264528 147454
rect 264208 147134 264528 147218
rect 264208 146898 264250 147134
rect 264486 146898 264528 147134
rect 264208 146866 264528 146898
rect 294928 147454 295248 147486
rect 294928 147218 294970 147454
rect 295206 147218 295248 147454
rect 294928 147134 295248 147218
rect 294928 146898 294970 147134
rect 295206 146898 295248 147134
rect 294928 146866 295248 146898
rect 325648 147454 325968 147486
rect 325648 147218 325690 147454
rect 325926 147218 325968 147454
rect 325648 147134 325968 147218
rect 325648 146898 325690 147134
rect 325926 146898 325968 147134
rect 325648 146866 325968 146898
rect 356368 147454 356688 147486
rect 356368 147218 356410 147454
rect 356646 147218 356688 147454
rect 356368 147134 356688 147218
rect 356368 146898 356410 147134
rect 356646 146898 356688 147134
rect 356368 146866 356688 146898
rect 387088 147454 387408 147486
rect 387088 147218 387130 147454
rect 387366 147218 387408 147454
rect 387088 147134 387408 147218
rect 387088 146898 387130 147134
rect 387366 146898 387408 147134
rect 387088 146866 387408 146898
rect 417808 147454 418128 147486
rect 417808 147218 417850 147454
rect 418086 147218 418128 147454
rect 417808 147134 418128 147218
rect 417808 146898 417850 147134
rect 418086 146898 418128 147134
rect 417808 146866 418128 146898
rect 448528 147454 448848 147486
rect 448528 147218 448570 147454
rect 448806 147218 448848 147454
rect 448528 147134 448848 147218
rect 448528 146898 448570 147134
rect 448806 146898 448848 147134
rect 448528 146866 448848 146898
rect 479248 147454 479568 147486
rect 479248 147218 479290 147454
rect 479526 147218 479568 147454
rect 479248 147134 479568 147218
rect 479248 146898 479290 147134
rect 479526 146898 479568 147134
rect 479248 146866 479568 146898
rect 509968 147454 510288 147486
rect 509968 147218 510010 147454
rect 510246 147218 510288 147454
rect 509968 147134 510288 147218
rect 509968 146898 510010 147134
rect 510246 146898 510288 147134
rect 509968 146866 510288 146898
rect 540688 147454 541008 147486
rect 540688 147218 540730 147454
rect 540966 147218 541008 147454
rect 540688 147134 541008 147218
rect 540688 146898 540730 147134
rect 540966 146898 541008 147134
rect 540688 146866 541008 146898
rect 552954 122614 553574 158058
rect 552954 122378 552986 122614
rect 553222 122378 553306 122614
rect 553542 122378 553574 122614
rect 552954 122294 553574 122378
rect 552954 122058 552986 122294
rect 553222 122058 553306 122294
rect 553542 122058 553574 122294
rect 257514 114938 257546 115174
rect 257782 114938 257866 115174
rect 258102 114938 258134 115174
rect 257514 114854 258134 114938
rect 257514 114618 257546 114854
rect 257782 114618 257866 114854
rect 258102 114618 258134 114854
rect 257514 79174 258134 114618
rect 279568 115174 279888 115206
rect 279568 114938 279610 115174
rect 279846 114938 279888 115174
rect 279568 114854 279888 114938
rect 279568 114618 279610 114854
rect 279846 114618 279888 114854
rect 279568 114586 279888 114618
rect 310288 115174 310608 115206
rect 310288 114938 310330 115174
rect 310566 114938 310608 115174
rect 310288 114854 310608 114938
rect 310288 114618 310330 114854
rect 310566 114618 310608 114854
rect 310288 114586 310608 114618
rect 341008 115174 341328 115206
rect 341008 114938 341050 115174
rect 341286 114938 341328 115174
rect 341008 114854 341328 114938
rect 341008 114618 341050 114854
rect 341286 114618 341328 114854
rect 341008 114586 341328 114618
rect 371728 115174 372048 115206
rect 371728 114938 371770 115174
rect 372006 114938 372048 115174
rect 371728 114854 372048 114938
rect 371728 114618 371770 114854
rect 372006 114618 372048 114854
rect 371728 114586 372048 114618
rect 402448 115174 402768 115206
rect 402448 114938 402490 115174
rect 402726 114938 402768 115174
rect 402448 114854 402768 114938
rect 402448 114618 402490 114854
rect 402726 114618 402768 114854
rect 402448 114586 402768 114618
rect 433168 115174 433488 115206
rect 433168 114938 433210 115174
rect 433446 114938 433488 115174
rect 433168 114854 433488 114938
rect 433168 114618 433210 114854
rect 433446 114618 433488 114854
rect 433168 114586 433488 114618
rect 463888 115174 464208 115206
rect 463888 114938 463930 115174
rect 464166 114938 464208 115174
rect 463888 114854 464208 114938
rect 463888 114618 463930 114854
rect 464166 114618 464208 114854
rect 463888 114586 464208 114618
rect 494608 115174 494928 115206
rect 494608 114938 494650 115174
rect 494886 114938 494928 115174
rect 494608 114854 494928 114938
rect 494608 114618 494650 114854
rect 494886 114618 494928 114854
rect 494608 114586 494928 114618
rect 525328 115174 525648 115206
rect 525328 114938 525370 115174
rect 525606 114938 525648 115174
rect 525328 114854 525648 114938
rect 525328 114618 525370 114854
rect 525606 114618 525648 114854
rect 525328 114586 525648 114618
rect 264208 111454 264528 111486
rect 264208 111218 264250 111454
rect 264486 111218 264528 111454
rect 264208 111134 264528 111218
rect 264208 110898 264250 111134
rect 264486 110898 264528 111134
rect 264208 110866 264528 110898
rect 294928 111454 295248 111486
rect 294928 111218 294970 111454
rect 295206 111218 295248 111454
rect 294928 111134 295248 111218
rect 294928 110898 294970 111134
rect 295206 110898 295248 111134
rect 294928 110866 295248 110898
rect 325648 111454 325968 111486
rect 325648 111218 325690 111454
rect 325926 111218 325968 111454
rect 325648 111134 325968 111218
rect 325648 110898 325690 111134
rect 325926 110898 325968 111134
rect 325648 110866 325968 110898
rect 356368 111454 356688 111486
rect 356368 111218 356410 111454
rect 356646 111218 356688 111454
rect 356368 111134 356688 111218
rect 356368 110898 356410 111134
rect 356646 110898 356688 111134
rect 356368 110866 356688 110898
rect 387088 111454 387408 111486
rect 387088 111218 387130 111454
rect 387366 111218 387408 111454
rect 387088 111134 387408 111218
rect 387088 110898 387130 111134
rect 387366 110898 387408 111134
rect 387088 110866 387408 110898
rect 417808 111454 418128 111486
rect 417808 111218 417850 111454
rect 418086 111218 418128 111454
rect 417808 111134 418128 111218
rect 417808 110898 417850 111134
rect 418086 110898 418128 111134
rect 417808 110866 418128 110898
rect 448528 111454 448848 111486
rect 448528 111218 448570 111454
rect 448806 111218 448848 111454
rect 448528 111134 448848 111218
rect 448528 110898 448570 111134
rect 448806 110898 448848 111134
rect 448528 110866 448848 110898
rect 479248 111454 479568 111486
rect 479248 111218 479290 111454
rect 479526 111218 479568 111454
rect 479248 111134 479568 111218
rect 479248 110898 479290 111134
rect 479526 110898 479568 111134
rect 479248 110866 479568 110898
rect 509968 111454 510288 111486
rect 509968 111218 510010 111454
rect 510246 111218 510288 111454
rect 509968 111134 510288 111218
rect 509968 110898 510010 111134
rect 510246 110898 510288 111134
rect 509968 110866 510288 110898
rect 540688 111454 541008 111486
rect 540688 111218 540730 111454
rect 540966 111218 541008 111454
rect 540688 111134 541008 111218
rect 540688 110898 540730 111134
rect 540966 110898 541008 111134
rect 540688 110866 541008 110898
rect 552954 86614 553574 122058
rect 552954 86378 552986 86614
rect 553222 86378 553306 86614
rect 553542 86378 553574 86614
rect 552954 86294 553574 86378
rect 552954 86058 552986 86294
rect 553222 86058 553306 86294
rect 553542 86058 553574 86294
rect 257514 78938 257546 79174
rect 257782 78938 257866 79174
rect 258102 78938 258134 79174
rect 257514 78854 258134 78938
rect 257514 78618 257546 78854
rect 257782 78618 257866 78854
rect 258102 78618 258134 78854
rect 257514 43174 258134 78618
rect 279568 79174 279888 79206
rect 279568 78938 279610 79174
rect 279846 78938 279888 79174
rect 279568 78854 279888 78938
rect 279568 78618 279610 78854
rect 279846 78618 279888 78854
rect 279568 78586 279888 78618
rect 310288 79174 310608 79206
rect 310288 78938 310330 79174
rect 310566 78938 310608 79174
rect 310288 78854 310608 78938
rect 310288 78618 310330 78854
rect 310566 78618 310608 78854
rect 310288 78586 310608 78618
rect 341008 79174 341328 79206
rect 341008 78938 341050 79174
rect 341286 78938 341328 79174
rect 341008 78854 341328 78938
rect 341008 78618 341050 78854
rect 341286 78618 341328 78854
rect 341008 78586 341328 78618
rect 371728 79174 372048 79206
rect 371728 78938 371770 79174
rect 372006 78938 372048 79174
rect 371728 78854 372048 78938
rect 371728 78618 371770 78854
rect 372006 78618 372048 78854
rect 371728 78586 372048 78618
rect 402448 79174 402768 79206
rect 402448 78938 402490 79174
rect 402726 78938 402768 79174
rect 402448 78854 402768 78938
rect 402448 78618 402490 78854
rect 402726 78618 402768 78854
rect 402448 78586 402768 78618
rect 433168 79174 433488 79206
rect 433168 78938 433210 79174
rect 433446 78938 433488 79174
rect 433168 78854 433488 78938
rect 433168 78618 433210 78854
rect 433446 78618 433488 78854
rect 433168 78586 433488 78618
rect 463888 79174 464208 79206
rect 463888 78938 463930 79174
rect 464166 78938 464208 79174
rect 463888 78854 464208 78938
rect 463888 78618 463930 78854
rect 464166 78618 464208 78854
rect 463888 78586 464208 78618
rect 494608 79174 494928 79206
rect 494608 78938 494650 79174
rect 494886 78938 494928 79174
rect 494608 78854 494928 78938
rect 494608 78618 494650 78854
rect 494886 78618 494928 78854
rect 494608 78586 494928 78618
rect 525328 79174 525648 79206
rect 525328 78938 525370 79174
rect 525606 78938 525648 79174
rect 525328 78854 525648 78938
rect 525328 78618 525370 78854
rect 525606 78618 525648 78854
rect 525328 78586 525648 78618
rect 264208 75454 264528 75486
rect 264208 75218 264250 75454
rect 264486 75218 264528 75454
rect 264208 75134 264528 75218
rect 264208 74898 264250 75134
rect 264486 74898 264528 75134
rect 264208 74866 264528 74898
rect 294928 75454 295248 75486
rect 294928 75218 294970 75454
rect 295206 75218 295248 75454
rect 294928 75134 295248 75218
rect 294928 74898 294970 75134
rect 295206 74898 295248 75134
rect 294928 74866 295248 74898
rect 325648 75454 325968 75486
rect 325648 75218 325690 75454
rect 325926 75218 325968 75454
rect 325648 75134 325968 75218
rect 325648 74898 325690 75134
rect 325926 74898 325968 75134
rect 325648 74866 325968 74898
rect 356368 75454 356688 75486
rect 356368 75218 356410 75454
rect 356646 75218 356688 75454
rect 356368 75134 356688 75218
rect 356368 74898 356410 75134
rect 356646 74898 356688 75134
rect 356368 74866 356688 74898
rect 387088 75454 387408 75486
rect 387088 75218 387130 75454
rect 387366 75218 387408 75454
rect 387088 75134 387408 75218
rect 387088 74898 387130 75134
rect 387366 74898 387408 75134
rect 387088 74866 387408 74898
rect 417808 75454 418128 75486
rect 417808 75218 417850 75454
rect 418086 75218 418128 75454
rect 417808 75134 418128 75218
rect 417808 74898 417850 75134
rect 418086 74898 418128 75134
rect 417808 74866 418128 74898
rect 448528 75454 448848 75486
rect 448528 75218 448570 75454
rect 448806 75218 448848 75454
rect 448528 75134 448848 75218
rect 448528 74898 448570 75134
rect 448806 74898 448848 75134
rect 448528 74866 448848 74898
rect 479248 75454 479568 75486
rect 479248 75218 479290 75454
rect 479526 75218 479568 75454
rect 479248 75134 479568 75218
rect 479248 74898 479290 75134
rect 479526 74898 479568 75134
rect 479248 74866 479568 74898
rect 509968 75454 510288 75486
rect 509968 75218 510010 75454
rect 510246 75218 510288 75454
rect 509968 75134 510288 75218
rect 509968 74898 510010 75134
rect 510246 74898 510288 75134
rect 509968 74866 510288 74898
rect 540688 75454 541008 75486
rect 540688 75218 540730 75454
rect 540966 75218 541008 75454
rect 540688 75134 541008 75218
rect 540688 74898 540730 75134
rect 540966 74898 541008 75134
rect 540688 74866 541008 74898
rect 552954 50614 553574 86058
rect 552954 50378 552986 50614
rect 553222 50378 553306 50614
rect 553542 50378 553574 50614
rect 552954 50294 553574 50378
rect 258579 50148 258645 50149
rect 258579 50084 258580 50148
rect 258644 50084 258645 50148
rect 258579 50083 258645 50084
rect 257514 42938 257546 43174
rect 257782 42938 257866 43174
rect 258102 42938 258134 43174
rect 257514 42854 258134 42938
rect 257514 42618 257546 42854
rect 257782 42618 257866 42854
rect 258102 42618 258134 42854
rect 257514 7174 258134 42618
rect 257514 6938 257546 7174
rect 257782 6938 257866 7174
rect 258102 6938 258134 7174
rect 257514 6854 258134 6938
rect 257514 6618 257546 6854
rect 257782 6618 257866 6854
rect 258102 6618 258134 6854
rect 257514 -1306 258134 6618
rect 258582 3501 258642 50083
rect 552954 50058 552986 50294
rect 553222 50058 553306 50294
rect 553542 50058 553574 50294
rect 279568 43174 279888 43206
rect 261234 10894 261854 43007
rect 261234 10658 261266 10894
rect 261502 10658 261586 10894
rect 261822 10658 261854 10894
rect 261234 10574 261854 10658
rect 261234 10338 261266 10574
rect 261502 10338 261586 10574
rect 261822 10338 261854 10574
rect 258579 3500 258645 3501
rect 258579 3436 258580 3500
rect 258644 3436 258645 3500
rect 258579 3435 258645 3436
rect 257514 -1542 257546 -1306
rect 257782 -1542 257866 -1306
rect 258102 -1542 258134 -1306
rect 257514 -1626 258134 -1542
rect 257514 -1862 257546 -1626
rect 257782 -1862 257866 -1626
rect 258102 -1862 258134 -1626
rect 257514 -7654 258134 -1862
rect 261234 -2266 261854 10338
rect 261234 -2502 261266 -2266
rect 261502 -2502 261586 -2266
rect 261822 -2502 261854 -2266
rect 261234 -2586 261854 -2502
rect 261234 -2822 261266 -2586
rect 261502 -2822 261586 -2586
rect 261822 -2822 261854 -2586
rect 261234 -7654 261854 -2822
rect 264954 14614 265574 43007
rect 264954 14378 264986 14614
rect 265222 14378 265306 14614
rect 265542 14378 265574 14614
rect 264954 14294 265574 14378
rect 264954 14058 264986 14294
rect 265222 14058 265306 14294
rect 265542 14058 265574 14294
rect 264954 -3226 265574 14058
rect 264954 -3462 264986 -3226
rect 265222 -3462 265306 -3226
rect 265542 -3462 265574 -3226
rect 264954 -3546 265574 -3462
rect 264954 -3782 264986 -3546
rect 265222 -3782 265306 -3546
rect 265542 -3782 265574 -3546
rect 264954 -7654 265574 -3782
rect 268674 18334 269294 43007
rect 268674 18098 268706 18334
rect 268942 18098 269026 18334
rect 269262 18098 269294 18334
rect 268674 18014 269294 18098
rect 268674 17778 268706 18014
rect 268942 17778 269026 18014
rect 269262 17778 269294 18014
rect 268674 -4186 269294 17778
rect 268674 -4422 268706 -4186
rect 268942 -4422 269026 -4186
rect 269262 -4422 269294 -4186
rect 268674 -4506 269294 -4422
rect 268674 -4742 268706 -4506
rect 268942 -4742 269026 -4506
rect 269262 -4742 269294 -4506
rect 268674 -7654 269294 -4742
rect 272394 22054 273014 43007
rect 272394 21818 272426 22054
rect 272662 21818 272746 22054
rect 272982 21818 273014 22054
rect 272394 21734 273014 21818
rect 272394 21498 272426 21734
rect 272662 21498 272746 21734
rect 272982 21498 273014 21734
rect 272394 -5146 273014 21498
rect 272394 -5382 272426 -5146
rect 272662 -5382 272746 -5146
rect 272982 -5382 273014 -5146
rect 272394 -5466 273014 -5382
rect 272394 -5702 272426 -5466
rect 272662 -5702 272746 -5466
rect 272982 -5702 273014 -5466
rect 272394 -7654 273014 -5702
rect 276114 25774 276734 43007
rect 279568 42938 279610 43174
rect 279846 42938 279888 43174
rect 310288 43174 310608 43206
rect 279568 42854 279888 42938
rect 279568 42618 279610 42854
rect 279846 42618 279888 42854
rect 279568 42586 279888 42618
rect 276114 25538 276146 25774
rect 276382 25538 276466 25774
rect 276702 25538 276734 25774
rect 276114 25454 276734 25538
rect 276114 25218 276146 25454
rect 276382 25218 276466 25454
rect 276702 25218 276734 25454
rect 276114 -6106 276734 25218
rect 276114 -6342 276146 -6106
rect 276382 -6342 276466 -6106
rect 276702 -6342 276734 -6106
rect 276114 -6426 276734 -6342
rect 276114 -6662 276146 -6426
rect 276382 -6662 276466 -6426
rect 276702 -6662 276734 -6426
rect 276114 -7654 276734 -6662
rect 279834 29494 280454 40068
rect 279834 29258 279866 29494
rect 280102 29258 280186 29494
rect 280422 29258 280454 29494
rect 279834 29174 280454 29258
rect 279834 28938 279866 29174
rect 280102 28938 280186 29174
rect 280422 28938 280454 29174
rect 279834 -7066 280454 28938
rect 279834 -7302 279866 -7066
rect 280102 -7302 280186 -7066
rect 280422 -7302 280454 -7066
rect 279834 -7386 280454 -7302
rect 279834 -7622 279866 -7386
rect 280102 -7622 280186 -7386
rect 280422 -7622 280454 -7386
rect 279834 -7654 280454 -7622
rect 289794 39454 290414 43007
rect 289794 39218 289826 39454
rect 290062 39218 290146 39454
rect 290382 39218 290414 39454
rect 289794 39134 290414 39218
rect 289794 38898 289826 39134
rect 290062 38898 290146 39134
rect 290382 38898 290414 39134
rect 289794 3454 290414 38898
rect 289794 3218 289826 3454
rect 290062 3218 290146 3454
rect 290382 3218 290414 3454
rect 289794 3134 290414 3218
rect 289794 2898 289826 3134
rect 290062 2898 290146 3134
rect 290382 2898 290414 3134
rect 289794 -346 290414 2898
rect 289794 -582 289826 -346
rect 290062 -582 290146 -346
rect 290382 -582 290414 -346
rect 289794 -666 290414 -582
rect 289794 -902 289826 -666
rect 290062 -902 290146 -666
rect 290382 -902 290414 -666
rect 289794 -7654 290414 -902
rect 293514 7174 294134 43007
rect 293514 6938 293546 7174
rect 293782 6938 293866 7174
rect 294102 6938 294134 7174
rect 293514 6854 294134 6938
rect 293514 6618 293546 6854
rect 293782 6618 293866 6854
rect 294102 6618 294134 6854
rect 293514 -1306 294134 6618
rect 293514 -1542 293546 -1306
rect 293782 -1542 293866 -1306
rect 294102 -1542 294134 -1306
rect 293514 -1626 294134 -1542
rect 293514 -1862 293546 -1626
rect 293782 -1862 293866 -1626
rect 294102 -1862 294134 -1626
rect 293514 -7654 294134 -1862
rect 297234 10894 297854 43007
rect 297234 10658 297266 10894
rect 297502 10658 297586 10894
rect 297822 10658 297854 10894
rect 297234 10574 297854 10658
rect 297234 10338 297266 10574
rect 297502 10338 297586 10574
rect 297822 10338 297854 10574
rect 297234 -2266 297854 10338
rect 297234 -2502 297266 -2266
rect 297502 -2502 297586 -2266
rect 297822 -2502 297854 -2266
rect 297234 -2586 297854 -2502
rect 297234 -2822 297266 -2586
rect 297502 -2822 297586 -2586
rect 297822 -2822 297854 -2586
rect 297234 -7654 297854 -2822
rect 300954 14614 301574 43007
rect 300954 14378 300986 14614
rect 301222 14378 301306 14614
rect 301542 14378 301574 14614
rect 300954 14294 301574 14378
rect 300954 14058 300986 14294
rect 301222 14058 301306 14294
rect 301542 14058 301574 14294
rect 300954 -3226 301574 14058
rect 300954 -3462 300986 -3226
rect 301222 -3462 301306 -3226
rect 301542 -3462 301574 -3226
rect 300954 -3546 301574 -3462
rect 300954 -3782 300986 -3546
rect 301222 -3782 301306 -3546
rect 301542 -3782 301574 -3546
rect 300954 -7654 301574 -3782
rect 304674 18334 305294 43007
rect 304674 18098 304706 18334
rect 304942 18098 305026 18334
rect 305262 18098 305294 18334
rect 304674 18014 305294 18098
rect 304674 17778 304706 18014
rect 304942 17778 305026 18014
rect 305262 17778 305294 18014
rect 304674 -4186 305294 17778
rect 304674 -4422 304706 -4186
rect 304942 -4422 305026 -4186
rect 305262 -4422 305294 -4186
rect 304674 -4506 305294 -4422
rect 304674 -4742 304706 -4506
rect 304942 -4742 305026 -4506
rect 305262 -4742 305294 -4506
rect 304674 -7654 305294 -4742
rect 308394 22054 309014 43007
rect 310288 42938 310330 43174
rect 310566 42938 310608 43174
rect 341008 43174 341328 43206
rect 310288 42854 310608 42938
rect 310288 42618 310330 42854
rect 310566 42618 310608 42854
rect 310288 42586 310608 42618
rect 308394 21818 308426 22054
rect 308662 21818 308746 22054
rect 308982 21818 309014 22054
rect 308394 21734 309014 21818
rect 308394 21498 308426 21734
rect 308662 21498 308746 21734
rect 308982 21498 309014 21734
rect 308394 -5146 309014 21498
rect 308394 -5382 308426 -5146
rect 308662 -5382 308746 -5146
rect 308982 -5382 309014 -5146
rect 308394 -5466 309014 -5382
rect 308394 -5702 308426 -5466
rect 308662 -5702 308746 -5466
rect 308982 -5702 309014 -5466
rect 308394 -7654 309014 -5702
rect 312114 25774 312734 43007
rect 312114 25538 312146 25774
rect 312382 25538 312466 25774
rect 312702 25538 312734 25774
rect 312114 25454 312734 25538
rect 312114 25218 312146 25454
rect 312382 25218 312466 25454
rect 312702 25218 312734 25454
rect 312114 -6106 312734 25218
rect 312114 -6342 312146 -6106
rect 312382 -6342 312466 -6106
rect 312702 -6342 312734 -6106
rect 312114 -6426 312734 -6342
rect 312114 -6662 312146 -6426
rect 312382 -6662 312466 -6426
rect 312702 -6662 312734 -6426
rect 312114 -7654 312734 -6662
rect 315834 29494 316454 43007
rect 315834 29258 315866 29494
rect 316102 29258 316186 29494
rect 316422 29258 316454 29494
rect 315834 29174 316454 29258
rect 315834 28938 315866 29174
rect 316102 28938 316186 29174
rect 316422 28938 316454 29174
rect 315834 -7066 316454 28938
rect 315834 -7302 315866 -7066
rect 316102 -7302 316186 -7066
rect 316422 -7302 316454 -7066
rect 315834 -7386 316454 -7302
rect 315834 -7622 315866 -7386
rect 316102 -7622 316186 -7386
rect 316422 -7622 316454 -7386
rect 315834 -7654 316454 -7622
rect 325794 39454 326414 40068
rect 325794 39218 325826 39454
rect 326062 39218 326146 39454
rect 326382 39218 326414 39454
rect 325794 39134 326414 39218
rect 325794 38898 325826 39134
rect 326062 38898 326146 39134
rect 326382 38898 326414 39134
rect 325794 3454 326414 38898
rect 325794 3218 325826 3454
rect 326062 3218 326146 3454
rect 326382 3218 326414 3454
rect 325794 3134 326414 3218
rect 325794 2898 325826 3134
rect 326062 2898 326146 3134
rect 326382 2898 326414 3134
rect 325794 -346 326414 2898
rect 325794 -582 325826 -346
rect 326062 -582 326146 -346
rect 326382 -582 326414 -346
rect 325794 -666 326414 -582
rect 325794 -902 325826 -666
rect 326062 -902 326146 -666
rect 326382 -902 326414 -666
rect 325794 -7654 326414 -902
rect 329514 7174 330134 43007
rect 329514 6938 329546 7174
rect 329782 6938 329866 7174
rect 330102 6938 330134 7174
rect 329514 6854 330134 6938
rect 329514 6618 329546 6854
rect 329782 6618 329866 6854
rect 330102 6618 330134 6854
rect 329514 -1306 330134 6618
rect 329514 -1542 329546 -1306
rect 329782 -1542 329866 -1306
rect 330102 -1542 330134 -1306
rect 329514 -1626 330134 -1542
rect 329514 -1862 329546 -1626
rect 329782 -1862 329866 -1626
rect 330102 -1862 330134 -1626
rect 329514 -7654 330134 -1862
rect 333234 10894 333854 43007
rect 333234 10658 333266 10894
rect 333502 10658 333586 10894
rect 333822 10658 333854 10894
rect 333234 10574 333854 10658
rect 333234 10338 333266 10574
rect 333502 10338 333586 10574
rect 333822 10338 333854 10574
rect 333234 -2266 333854 10338
rect 333234 -2502 333266 -2266
rect 333502 -2502 333586 -2266
rect 333822 -2502 333854 -2266
rect 333234 -2586 333854 -2502
rect 333234 -2822 333266 -2586
rect 333502 -2822 333586 -2586
rect 333822 -2822 333854 -2586
rect 333234 -7654 333854 -2822
rect 336954 14614 337574 43007
rect 341008 42938 341050 43174
rect 341286 42938 341328 43174
rect 371728 43174 372048 43206
rect 341008 42854 341328 42938
rect 341008 42618 341050 42854
rect 341286 42618 341328 42854
rect 341008 42586 341328 42618
rect 336954 14378 336986 14614
rect 337222 14378 337306 14614
rect 337542 14378 337574 14614
rect 336954 14294 337574 14378
rect 336954 14058 336986 14294
rect 337222 14058 337306 14294
rect 337542 14058 337574 14294
rect 336954 -3226 337574 14058
rect 336954 -3462 336986 -3226
rect 337222 -3462 337306 -3226
rect 337542 -3462 337574 -3226
rect 336954 -3546 337574 -3462
rect 336954 -3782 336986 -3546
rect 337222 -3782 337306 -3546
rect 337542 -3782 337574 -3546
rect 336954 -7654 337574 -3782
rect 340674 18334 341294 40068
rect 340674 18098 340706 18334
rect 340942 18098 341026 18334
rect 341262 18098 341294 18334
rect 340674 18014 341294 18098
rect 340674 17778 340706 18014
rect 340942 17778 341026 18014
rect 341262 17778 341294 18014
rect 340674 -4186 341294 17778
rect 340674 -4422 340706 -4186
rect 340942 -4422 341026 -4186
rect 341262 -4422 341294 -4186
rect 340674 -4506 341294 -4422
rect 340674 -4742 340706 -4506
rect 340942 -4742 341026 -4506
rect 341262 -4742 341294 -4506
rect 340674 -7654 341294 -4742
rect 344394 22054 345014 43007
rect 344394 21818 344426 22054
rect 344662 21818 344746 22054
rect 344982 21818 345014 22054
rect 344394 21734 345014 21818
rect 344394 21498 344426 21734
rect 344662 21498 344746 21734
rect 344982 21498 345014 21734
rect 344394 -5146 345014 21498
rect 344394 -5382 344426 -5146
rect 344662 -5382 344746 -5146
rect 344982 -5382 345014 -5146
rect 344394 -5466 345014 -5382
rect 344394 -5702 344426 -5466
rect 344662 -5702 344746 -5466
rect 344982 -5702 345014 -5466
rect 344394 -7654 345014 -5702
rect 348114 25774 348734 43007
rect 348114 25538 348146 25774
rect 348382 25538 348466 25774
rect 348702 25538 348734 25774
rect 348114 25454 348734 25538
rect 348114 25218 348146 25454
rect 348382 25218 348466 25454
rect 348702 25218 348734 25454
rect 348114 -6106 348734 25218
rect 348114 -6342 348146 -6106
rect 348382 -6342 348466 -6106
rect 348702 -6342 348734 -6106
rect 348114 -6426 348734 -6342
rect 348114 -6662 348146 -6426
rect 348382 -6662 348466 -6426
rect 348702 -6662 348734 -6426
rect 348114 -7654 348734 -6662
rect 351834 29494 352454 43007
rect 351834 29258 351866 29494
rect 352102 29258 352186 29494
rect 352422 29258 352454 29494
rect 351834 29174 352454 29258
rect 351834 28938 351866 29174
rect 352102 28938 352186 29174
rect 352422 28938 352454 29174
rect 351834 -7066 352454 28938
rect 351834 -7302 351866 -7066
rect 352102 -7302 352186 -7066
rect 352422 -7302 352454 -7066
rect 351834 -7386 352454 -7302
rect 351834 -7622 351866 -7386
rect 352102 -7622 352186 -7386
rect 352422 -7622 352454 -7386
rect 351834 -7654 352454 -7622
rect 361794 39454 362414 43007
rect 361794 39218 361826 39454
rect 362062 39218 362146 39454
rect 362382 39218 362414 39454
rect 361794 39134 362414 39218
rect 361794 38898 361826 39134
rect 362062 38898 362146 39134
rect 362382 38898 362414 39134
rect 361794 3454 362414 38898
rect 361794 3218 361826 3454
rect 362062 3218 362146 3454
rect 362382 3218 362414 3454
rect 361794 3134 362414 3218
rect 361794 2898 361826 3134
rect 362062 2898 362146 3134
rect 362382 2898 362414 3134
rect 361794 -346 362414 2898
rect 361794 -582 361826 -346
rect 362062 -582 362146 -346
rect 362382 -582 362414 -346
rect 361794 -666 362414 -582
rect 361794 -902 361826 -666
rect 362062 -902 362146 -666
rect 362382 -902 362414 -666
rect 361794 -7654 362414 -902
rect 365514 7174 366134 43007
rect 365514 6938 365546 7174
rect 365782 6938 365866 7174
rect 366102 6938 366134 7174
rect 365514 6854 366134 6938
rect 365514 6618 365546 6854
rect 365782 6618 365866 6854
rect 366102 6618 366134 6854
rect 365514 -1306 366134 6618
rect 365514 -1542 365546 -1306
rect 365782 -1542 365866 -1306
rect 366102 -1542 366134 -1306
rect 365514 -1626 366134 -1542
rect 365514 -1862 365546 -1626
rect 365782 -1862 365866 -1626
rect 366102 -1862 366134 -1626
rect 365514 -7654 366134 -1862
rect 369234 10894 369854 43007
rect 371728 42938 371770 43174
rect 372006 42938 372048 43174
rect 402448 43174 402768 43206
rect 371728 42854 372048 42938
rect 371728 42618 371770 42854
rect 372006 42618 372048 42854
rect 371728 42586 372048 42618
rect 369234 10658 369266 10894
rect 369502 10658 369586 10894
rect 369822 10658 369854 10894
rect 369234 10574 369854 10658
rect 369234 10338 369266 10574
rect 369502 10338 369586 10574
rect 369822 10338 369854 10574
rect 369234 -2266 369854 10338
rect 369234 -2502 369266 -2266
rect 369502 -2502 369586 -2266
rect 369822 -2502 369854 -2266
rect 369234 -2586 369854 -2502
rect 369234 -2822 369266 -2586
rect 369502 -2822 369586 -2586
rect 369822 -2822 369854 -2586
rect 369234 -7654 369854 -2822
rect 372954 14614 373574 43007
rect 372954 14378 372986 14614
rect 373222 14378 373306 14614
rect 373542 14378 373574 14614
rect 372954 14294 373574 14378
rect 372954 14058 372986 14294
rect 373222 14058 373306 14294
rect 373542 14058 373574 14294
rect 372954 -3226 373574 14058
rect 372954 -3462 372986 -3226
rect 373222 -3462 373306 -3226
rect 373542 -3462 373574 -3226
rect 372954 -3546 373574 -3462
rect 372954 -3782 372986 -3546
rect 373222 -3782 373306 -3546
rect 373542 -3782 373574 -3546
rect 372954 -7654 373574 -3782
rect 376674 18334 377294 43007
rect 376674 18098 376706 18334
rect 376942 18098 377026 18334
rect 377262 18098 377294 18334
rect 376674 18014 377294 18098
rect 376674 17778 376706 18014
rect 376942 17778 377026 18014
rect 377262 17778 377294 18014
rect 376674 -4186 377294 17778
rect 376674 -4422 376706 -4186
rect 376942 -4422 377026 -4186
rect 377262 -4422 377294 -4186
rect 376674 -4506 377294 -4422
rect 376674 -4742 376706 -4506
rect 376942 -4742 377026 -4506
rect 377262 -4742 377294 -4506
rect 376674 -7654 377294 -4742
rect 380394 22054 381014 43007
rect 380394 21818 380426 22054
rect 380662 21818 380746 22054
rect 380982 21818 381014 22054
rect 380394 21734 381014 21818
rect 380394 21498 380426 21734
rect 380662 21498 380746 21734
rect 380982 21498 381014 21734
rect 380394 -5146 381014 21498
rect 380394 -5382 380426 -5146
rect 380662 -5382 380746 -5146
rect 380982 -5382 381014 -5146
rect 380394 -5466 381014 -5382
rect 380394 -5702 380426 -5466
rect 380662 -5702 380746 -5466
rect 380982 -5702 381014 -5466
rect 380394 -7654 381014 -5702
rect 384114 25774 384734 43007
rect 384114 25538 384146 25774
rect 384382 25538 384466 25774
rect 384702 25538 384734 25774
rect 384114 25454 384734 25538
rect 384114 25218 384146 25454
rect 384382 25218 384466 25454
rect 384702 25218 384734 25454
rect 384114 -6106 384734 25218
rect 384114 -6342 384146 -6106
rect 384382 -6342 384466 -6106
rect 384702 -6342 384734 -6106
rect 384114 -6426 384734 -6342
rect 384114 -6662 384146 -6426
rect 384382 -6662 384466 -6426
rect 384702 -6662 384734 -6426
rect 384114 -7654 384734 -6662
rect 387834 29494 388454 43007
rect 387834 29258 387866 29494
rect 388102 29258 388186 29494
rect 388422 29258 388454 29494
rect 387834 29174 388454 29258
rect 387834 28938 387866 29174
rect 388102 28938 388186 29174
rect 388422 28938 388454 29174
rect 387834 -7066 388454 28938
rect 387834 -7302 387866 -7066
rect 388102 -7302 388186 -7066
rect 388422 -7302 388454 -7066
rect 387834 -7386 388454 -7302
rect 387834 -7622 387866 -7386
rect 388102 -7622 388186 -7386
rect 388422 -7622 388454 -7386
rect 387834 -7654 388454 -7622
rect 397794 39454 398414 43007
rect 397794 39218 397826 39454
rect 398062 39218 398146 39454
rect 398382 39218 398414 39454
rect 397794 39134 398414 39218
rect 397794 38898 397826 39134
rect 398062 38898 398146 39134
rect 398382 38898 398414 39134
rect 397794 3454 398414 38898
rect 397794 3218 397826 3454
rect 398062 3218 398146 3454
rect 398382 3218 398414 3454
rect 397794 3134 398414 3218
rect 397794 2898 397826 3134
rect 398062 2898 398146 3134
rect 398382 2898 398414 3134
rect 397794 -346 398414 2898
rect 397794 -582 397826 -346
rect 398062 -582 398146 -346
rect 398382 -582 398414 -346
rect 397794 -666 398414 -582
rect 397794 -902 397826 -666
rect 398062 -902 398146 -666
rect 398382 -902 398414 -666
rect 397794 -7654 398414 -902
rect 401514 7174 402134 43007
rect 402448 42938 402490 43174
rect 402726 42938 402768 43174
rect 433168 43174 433488 43206
rect 402448 42854 402768 42938
rect 402448 42618 402490 42854
rect 402726 42618 402768 42854
rect 402448 42586 402768 42618
rect 401514 6938 401546 7174
rect 401782 6938 401866 7174
rect 402102 6938 402134 7174
rect 401514 6854 402134 6938
rect 401514 6618 401546 6854
rect 401782 6618 401866 6854
rect 402102 6618 402134 6854
rect 401514 -1306 402134 6618
rect 401514 -1542 401546 -1306
rect 401782 -1542 401866 -1306
rect 402102 -1542 402134 -1306
rect 401514 -1626 402134 -1542
rect 401514 -1862 401546 -1626
rect 401782 -1862 401866 -1626
rect 402102 -1862 402134 -1626
rect 401514 -7654 402134 -1862
rect 405234 10894 405854 43007
rect 405234 10658 405266 10894
rect 405502 10658 405586 10894
rect 405822 10658 405854 10894
rect 405234 10574 405854 10658
rect 405234 10338 405266 10574
rect 405502 10338 405586 10574
rect 405822 10338 405854 10574
rect 405234 -2266 405854 10338
rect 405234 -2502 405266 -2266
rect 405502 -2502 405586 -2266
rect 405822 -2502 405854 -2266
rect 405234 -2586 405854 -2502
rect 405234 -2822 405266 -2586
rect 405502 -2822 405586 -2586
rect 405822 -2822 405854 -2586
rect 405234 -7654 405854 -2822
rect 408954 14614 409574 43007
rect 408954 14378 408986 14614
rect 409222 14378 409306 14614
rect 409542 14378 409574 14614
rect 408954 14294 409574 14378
rect 408954 14058 408986 14294
rect 409222 14058 409306 14294
rect 409542 14058 409574 14294
rect 408954 -3226 409574 14058
rect 408954 -3462 408986 -3226
rect 409222 -3462 409306 -3226
rect 409542 -3462 409574 -3226
rect 408954 -3546 409574 -3462
rect 408954 -3782 408986 -3546
rect 409222 -3782 409306 -3546
rect 409542 -3782 409574 -3546
rect 408954 -7654 409574 -3782
rect 412674 18334 413294 43007
rect 412674 18098 412706 18334
rect 412942 18098 413026 18334
rect 413262 18098 413294 18334
rect 412674 18014 413294 18098
rect 412674 17778 412706 18014
rect 412942 17778 413026 18014
rect 413262 17778 413294 18014
rect 412674 -4186 413294 17778
rect 412674 -4422 412706 -4186
rect 412942 -4422 413026 -4186
rect 413262 -4422 413294 -4186
rect 412674 -4506 413294 -4422
rect 412674 -4742 412706 -4506
rect 412942 -4742 413026 -4506
rect 413262 -4742 413294 -4506
rect 412674 -7654 413294 -4742
rect 416394 22054 417014 43007
rect 416394 21818 416426 22054
rect 416662 21818 416746 22054
rect 416982 21818 417014 22054
rect 416394 21734 417014 21818
rect 416394 21498 416426 21734
rect 416662 21498 416746 21734
rect 416982 21498 417014 21734
rect 416394 -5146 417014 21498
rect 416394 -5382 416426 -5146
rect 416662 -5382 416746 -5146
rect 416982 -5382 417014 -5146
rect 416394 -5466 417014 -5382
rect 416394 -5702 416426 -5466
rect 416662 -5702 416746 -5466
rect 416982 -5702 417014 -5466
rect 416394 -7654 417014 -5702
rect 420114 25774 420734 43007
rect 420114 25538 420146 25774
rect 420382 25538 420466 25774
rect 420702 25538 420734 25774
rect 420114 25454 420734 25538
rect 420114 25218 420146 25454
rect 420382 25218 420466 25454
rect 420702 25218 420734 25454
rect 420114 -6106 420734 25218
rect 420114 -6342 420146 -6106
rect 420382 -6342 420466 -6106
rect 420702 -6342 420734 -6106
rect 420114 -6426 420734 -6342
rect 420114 -6662 420146 -6426
rect 420382 -6662 420466 -6426
rect 420702 -6662 420734 -6426
rect 420114 -7654 420734 -6662
rect 423834 29494 424454 43007
rect 433168 42938 433210 43174
rect 433446 42938 433488 43174
rect 463888 43174 464208 43206
rect 433168 42854 433488 42938
rect 433168 42618 433210 42854
rect 433446 42618 433488 42854
rect 433168 42586 433488 42618
rect 423834 29258 423866 29494
rect 424102 29258 424186 29494
rect 424422 29258 424454 29494
rect 423834 29174 424454 29258
rect 423834 28938 423866 29174
rect 424102 28938 424186 29174
rect 424422 28938 424454 29174
rect 423834 -7066 424454 28938
rect 423834 -7302 423866 -7066
rect 424102 -7302 424186 -7066
rect 424422 -7302 424454 -7066
rect 423834 -7386 424454 -7302
rect 423834 -7622 423866 -7386
rect 424102 -7622 424186 -7386
rect 424422 -7622 424454 -7386
rect 423834 -7654 424454 -7622
rect 433794 39454 434414 43007
rect 433794 39218 433826 39454
rect 434062 39218 434146 39454
rect 434382 39218 434414 39454
rect 433794 39134 434414 39218
rect 433794 38898 433826 39134
rect 434062 38898 434146 39134
rect 434382 38898 434414 39134
rect 433794 3454 434414 38898
rect 433794 3218 433826 3454
rect 434062 3218 434146 3454
rect 434382 3218 434414 3454
rect 433794 3134 434414 3218
rect 433794 2898 433826 3134
rect 434062 2898 434146 3134
rect 434382 2898 434414 3134
rect 433794 -346 434414 2898
rect 433794 -582 433826 -346
rect 434062 -582 434146 -346
rect 434382 -582 434414 -346
rect 433794 -666 434414 -582
rect 433794 -902 433826 -666
rect 434062 -902 434146 -666
rect 434382 -902 434414 -666
rect 433794 -7654 434414 -902
rect 437514 7174 438134 43007
rect 437514 6938 437546 7174
rect 437782 6938 437866 7174
rect 438102 6938 438134 7174
rect 437514 6854 438134 6938
rect 437514 6618 437546 6854
rect 437782 6618 437866 6854
rect 438102 6618 438134 6854
rect 437514 -1306 438134 6618
rect 437514 -1542 437546 -1306
rect 437782 -1542 437866 -1306
rect 438102 -1542 438134 -1306
rect 437514 -1626 438134 -1542
rect 437514 -1862 437546 -1626
rect 437782 -1862 437866 -1626
rect 438102 -1862 438134 -1626
rect 437514 -7654 438134 -1862
rect 441234 10894 441854 43007
rect 441234 10658 441266 10894
rect 441502 10658 441586 10894
rect 441822 10658 441854 10894
rect 441234 10574 441854 10658
rect 441234 10338 441266 10574
rect 441502 10338 441586 10574
rect 441822 10338 441854 10574
rect 441234 -2266 441854 10338
rect 441234 -2502 441266 -2266
rect 441502 -2502 441586 -2266
rect 441822 -2502 441854 -2266
rect 441234 -2586 441854 -2502
rect 441234 -2822 441266 -2586
rect 441502 -2822 441586 -2586
rect 441822 -2822 441854 -2586
rect 441234 -7654 441854 -2822
rect 444954 14614 445574 43007
rect 444954 14378 444986 14614
rect 445222 14378 445306 14614
rect 445542 14378 445574 14614
rect 444954 14294 445574 14378
rect 444954 14058 444986 14294
rect 445222 14058 445306 14294
rect 445542 14058 445574 14294
rect 444954 -3226 445574 14058
rect 444954 -3462 444986 -3226
rect 445222 -3462 445306 -3226
rect 445542 -3462 445574 -3226
rect 444954 -3546 445574 -3462
rect 444954 -3782 444986 -3546
rect 445222 -3782 445306 -3546
rect 445542 -3782 445574 -3546
rect 444954 -7654 445574 -3782
rect 448674 18334 449294 40068
rect 448674 18098 448706 18334
rect 448942 18098 449026 18334
rect 449262 18098 449294 18334
rect 448674 18014 449294 18098
rect 448674 17778 448706 18014
rect 448942 17778 449026 18014
rect 449262 17778 449294 18014
rect 448674 -4186 449294 17778
rect 448674 -4422 448706 -4186
rect 448942 -4422 449026 -4186
rect 449262 -4422 449294 -4186
rect 448674 -4506 449294 -4422
rect 448674 -4742 448706 -4506
rect 448942 -4742 449026 -4506
rect 449262 -4742 449294 -4506
rect 448674 -7654 449294 -4742
rect 452394 22054 453014 43007
rect 452394 21818 452426 22054
rect 452662 21818 452746 22054
rect 452982 21818 453014 22054
rect 452394 21734 453014 21818
rect 452394 21498 452426 21734
rect 452662 21498 452746 21734
rect 452982 21498 453014 21734
rect 452394 -5146 453014 21498
rect 452394 -5382 452426 -5146
rect 452662 -5382 452746 -5146
rect 452982 -5382 453014 -5146
rect 452394 -5466 453014 -5382
rect 452394 -5702 452426 -5466
rect 452662 -5702 452746 -5466
rect 452982 -5702 453014 -5466
rect 452394 -7654 453014 -5702
rect 456114 25774 456734 43007
rect 456114 25538 456146 25774
rect 456382 25538 456466 25774
rect 456702 25538 456734 25774
rect 456114 25454 456734 25538
rect 456114 25218 456146 25454
rect 456382 25218 456466 25454
rect 456702 25218 456734 25454
rect 456114 -6106 456734 25218
rect 456114 -6342 456146 -6106
rect 456382 -6342 456466 -6106
rect 456702 -6342 456734 -6106
rect 456114 -6426 456734 -6342
rect 456114 -6662 456146 -6426
rect 456382 -6662 456466 -6426
rect 456702 -6662 456734 -6426
rect 456114 -7654 456734 -6662
rect 459834 29494 460454 43007
rect 463888 42938 463930 43174
rect 464166 42938 464208 43174
rect 494608 43174 494928 43206
rect 463888 42854 464208 42938
rect 463888 42618 463930 42854
rect 464166 42618 464208 42854
rect 463888 42586 464208 42618
rect 459834 29258 459866 29494
rect 460102 29258 460186 29494
rect 460422 29258 460454 29494
rect 459834 29174 460454 29258
rect 459834 28938 459866 29174
rect 460102 28938 460186 29174
rect 460422 28938 460454 29174
rect 459834 -7066 460454 28938
rect 459834 -7302 459866 -7066
rect 460102 -7302 460186 -7066
rect 460422 -7302 460454 -7066
rect 459834 -7386 460454 -7302
rect 459834 -7622 459866 -7386
rect 460102 -7622 460186 -7386
rect 460422 -7622 460454 -7386
rect 459834 -7654 460454 -7622
rect 469794 39454 470414 43007
rect 469794 39218 469826 39454
rect 470062 39218 470146 39454
rect 470382 39218 470414 39454
rect 469794 39134 470414 39218
rect 469794 38898 469826 39134
rect 470062 38898 470146 39134
rect 470382 38898 470414 39134
rect 469794 3454 470414 38898
rect 469794 3218 469826 3454
rect 470062 3218 470146 3454
rect 470382 3218 470414 3454
rect 469794 3134 470414 3218
rect 469794 2898 469826 3134
rect 470062 2898 470146 3134
rect 470382 2898 470414 3134
rect 469794 -346 470414 2898
rect 469794 -582 469826 -346
rect 470062 -582 470146 -346
rect 470382 -582 470414 -346
rect 469794 -666 470414 -582
rect 469794 -902 469826 -666
rect 470062 -902 470146 -666
rect 470382 -902 470414 -666
rect 469794 -7654 470414 -902
rect 473514 7174 474134 43007
rect 473514 6938 473546 7174
rect 473782 6938 473866 7174
rect 474102 6938 474134 7174
rect 473514 6854 474134 6938
rect 473514 6618 473546 6854
rect 473782 6618 473866 6854
rect 474102 6618 474134 6854
rect 473514 -1306 474134 6618
rect 473514 -1542 473546 -1306
rect 473782 -1542 473866 -1306
rect 474102 -1542 474134 -1306
rect 473514 -1626 474134 -1542
rect 473514 -1862 473546 -1626
rect 473782 -1862 473866 -1626
rect 474102 -1862 474134 -1626
rect 473514 -7654 474134 -1862
rect 477234 10894 477854 43007
rect 477234 10658 477266 10894
rect 477502 10658 477586 10894
rect 477822 10658 477854 10894
rect 477234 10574 477854 10658
rect 477234 10338 477266 10574
rect 477502 10338 477586 10574
rect 477822 10338 477854 10574
rect 477234 -2266 477854 10338
rect 477234 -2502 477266 -2266
rect 477502 -2502 477586 -2266
rect 477822 -2502 477854 -2266
rect 477234 -2586 477854 -2502
rect 477234 -2822 477266 -2586
rect 477502 -2822 477586 -2586
rect 477822 -2822 477854 -2586
rect 477234 -7654 477854 -2822
rect 480954 14614 481574 43007
rect 480954 14378 480986 14614
rect 481222 14378 481306 14614
rect 481542 14378 481574 14614
rect 480954 14294 481574 14378
rect 480954 14058 480986 14294
rect 481222 14058 481306 14294
rect 481542 14058 481574 14294
rect 480954 -3226 481574 14058
rect 480954 -3462 480986 -3226
rect 481222 -3462 481306 -3226
rect 481542 -3462 481574 -3226
rect 480954 -3546 481574 -3462
rect 480954 -3782 480986 -3546
rect 481222 -3782 481306 -3546
rect 481542 -3782 481574 -3546
rect 480954 -7654 481574 -3782
rect 484674 18334 485294 43007
rect 484674 18098 484706 18334
rect 484942 18098 485026 18334
rect 485262 18098 485294 18334
rect 484674 18014 485294 18098
rect 484674 17778 484706 18014
rect 484942 17778 485026 18014
rect 485262 17778 485294 18014
rect 484674 -4186 485294 17778
rect 484674 -4422 484706 -4186
rect 484942 -4422 485026 -4186
rect 485262 -4422 485294 -4186
rect 484674 -4506 485294 -4422
rect 484674 -4742 484706 -4506
rect 484942 -4742 485026 -4506
rect 485262 -4742 485294 -4506
rect 484674 -7654 485294 -4742
rect 488394 22054 489014 43007
rect 488394 21818 488426 22054
rect 488662 21818 488746 22054
rect 488982 21818 489014 22054
rect 488394 21734 489014 21818
rect 488394 21498 488426 21734
rect 488662 21498 488746 21734
rect 488982 21498 489014 21734
rect 488394 -5146 489014 21498
rect 488394 -5382 488426 -5146
rect 488662 -5382 488746 -5146
rect 488982 -5382 489014 -5146
rect 488394 -5466 489014 -5382
rect 488394 -5702 488426 -5466
rect 488662 -5702 488746 -5466
rect 488982 -5702 489014 -5466
rect 488394 -7654 489014 -5702
rect 492114 25774 492734 43007
rect 494608 42938 494650 43174
rect 494886 42938 494928 43174
rect 525328 43174 525648 43206
rect 494608 42854 494928 42938
rect 494608 42618 494650 42854
rect 494886 42618 494928 42854
rect 494608 42586 494928 42618
rect 492114 25538 492146 25774
rect 492382 25538 492466 25774
rect 492702 25538 492734 25774
rect 492114 25454 492734 25538
rect 492114 25218 492146 25454
rect 492382 25218 492466 25454
rect 492702 25218 492734 25454
rect 492114 -6106 492734 25218
rect 492114 -6342 492146 -6106
rect 492382 -6342 492466 -6106
rect 492702 -6342 492734 -6106
rect 492114 -6426 492734 -6342
rect 492114 -6662 492146 -6426
rect 492382 -6662 492466 -6426
rect 492702 -6662 492734 -6426
rect 492114 -7654 492734 -6662
rect 495834 29494 496454 43007
rect 495834 29258 495866 29494
rect 496102 29258 496186 29494
rect 496422 29258 496454 29494
rect 495834 29174 496454 29258
rect 495834 28938 495866 29174
rect 496102 28938 496186 29174
rect 496422 28938 496454 29174
rect 495834 -7066 496454 28938
rect 495834 -7302 495866 -7066
rect 496102 -7302 496186 -7066
rect 496422 -7302 496454 -7066
rect 495834 -7386 496454 -7302
rect 495834 -7622 495866 -7386
rect 496102 -7622 496186 -7386
rect 496422 -7622 496454 -7386
rect 495834 -7654 496454 -7622
rect 505794 39454 506414 43007
rect 505794 39218 505826 39454
rect 506062 39218 506146 39454
rect 506382 39218 506414 39454
rect 505794 39134 506414 39218
rect 505794 38898 505826 39134
rect 506062 38898 506146 39134
rect 506382 38898 506414 39134
rect 505794 3454 506414 38898
rect 505794 3218 505826 3454
rect 506062 3218 506146 3454
rect 506382 3218 506414 3454
rect 505794 3134 506414 3218
rect 505794 2898 505826 3134
rect 506062 2898 506146 3134
rect 506382 2898 506414 3134
rect 505794 -346 506414 2898
rect 505794 -582 505826 -346
rect 506062 -582 506146 -346
rect 506382 -582 506414 -346
rect 505794 -666 506414 -582
rect 505794 -902 505826 -666
rect 506062 -902 506146 -666
rect 506382 -902 506414 -666
rect 505794 -7654 506414 -902
rect 509514 7174 510134 40068
rect 509514 6938 509546 7174
rect 509782 6938 509866 7174
rect 510102 6938 510134 7174
rect 509514 6854 510134 6938
rect 509514 6618 509546 6854
rect 509782 6618 509866 6854
rect 510102 6618 510134 6854
rect 509514 -1306 510134 6618
rect 509514 -1542 509546 -1306
rect 509782 -1542 509866 -1306
rect 510102 -1542 510134 -1306
rect 509514 -1626 510134 -1542
rect 509514 -1862 509546 -1626
rect 509782 -1862 509866 -1626
rect 510102 -1862 510134 -1626
rect 509514 -7654 510134 -1862
rect 513234 10894 513854 43007
rect 513234 10658 513266 10894
rect 513502 10658 513586 10894
rect 513822 10658 513854 10894
rect 513234 10574 513854 10658
rect 513234 10338 513266 10574
rect 513502 10338 513586 10574
rect 513822 10338 513854 10574
rect 513234 -2266 513854 10338
rect 513234 -2502 513266 -2266
rect 513502 -2502 513586 -2266
rect 513822 -2502 513854 -2266
rect 513234 -2586 513854 -2502
rect 513234 -2822 513266 -2586
rect 513502 -2822 513586 -2586
rect 513822 -2822 513854 -2586
rect 513234 -7654 513854 -2822
rect 516954 14614 517574 43007
rect 516954 14378 516986 14614
rect 517222 14378 517306 14614
rect 517542 14378 517574 14614
rect 516954 14294 517574 14378
rect 516954 14058 516986 14294
rect 517222 14058 517306 14294
rect 517542 14058 517574 14294
rect 516954 -3226 517574 14058
rect 516954 -3462 516986 -3226
rect 517222 -3462 517306 -3226
rect 517542 -3462 517574 -3226
rect 516954 -3546 517574 -3462
rect 516954 -3782 516986 -3546
rect 517222 -3782 517306 -3546
rect 517542 -3782 517574 -3546
rect 516954 -7654 517574 -3782
rect 520674 18334 521294 43007
rect 520674 18098 520706 18334
rect 520942 18098 521026 18334
rect 521262 18098 521294 18334
rect 520674 18014 521294 18098
rect 520674 17778 520706 18014
rect 520942 17778 521026 18014
rect 521262 17778 521294 18014
rect 520674 -4186 521294 17778
rect 520674 -4422 520706 -4186
rect 520942 -4422 521026 -4186
rect 521262 -4422 521294 -4186
rect 520674 -4506 521294 -4422
rect 520674 -4742 520706 -4506
rect 520942 -4742 521026 -4506
rect 521262 -4742 521294 -4506
rect 520674 -7654 521294 -4742
rect 524394 22054 525014 43007
rect 525328 42938 525370 43174
rect 525606 42938 525648 43174
rect 525328 42854 525648 42938
rect 525328 42618 525370 42854
rect 525606 42618 525648 42854
rect 525328 42586 525648 42618
rect 524394 21818 524426 22054
rect 524662 21818 524746 22054
rect 524982 21818 525014 22054
rect 524394 21734 525014 21818
rect 524394 21498 524426 21734
rect 524662 21498 524746 21734
rect 524982 21498 525014 21734
rect 524394 -5146 525014 21498
rect 524394 -5382 524426 -5146
rect 524662 -5382 524746 -5146
rect 524982 -5382 525014 -5146
rect 524394 -5466 525014 -5382
rect 524394 -5702 524426 -5466
rect 524662 -5702 524746 -5466
rect 524982 -5702 525014 -5466
rect 524394 -7654 525014 -5702
rect 528114 25774 528734 43007
rect 528114 25538 528146 25774
rect 528382 25538 528466 25774
rect 528702 25538 528734 25774
rect 528114 25454 528734 25538
rect 528114 25218 528146 25454
rect 528382 25218 528466 25454
rect 528702 25218 528734 25454
rect 528114 -6106 528734 25218
rect 528114 -6342 528146 -6106
rect 528382 -6342 528466 -6106
rect 528702 -6342 528734 -6106
rect 528114 -6426 528734 -6342
rect 528114 -6662 528146 -6426
rect 528382 -6662 528466 -6426
rect 528702 -6662 528734 -6426
rect 528114 -7654 528734 -6662
rect 531834 29494 532454 43007
rect 531834 29258 531866 29494
rect 532102 29258 532186 29494
rect 532422 29258 532454 29494
rect 531834 29174 532454 29258
rect 531834 28938 531866 29174
rect 532102 28938 532186 29174
rect 532422 28938 532454 29174
rect 531834 -7066 532454 28938
rect 531834 -7302 531866 -7066
rect 532102 -7302 532186 -7066
rect 532422 -7302 532454 -7066
rect 531834 -7386 532454 -7302
rect 531834 -7622 531866 -7386
rect 532102 -7622 532186 -7386
rect 532422 -7622 532454 -7386
rect 531834 -7654 532454 -7622
rect 541794 39454 542414 43007
rect 541794 39218 541826 39454
rect 542062 39218 542146 39454
rect 542382 39218 542414 39454
rect 541794 39134 542414 39218
rect 541794 38898 541826 39134
rect 542062 38898 542146 39134
rect 542382 38898 542414 39134
rect 541794 3454 542414 38898
rect 541794 3218 541826 3454
rect 542062 3218 542146 3454
rect 542382 3218 542414 3454
rect 541794 3134 542414 3218
rect 541794 2898 541826 3134
rect 542062 2898 542146 3134
rect 542382 2898 542414 3134
rect 541794 -346 542414 2898
rect 541794 -582 541826 -346
rect 542062 -582 542146 -346
rect 542382 -582 542414 -346
rect 541794 -666 542414 -582
rect 541794 -902 541826 -666
rect 542062 -902 542146 -666
rect 542382 -902 542414 -666
rect 541794 -7654 542414 -902
rect 545514 7174 546134 43007
rect 545514 6938 545546 7174
rect 545782 6938 545866 7174
rect 546102 6938 546134 7174
rect 545514 6854 546134 6938
rect 545514 6618 545546 6854
rect 545782 6618 545866 6854
rect 546102 6618 546134 6854
rect 545514 -1306 546134 6618
rect 545514 -1542 545546 -1306
rect 545782 -1542 545866 -1306
rect 546102 -1542 546134 -1306
rect 545514 -1626 546134 -1542
rect 545514 -1862 545546 -1626
rect 545782 -1862 545866 -1626
rect 546102 -1862 546134 -1626
rect 545514 -7654 546134 -1862
rect 549234 10894 549854 43007
rect 549234 10658 549266 10894
rect 549502 10658 549586 10894
rect 549822 10658 549854 10894
rect 549234 10574 549854 10658
rect 549234 10338 549266 10574
rect 549502 10338 549586 10574
rect 549822 10338 549854 10574
rect 549234 -2266 549854 10338
rect 549234 -2502 549266 -2266
rect 549502 -2502 549586 -2266
rect 549822 -2502 549854 -2266
rect 549234 -2586 549854 -2502
rect 549234 -2822 549266 -2586
rect 549502 -2822 549586 -2586
rect 549822 -2822 549854 -2586
rect 549234 -7654 549854 -2822
rect 552954 14614 553574 50058
rect 552954 14378 552986 14614
rect 553222 14378 553306 14614
rect 553542 14378 553574 14614
rect 552954 14294 553574 14378
rect 552954 14058 552986 14294
rect 553222 14058 553306 14294
rect 553542 14058 553574 14294
rect 552954 -3226 553574 14058
rect 552954 -3462 552986 -3226
rect 553222 -3462 553306 -3226
rect 553542 -3462 553574 -3226
rect 552954 -3546 553574 -3462
rect 552954 -3782 552986 -3546
rect 553222 -3782 553306 -3546
rect 553542 -3782 553574 -3546
rect 552954 -7654 553574 -3782
rect 556674 708678 557294 711590
rect 556674 708442 556706 708678
rect 556942 708442 557026 708678
rect 557262 708442 557294 708678
rect 556674 708358 557294 708442
rect 556674 708122 556706 708358
rect 556942 708122 557026 708358
rect 557262 708122 557294 708358
rect 556674 666334 557294 708122
rect 556674 666098 556706 666334
rect 556942 666098 557026 666334
rect 557262 666098 557294 666334
rect 556674 666014 557294 666098
rect 556674 665778 556706 666014
rect 556942 665778 557026 666014
rect 557262 665778 557294 666014
rect 556674 630334 557294 665778
rect 556674 630098 556706 630334
rect 556942 630098 557026 630334
rect 557262 630098 557294 630334
rect 556674 630014 557294 630098
rect 556674 629778 556706 630014
rect 556942 629778 557026 630014
rect 557262 629778 557294 630014
rect 556674 594334 557294 629778
rect 556674 594098 556706 594334
rect 556942 594098 557026 594334
rect 557262 594098 557294 594334
rect 556674 594014 557294 594098
rect 556674 593778 556706 594014
rect 556942 593778 557026 594014
rect 557262 593778 557294 594014
rect 556674 558334 557294 593778
rect 556674 558098 556706 558334
rect 556942 558098 557026 558334
rect 557262 558098 557294 558334
rect 556674 558014 557294 558098
rect 556674 557778 556706 558014
rect 556942 557778 557026 558014
rect 557262 557778 557294 558014
rect 556674 522334 557294 557778
rect 556674 522098 556706 522334
rect 556942 522098 557026 522334
rect 557262 522098 557294 522334
rect 556674 522014 557294 522098
rect 556674 521778 556706 522014
rect 556942 521778 557026 522014
rect 557262 521778 557294 522014
rect 556674 486334 557294 521778
rect 556674 486098 556706 486334
rect 556942 486098 557026 486334
rect 557262 486098 557294 486334
rect 556674 486014 557294 486098
rect 556674 485778 556706 486014
rect 556942 485778 557026 486014
rect 557262 485778 557294 486014
rect 556674 450334 557294 485778
rect 556674 450098 556706 450334
rect 556942 450098 557026 450334
rect 557262 450098 557294 450334
rect 556674 450014 557294 450098
rect 556674 449778 556706 450014
rect 556942 449778 557026 450014
rect 557262 449778 557294 450014
rect 556674 414334 557294 449778
rect 556674 414098 556706 414334
rect 556942 414098 557026 414334
rect 557262 414098 557294 414334
rect 556674 414014 557294 414098
rect 556674 413778 556706 414014
rect 556942 413778 557026 414014
rect 557262 413778 557294 414014
rect 556674 378334 557294 413778
rect 556674 378098 556706 378334
rect 556942 378098 557026 378334
rect 557262 378098 557294 378334
rect 556674 378014 557294 378098
rect 556674 377778 556706 378014
rect 556942 377778 557026 378014
rect 557262 377778 557294 378014
rect 556674 342334 557294 377778
rect 556674 342098 556706 342334
rect 556942 342098 557026 342334
rect 557262 342098 557294 342334
rect 556674 342014 557294 342098
rect 556674 341778 556706 342014
rect 556942 341778 557026 342014
rect 557262 341778 557294 342014
rect 556674 306334 557294 341778
rect 556674 306098 556706 306334
rect 556942 306098 557026 306334
rect 557262 306098 557294 306334
rect 556674 306014 557294 306098
rect 556674 305778 556706 306014
rect 556942 305778 557026 306014
rect 557262 305778 557294 306014
rect 556674 270334 557294 305778
rect 556674 270098 556706 270334
rect 556942 270098 557026 270334
rect 557262 270098 557294 270334
rect 556674 270014 557294 270098
rect 556674 269778 556706 270014
rect 556942 269778 557026 270014
rect 557262 269778 557294 270014
rect 556674 234334 557294 269778
rect 556674 234098 556706 234334
rect 556942 234098 557026 234334
rect 557262 234098 557294 234334
rect 556674 234014 557294 234098
rect 556674 233778 556706 234014
rect 556942 233778 557026 234014
rect 557262 233778 557294 234014
rect 556674 198334 557294 233778
rect 556674 198098 556706 198334
rect 556942 198098 557026 198334
rect 557262 198098 557294 198334
rect 556674 198014 557294 198098
rect 556674 197778 556706 198014
rect 556942 197778 557026 198014
rect 557262 197778 557294 198014
rect 556674 162334 557294 197778
rect 556674 162098 556706 162334
rect 556942 162098 557026 162334
rect 557262 162098 557294 162334
rect 556674 162014 557294 162098
rect 556674 161778 556706 162014
rect 556942 161778 557026 162014
rect 557262 161778 557294 162014
rect 556674 126334 557294 161778
rect 556674 126098 556706 126334
rect 556942 126098 557026 126334
rect 557262 126098 557294 126334
rect 556674 126014 557294 126098
rect 556674 125778 556706 126014
rect 556942 125778 557026 126014
rect 557262 125778 557294 126014
rect 556674 90334 557294 125778
rect 556674 90098 556706 90334
rect 556942 90098 557026 90334
rect 557262 90098 557294 90334
rect 556674 90014 557294 90098
rect 556674 89778 556706 90014
rect 556942 89778 557026 90014
rect 557262 89778 557294 90014
rect 556674 54334 557294 89778
rect 556674 54098 556706 54334
rect 556942 54098 557026 54334
rect 557262 54098 557294 54334
rect 556674 54014 557294 54098
rect 556674 53778 556706 54014
rect 556942 53778 557026 54014
rect 557262 53778 557294 54014
rect 556674 18334 557294 53778
rect 556674 18098 556706 18334
rect 556942 18098 557026 18334
rect 557262 18098 557294 18334
rect 556674 18014 557294 18098
rect 556674 17778 556706 18014
rect 556942 17778 557026 18014
rect 557262 17778 557294 18014
rect 556674 -4186 557294 17778
rect 556674 -4422 556706 -4186
rect 556942 -4422 557026 -4186
rect 557262 -4422 557294 -4186
rect 556674 -4506 557294 -4422
rect 556674 -4742 556706 -4506
rect 556942 -4742 557026 -4506
rect 557262 -4742 557294 -4506
rect 556674 -7654 557294 -4742
rect 560394 709638 561014 711590
rect 560394 709402 560426 709638
rect 560662 709402 560746 709638
rect 560982 709402 561014 709638
rect 560394 709318 561014 709402
rect 560394 709082 560426 709318
rect 560662 709082 560746 709318
rect 560982 709082 561014 709318
rect 560394 670054 561014 709082
rect 560394 669818 560426 670054
rect 560662 669818 560746 670054
rect 560982 669818 561014 670054
rect 560394 669734 561014 669818
rect 560394 669498 560426 669734
rect 560662 669498 560746 669734
rect 560982 669498 561014 669734
rect 560394 634054 561014 669498
rect 560394 633818 560426 634054
rect 560662 633818 560746 634054
rect 560982 633818 561014 634054
rect 560394 633734 561014 633818
rect 560394 633498 560426 633734
rect 560662 633498 560746 633734
rect 560982 633498 561014 633734
rect 560394 598054 561014 633498
rect 560394 597818 560426 598054
rect 560662 597818 560746 598054
rect 560982 597818 561014 598054
rect 560394 597734 561014 597818
rect 560394 597498 560426 597734
rect 560662 597498 560746 597734
rect 560982 597498 561014 597734
rect 560394 562054 561014 597498
rect 560394 561818 560426 562054
rect 560662 561818 560746 562054
rect 560982 561818 561014 562054
rect 560394 561734 561014 561818
rect 560394 561498 560426 561734
rect 560662 561498 560746 561734
rect 560982 561498 561014 561734
rect 560394 526054 561014 561498
rect 560394 525818 560426 526054
rect 560662 525818 560746 526054
rect 560982 525818 561014 526054
rect 560394 525734 561014 525818
rect 560394 525498 560426 525734
rect 560662 525498 560746 525734
rect 560982 525498 561014 525734
rect 560394 490054 561014 525498
rect 560394 489818 560426 490054
rect 560662 489818 560746 490054
rect 560982 489818 561014 490054
rect 560394 489734 561014 489818
rect 560394 489498 560426 489734
rect 560662 489498 560746 489734
rect 560982 489498 561014 489734
rect 560394 454054 561014 489498
rect 560394 453818 560426 454054
rect 560662 453818 560746 454054
rect 560982 453818 561014 454054
rect 560394 453734 561014 453818
rect 560394 453498 560426 453734
rect 560662 453498 560746 453734
rect 560982 453498 561014 453734
rect 560394 418054 561014 453498
rect 560394 417818 560426 418054
rect 560662 417818 560746 418054
rect 560982 417818 561014 418054
rect 560394 417734 561014 417818
rect 560394 417498 560426 417734
rect 560662 417498 560746 417734
rect 560982 417498 561014 417734
rect 560394 382054 561014 417498
rect 560394 381818 560426 382054
rect 560662 381818 560746 382054
rect 560982 381818 561014 382054
rect 560394 381734 561014 381818
rect 560394 381498 560426 381734
rect 560662 381498 560746 381734
rect 560982 381498 561014 381734
rect 560394 346054 561014 381498
rect 560394 345818 560426 346054
rect 560662 345818 560746 346054
rect 560982 345818 561014 346054
rect 560394 345734 561014 345818
rect 560394 345498 560426 345734
rect 560662 345498 560746 345734
rect 560982 345498 561014 345734
rect 560394 310054 561014 345498
rect 560394 309818 560426 310054
rect 560662 309818 560746 310054
rect 560982 309818 561014 310054
rect 560394 309734 561014 309818
rect 560394 309498 560426 309734
rect 560662 309498 560746 309734
rect 560982 309498 561014 309734
rect 560394 274054 561014 309498
rect 560394 273818 560426 274054
rect 560662 273818 560746 274054
rect 560982 273818 561014 274054
rect 560394 273734 561014 273818
rect 560394 273498 560426 273734
rect 560662 273498 560746 273734
rect 560982 273498 561014 273734
rect 560394 238054 561014 273498
rect 560394 237818 560426 238054
rect 560662 237818 560746 238054
rect 560982 237818 561014 238054
rect 560394 237734 561014 237818
rect 560394 237498 560426 237734
rect 560662 237498 560746 237734
rect 560982 237498 561014 237734
rect 560394 202054 561014 237498
rect 560394 201818 560426 202054
rect 560662 201818 560746 202054
rect 560982 201818 561014 202054
rect 560394 201734 561014 201818
rect 560394 201498 560426 201734
rect 560662 201498 560746 201734
rect 560982 201498 561014 201734
rect 560394 166054 561014 201498
rect 560394 165818 560426 166054
rect 560662 165818 560746 166054
rect 560982 165818 561014 166054
rect 560394 165734 561014 165818
rect 560394 165498 560426 165734
rect 560662 165498 560746 165734
rect 560982 165498 561014 165734
rect 560394 130054 561014 165498
rect 560394 129818 560426 130054
rect 560662 129818 560746 130054
rect 560982 129818 561014 130054
rect 560394 129734 561014 129818
rect 560394 129498 560426 129734
rect 560662 129498 560746 129734
rect 560982 129498 561014 129734
rect 560394 94054 561014 129498
rect 560394 93818 560426 94054
rect 560662 93818 560746 94054
rect 560982 93818 561014 94054
rect 560394 93734 561014 93818
rect 560394 93498 560426 93734
rect 560662 93498 560746 93734
rect 560982 93498 561014 93734
rect 560394 58054 561014 93498
rect 560394 57818 560426 58054
rect 560662 57818 560746 58054
rect 560982 57818 561014 58054
rect 560394 57734 561014 57818
rect 560394 57498 560426 57734
rect 560662 57498 560746 57734
rect 560982 57498 561014 57734
rect 560394 22054 561014 57498
rect 560394 21818 560426 22054
rect 560662 21818 560746 22054
rect 560982 21818 561014 22054
rect 560394 21734 561014 21818
rect 560394 21498 560426 21734
rect 560662 21498 560746 21734
rect 560982 21498 561014 21734
rect 560394 -5146 561014 21498
rect 560394 -5382 560426 -5146
rect 560662 -5382 560746 -5146
rect 560982 -5382 561014 -5146
rect 560394 -5466 561014 -5382
rect 560394 -5702 560426 -5466
rect 560662 -5702 560746 -5466
rect 560982 -5702 561014 -5466
rect 560394 -7654 561014 -5702
rect 564114 710598 564734 711590
rect 564114 710362 564146 710598
rect 564382 710362 564466 710598
rect 564702 710362 564734 710598
rect 564114 710278 564734 710362
rect 564114 710042 564146 710278
rect 564382 710042 564466 710278
rect 564702 710042 564734 710278
rect 564114 673774 564734 710042
rect 564114 673538 564146 673774
rect 564382 673538 564466 673774
rect 564702 673538 564734 673774
rect 564114 673454 564734 673538
rect 564114 673218 564146 673454
rect 564382 673218 564466 673454
rect 564702 673218 564734 673454
rect 564114 637774 564734 673218
rect 564114 637538 564146 637774
rect 564382 637538 564466 637774
rect 564702 637538 564734 637774
rect 564114 637454 564734 637538
rect 564114 637218 564146 637454
rect 564382 637218 564466 637454
rect 564702 637218 564734 637454
rect 564114 601774 564734 637218
rect 567834 711558 568454 711590
rect 567834 711322 567866 711558
rect 568102 711322 568186 711558
rect 568422 711322 568454 711558
rect 567834 711238 568454 711322
rect 567834 711002 567866 711238
rect 568102 711002 568186 711238
rect 568422 711002 568454 711238
rect 567834 677494 568454 711002
rect 567834 677258 567866 677494
rect 568102 677258 568186 677494
rect 568422 677258 568454 677494
rect 567834 677174 568454 677258
rect 567834 676938 567866 677174
rect 568102 676938 568186 677174
rect 568422 676938 568454 677174
rect 567834 641494 568454 676938
rect 567834 641258 567866 641494
rect 568102 641258 568186 641494
rect 568422 641258 568454 641494
rect 567834 641174 568454 641258
rect 567834 640938 567866 641174
rect 568102 640938 568186 641174
rect 568422 640938 568454 641174
rect 565008 615454 565328 615486
rect 565008 615218 565050 615454
rect 565286 615218 565328 615454
rect 565008 615134 565328 615218
rect 565008 614898 565050 615134
rect 565286 614898 565328 615134
rect 565008 614866 565328 614898
rect 564114 601538 564146 601774
rect 564382 601538 564466 601774
rect 564702 601538 564734 601774
rect 564114 601454 564734 601538
rect 564114 601218 564146 601454
rect 564382 601218 564466 601454
rect 564702 601218 564734 601454
rect 564114 565774 564734 601218
rect 567834 605494 568454 640938
rect 567834 605258 567866 605494
rect 568102 605258 568186 605494
rect 568422 605258 568454 605494
rect 567834 605174 568454 605258
rect 567834 604938 567866 605174
rect 568102 604938 568186 605174
rect 568422 604938 568454 605174
rect 565008 579454 565328 579486
rect 565008 579218 565050 579454
rect 565286 579218 565328 579454
rect 565008 579134 565328 579218
rect 565008 578898 565050 579134
rect 565286 578898 565328 579134
rect 565008 578866 565328 578898
rect 564114 565538 564146 565774
rect 564382 565538 564466 565774
rect 564702 565538 564734 565774
rect 564114 565454 564734 565538
rect 564114 565218 564146 565454
rect 564382 565218 564466 565454
rect 564702 565218 564734 565454
rect 564114 529774 564734 565218
rect 567834 569494 568454 604938
rect 567834 569258 567866 569494
rect 568102 569258 568186 569494
rect 568422 569258 568454 569494
rect 567834 569174 568454 569258
rect 567834 568938 567866 569174
rect 568102 568938 568186 569174
rect 568422 568938 568454 569174
rect 565008 543454 565328 543486
rect 565008 543218 565050 543454
rect 565286 543218 565328 543454
rect 565008 543134 565328 543218
rect 565008 542898 565050 543134
rect 565286 542898 565328 543134
rect 565008 542866 565328 542898
rect 564114 529538 564146 529774
rect 564382 529538 564466 529774
rect 564702 529538 564734 529774
rect 564114 529454 564734 529538
rect 564114 529218 564146 529454
rect 564382 529218 564466 529454
rect 564702 529218 564734 529454
rect 564114 493774 564734 529218
rect 564114 493538 564146 493774
rect 564382 493538 564466 493774
rect 564702 493538 564734 493774
rect 564114 493454 564734 493538
rect 564114 493218 564146 493454
rect 564382 493218 564466 493454
rect 564702 493218 564734 493454
rect 564114 457774 564734 493218
rect 567834 533494 568454 568938
rect 567834 533258 567866 533494
rect 568102 533258 568186 533494
rect 568422 533258 568454 533494
rect 567834 533174 568454 533258
rect 567834 532938 567866 533174
rect 568102 532938 568186 533174
rect 568422 532938 568454 533174
rect 567834 497494 568454 532938
rect 567834 497258 567866 497494
rect 568102 497258 568186 497494
rect 568422 497258 568454 497494
rect 567834 497174 568454 497258
rect 567834 496938 567866 497174
rect 568102 496938 568186 497174
rect 568422 496938 568454 497174
rect 565008 471454 565328 471486
rect 565008 471218 565050 471454
rect 565286 471218 565328 471454
rect 565008 471134 565328 471218
rect 565008 470898 565050 471134
rect 565286 470898 565328 471134
rect 565008 470866 565328 470898
rect 564114 457538 564146 457774
rect 564382 457538 564466 457774
rect 564702 457538 564734 457774
rect 564114 457454 564734 457538
rect 564114 457218 564146 457454
rect 564382 457218 564466 457454
rect 564702 457218 564734 457454
rect 564114 421774 564734 457218
rect 567834 461494 568454 496938
rect 567834 461258 567866 461494
rect 568102 461258 568186 461494
rect 568422 461258 568454 461494
rect 567834 461174 568454 461258
rect 567834 460938 567866 461174
rect 568102 460938 568186 461174
rect 568422 460938 568454 461174
rect 565008 435454 565328 435486
rect 565008 435218 565050 435454
rect 565286 435218 565328 435454
rect 565008 435134 565328 435218
rect 565008 434898 565050 435134
rect 565286 434898 565328 435134
rect 565008 434866 565328 434898
rect 564114 421538 564146 421774
rect 564382 421538 564466 421774
rect 564702 421538 564734 421774
rect 564114 421454 564734 421538
rect 564114 421218 564146 421454
rect 564382 421218 564466 421454
rect 564702 421218 564734 421454
rect 564114 385774 564734 421218
rect 567834 425494 568454 460938
rect 567834 425258 567866 425494
rect 568102 425258 568186 425494
rect 568422 425258 568454 425494
rect 567834 425174 568454 425258
rect 567834 424938 567866 425174
rect 568102 424938 568186 425174
rect 568422 424938 568454 425174
rect 565008 399454 565328 399486
rect 565008 399218 565050 399454
rect 565286 399218 565328 399454
rect 565008 399134 565328 399218
rect 565008 398898 565050 399134
rect 565286 398898 565328 399134
rect 565008 398866 565328 398898
rect 564114 385538 564146 385774
rect 564382 385538 564466 385774
rect 564702 385538 564734 385774
rect 564114 385454 564734 385538
rect 564114 385218 564146 385454
rect 564382 385218 564466 385454
rect 564702 385218 564734 385454
rect 564114 349774 564734 385218
rect 564114 349538 564146 349774
rect 564382 349538 564466 349774
rect 564702 349538 564734 349774
rect 564114 349454 564734 349538
rect 564114 349218 564146 349454
rect 564382 349218 564466 349454
rect 564702 349218 564734 349454
rect 564114 313774 564734 349218
rect 564114 313538 564146 313774
rect 564382 313538 564466 313774
rect 564702 313538 564734 313774
rect 564114 313454 564734 313538
rect 564114 313218 564146 313454
rect 564382 313218 564466 313454
rect 564702 313218 564734 313454
rect 564114 277774 564734 313218
rect 564114 277538 564146 277774
rect 564382 277538 564466 277774
rect 564702 277538 564734 277774
rect 564114 277454 564734 277538
rect 564114 277218 564146 277454
rect 564382 277218 564466 277454
rect 564702 277218 564734 277454
rect 564114 241774 564734 277218
rect 564114 241538 564146 241774
rect 564382 241538 564466 241774
rect 564702 241538 564734 241774
rect 564114 241454 564734 241538
rect 564114 241218 564146 241454
rect 564382 241218 564466 241454
rect 564702 241218 564734 241454
rect 564114 205774 564734 241218
rect 564114 205538 564146 205774
rect 564382 205538 564466 205774
rect 564702 205538 564734 205774
rect 564114 205454 564734 205538
rect 564114 205218 564146 205454
rect 564382 205218 564466 205454
rect 564702 205218 564734 205454
rect 564114 169774 564734 205218
rect 564114 169538 564146 169774
rect 564382 169538 564466 169774
rect 564702 169538 564734 169774
rect 564114 169454 564734 169538
rect 564114 169218 564146 169454
rect 564382 169218 564466 169454
rect 564702 169218 564734 169454
rect 564114 133774 564734 169218
rect 564114 133538 564146 133774
rect 564382 133538 564466 133774
rect 564702 133538 564734 133774
rect 564114 133454 564734 133538
rect 564114 133218 564146 133454
rect 564382 133218 564466 133454
rect 564702 133218 564734 133454
rect 564114 97774 564734 133218
rect 564114 97538 564146 97774
rect 564382 97538 564466 97774
rect 564702 97538 564734 97774
rect 564114 97454 564734 97538
rect 564114 97218 564146 97454
rect 564382 97218 564466 97454
rect 564702 97218 564734 97454
rect 564114 61774 564734 97218
rect 564114 61538 564146 61774
rect 564382 61538 564466 61774
rect 564702 61538 564734 61774
rect 564114 61454 564734 61538
rect 564114 61218 564146 61454
rect 564382 61218 564466 61454
rect 564702 61218 564734 61454
rect 564114 25774 564734 61218
rect 564114 25538 564146 25774
rect 564382 25538 564466 25774
rect 564702 25538 564734 25774
rect 564114 25454 564734 25538
rect 564114 25218 564146 25454
rect 564382 25218 564466 25454
rect 564702 25218 564734 25454
rect 564114 -6106 564734 25218
rect 564114 -6342 564146 -6106
rect 564382 -6342 564466 -6106
rect 564702 -6342 564734 -6106
rect 564114 -6426 564734 -6342
rect 564114 -6662 564146 -6426
rect 564382 -6662 564466 -6426
rect 564702 -6662 564734 -6426
rect 564114 -7654 564734 -6662
rect 567834 389494 568454 424938
rect 567834 389258 567866 389494
rect 568102 389258 568186 389494
rect 568422 389258 568454 389494
rect 567834 389174 568454 389258
rect 567834 388938 567866 389174
rect 568102 388938 568186 389174
rect 568422 388938 568454 389174
rect 567834 353494 568454 388938
rect 567834 353258 567866 353494
rect 568102 353258 568186 353494
rect 568422 353258 568454 353494
rect 567834 353174 568454 353258
rect 567834 352938 567866 353174
rect 568102 352938 568186 353174
rect 568422 352938 568454 353174
rect 567834 317494 568454 352938
rect 567834 317258 567866 317494
rect 568102 317258 568186 317494
rect 568422 317258 568454 317494
rect 567834 317174 568454 317258
rect 567834 316938 567866 317174
rect 568102 316938 568186 317174
rect 568422 316938 568454 317174
rect 567834 281494 568454 316938
rect 567834 281258 567866 281494
rect 568102 281258 568186 281494
rect 568422 281258 568454 281494
rect 567834 281174 568454 281258
rect 567834 280938 567866 281174
rect 568102 280938 568186 281174
rect 568422 280938 568454 281174
rect 567834 245494 568454 280938
rect 567834 245258 567866 245494
rect 568102 245258 568186 245494
rect 568422 245258 568454 245494
rect 567834 245174 568454 245258
rect 567834 244938 567866 245174
rect 568102 244938 568186 245174
rect 568422 244938 568454 245174
rect 567834 209494 568454 244938
rect 567834 209258 567866 209494
rect 568102 209258 568186 209494
rect 568422 209258 568454 209494
rect 567834 209174 568454 209258
rect 567834 208938 567866 209174
rect 568102 208938 568186 209174
rect 568422 208938 568454 209174
rect 567834 173494 568454 208938
rect 567834 173258 567866 173494
rect 568102 173258 568186 173494
rect 568422 173258 568454 173494
rect 567834 173174 568454 173258
rect 567834 172938 567866 173174
rect 568102 172938 568186 173174
rect 568422 172938 568454 173174
rect 567834 137494 568454 172938
rect 567834 137258 567866 137494
rect 568102 137258 568186 137494
rect 568422 137258 568454 137494
rect 567834 137174 568454 137258
rect 567834 136938 567866 137174
rect 568102 136938 568186 137174
rect 568422 136938 568454 137174
rect 567834 101494 568454 136938
rect 567834 101258 567866 101494
rect 568102 101258 568186 101494
rect 568422 101258 568454 101494
rect 567834 101174 568454 101258
rect 567834 100938 567866 101174
rect 568102 100938 568186 101174
rect 568422 100938 568454 101174
rect 567834 65494 568454 100938
rect 567834 65258 567866 65494
rect 568102 65258 568186 65494
rect 568422 65258 568454 65494
rect 567834 65174 568454 65258
rect 567834 64938 567866 65174
rect 568102 64938 568186 65174
rect 568422 64938 568454 65174
rect 567834 29494 568454 64938
rect 567834 29258 567866 29494
rect 568102 29258 568186 29494
rect 568422 29258 568454 29494
rect 567834 29174 568454 29258
rect 567834 28938 567866 29174
rect 568102 28938 568186 29174
rect 568422 28938 568454 29174
rect 567834 -7066 568454 28938
rect 567834 -7302 567866 -7066
rect 568102 -7302 568186 -7066
rect 568422 -7302 568454 -7066
rect 567834 -7386 568454 -7302
rect 567834 -7622 567866 -7386
rect 568102 -7622 568186 -7386
rect 568422 -7622 568454 -7386
rect 567834 -7654 568454 -7622
rect 577794 704838 578414 711590
rect 577794 704602 577826 704838
rect 578062 704602 578146 704838
rect 578382 704602 578414 704838
rect 577794 704518 578414 704602
rect 577794 704282 577826 704518
rect 578062 704282 578146 704518
rect 578382 704282 578414 704518
rect 577794 687454 578414 704282
rect 577794 687218 577826 687454
rect 578062 687218 578146 687454
rect 578382 687218 578414 687454
rect 577794 687134 578414 687218
rect 577794 686898 577826 687134
rect 578062 686898 578146 687134
rect 578382 686898 578414 687134
rect 577794 651454 578414 686898
rect 577794 651218 577826 651454
rect 578062 651218 578146 651454
rect 578382 651218 578414 651454
rect 577794 651134 578414 651218
rect 577794 650898 577826 651134
rect 578062 650898 578146 651134
rect 578382 650898 578414 651134
rect 577794 615454 578414 650898
rect 577794 615218 577826 615454
rect 578062 615218 578146 615454
rect 578382 615218 578414 615454
rect 577794 615134 578414 615218
rect 577794 614898 577826 615134
rect 578062 614898 578146 615134
rect 578382 614898 578414 615134
rect 577794 579454 578414 614898
rect 577794 579218 577826 579454
rect 578062 579218 578146 579454
rect 578382 579218 578414 579454
rect 577794 579134 578414 579218
rect 577794 578898 577826 579134
rect 578062 578898 578146 579134
rect 578382 578898 578414 579134
rect 577794 543454 578414 578898
rect 577794 543218 577826 543454
rect 578062 543218 578146 543454
rect 578382 543218 578414 543454
rect 577794 543134 578414 543218
rect 577794 542898 577826 543134
rect 578062 542898 578146 543134
rect 578382 542898 578414 543134
rect 577794 507454 578414 542898
rect 577794 507218 577826 507454
rect 578062 507218 578146 507454
rect 578382 507218 578414 507454
rect 577794 507134 578414 507218
rect 577794 506898 577826 507134
rect 578062 506898 578146 507134
rect 578382 506898 578414 507134
rect 577794 471454 578414 506898
rect 577794 471218 577826 471454
rect 578062 471218 578146 471454
rect 578382 471218 578414 471454
rect 577794 471134 578414 471218
rect 577794 470898 577826 471134
rect 578062 470898 578146 471134
rect 578382 470898 578414 471134
rect 577794 435454 578414 470898
rect 577794 435218 577826 435454
rect 578062 435218 578146 435454
rect 578382 435218 578414 435454
rect 577794 435134 578414 435218
rect 577794 434898 577826 435134
rect 578062 434898 578146 435134
rect 578382 434898 578414 435134
rect 577794 399454 578414 434898
rect 577794 399218 577826 399454
rect 578062 399218 578146 399454
rect 578382 399218 578414 399454
rect 577794 399134 578414 399218
rect 577794 398898 577826 399134
rect 578062 398898 578146 399134
rect 578382 398898 578414 399134
rect 577794 363454 578414 398898
rect 577794 363218 577826 363454
rect 578062 363218 578146 363454
rect 578382 363218 578414 363454
rect 577794 363134 578414 363218
rect 577794 362898 577826 363134
rect 578062 362898 578146 363134
rect 578382 362898 578414 363134
rect 577794 327454 578414 362898
rect 577794 327218 577826 327454
rect 578062 327218 578146 327454
rect 578382 327218 578414 327454
rect 577794 327134 578414 327218
rect 577794 326898 577826 327134
rect 578062 326898 578146 327134
rect 578382 326898 578414 327134
rect 577794 291454 578414 326898
rect 577794 291218 577826 291454
rect 578062 291218 578146 291454
rect 578382 291218 578414 291454
rect 577794 291134 578414 291218
rect 577794 290898 577826 291134
rect 578062 290898 578146 291134
rect 578382 290898 578414 291134
rect 577794 255454 578414 290898
rect 577794 255218 577826 255454
rect 578062 255218 578146 255454
rect 578382 255218 578414 255454
rect 577794 255134 578414 255218
rect 577794 254898 577826 255134
rect 578062 254898 578146 255134
rect 578382 254898 578414 255134
rect 577794 219454 578414 254898
rect 577794 219218 577826 219454
rect 578062 219218 578146 219454
rect 578382 219218 578414 219454
rect 577794 219134 578414 219218
rect 577794 218898 577826 219134
rect 578062 218898 578146 219134
rect 578382 218898 578414 219134
rect 577794 183454 578414 218898
rect 577794 183218 577826 183454
rect 578062 183218 578146 183454
rect 578382 183218 578414 183454
rect 577794 183134 578414 183218
rect 577794 182898 577826 183134
rect 578062 182898 578146 183134
rect 578382 182898 578414 183134
rect 577794 147454 578414 182898
rect 577794 147218 577826 147454
rect 578062 147218 578146 147454
rect 578382 147218 578414 147454
rect 577794 147134 578414 147218
rect 577794 146898 577826 147134
rect 578062 146898 578146 147134
rect 578382 146898 578414 147134
rect 577794 111454 578414 146898
rect 577794 111218 577826 111454
rect 578062 111218 578146 111454
rect 578382 111218 578414 111454
rect 577794 111134 578414 111218
rect 577794 110898 577826 111134
rect 578062 110898 578146 111134
rect 578382 110898 578414 111134
rect 577794 75454 578414 110898
rect 577794 75218 577826 75454
rect 578062 75218 578146 75454
rect 578382 75218 578414 75454
rect 577794 75134 578414 75218
rect 577794 74898 577826 75134
rect 578062 74898 578146 75134
rect 578382 74898 578414 75134
rect 577794 39454 578414 74898
rect 577794 39218 577826 39454
rect 578062 39218 578146 39454
rect 578382 39218 578414 39454
rect 577794 39134 578414 39218
rect 577794 38898 577826 39134
rect 578062 38898 578146 39134
rect 578382 38898 578414 39134
rect 577794 3454 578414 38898
rect 577794 3218 577826 3454
rect 578062 3218 578146 3454
rect 578382 3218 578414 3454
rect 577794 3134 578414 3218
rect 577794 2898 577826 3134
rect 578062 2898 578146 3134
rect 578382 2898 578414 3134
rect 577794 -346 578414 2898
rect 577794 -582 577826 -346
rect 578062 -582 578146 -346
rect 578382 -582 578414 -346
rect 577794 -666 578414 -582
rect 577794 -902 577826 -666
rect 578062 -902 578146 -666
rect 578382 -902 578414 -666
rect 577794 -7654 578414 -902
rect 581514 705798 582134 711590
rect 592030 711558 592650 711590
rect 592030 711322 592062 711558
rect 592298 711322 592382 711558
rect 592618 711322 592650 711558
rect 592030 711238 592650 711322
rect 592030 711002 592062 711238
rect 592298 711002 592382 711238
rect 592618 711002 592650 711238
rect 591070 710598 591690 710630
rect 591070 710362 591102 710598
rect 591338 710362 591422 710598
rect 591658 710362 591690 710598
rect 591070 710278 591690 710362
rect 591070 710042 591102 710278
rect 591338 710042 591422 710278
rect 591658 710042 591690 710278
rect 590110 709638 590730 709670
rect 590110 709402 590142 709638
rect 590378 709402 590462 709638
rect 590698 709402 590730 709638
rect 590110 709318 590730 709402
rect 590110 709082 590142 709318
rect 590378 709082 590462 709318
rect 590698 709082 590730 709318
rect 589150 708678 589770 708710
rect 589150 708442 589182 708678
rect 589418 708442 589502 708678
rect 589738 708442 589770 708678
rect 589150 708358 589770 708442
rect 589150 708122 589182 708358
rect 589418 708122 589502 708358
rect 589738 708122 589770 708358
rect 588190 707718 588810 707750
rect 588190 707482 588222 707718
rect 588458 707482 588542 707718
rect 588778 707482 588810 707718
rect 588190 707398 588810 707482
rect 588190 707162 588222 707398
rect 588458 707162 588542 707398
rect 588778 707162 588810 707398
rect 587230 706758 587850 706790
rect 587230 706522 587262 706758
rect 587498 706522 587582 706758
rect 587818 706522 587850 706758
rect 587230 706438 587850 706522
rect 587230 706202 587262 706438
rect 587498 706202 587582 706438
rect 587818 706202 587850 706438
rect 581514 705562 581546 705798
rect 581782 705562 581866 705798
rect 582102 705562 582134 705798
rect 581514 705478 582134 705562
rect 581514 705242 581546 705478
rect 581782 705242 581866 705478
rect 582102 705242 582134 705478
rect 581514 691174 582134 705242
rect 586270 705798 586890 705830
rect 586270 705562 586302 705798
rect 586538 705562 586622 705798
rect 586858 705562 586890 705798
rect 586270 705478 586890 705562
rect 586270 705242 586302 705478
rect 586538 705242 586622 705478
rect 586858 705242 586890 705478
rect 581514 690938 581546 691174
rect 581782 690938 581866 691174
rect 582102 690938 582134 691174
rect 581514 690854 582134 690938
rect 581514 690618 581546 690854
rect 581782 690618 581866 690854
rect 582102 690618 582134 690854
rect 581514 655174 582134 690618
rect 581514 654938 581546 655174
rect 581782 654938 581866 655174
rect 582102 654938 582134 655174
rect 581514 654854 582134 654938
rect 581514 654618 581546 654854
rect 581782 654618 581866 654854
rect 582102 654618 582134 654854
rect 581514 619174 582134 654618
rect 581514 618938 581546 619174
rect 581782 618938 581866 619174
rect 582102 618938 582134 619174
rect 581514 618854 582134 618938
rect 581514 618618 581546 618854
rect 581782 618618 581866 618854
rect 582102 618618 582134 618854
rect 581514 583174 582134 618618
rect 581514 582938 581546 583174
rect 581782 582938 581866 583174
rect 582102 582938 582134 583174
rect 581514 582854 582134 582938
rect 581514 582618 581546 582854
rect 581782 582618 581866 582854
rect 582102 582618 582134 582854
rect 581514 547174 582134 582618
rect 581514 546938 581546 547174
rect 581782 546938 581866 547174
rect 582102 546938 582134 547174
rect 581514 546854 582134 546938
rect 581514 546618 581546 546854
rect 581782 546618 581866 546854
rect 582102 546618 582134 546854
rect 581514 511174 582134 546618
rect 581514 510938 581546 511174
rect 581782 510938 581866 511174
rect 582102 510938 582134 511174
rect 581514 510854 582134 510938
rect 581514 510618 581546 510854
rect 581782 510618 581866 510854
rect 582102 510618 582134 510854
rect 581514 475174 582134 510618
rect 581514 474938 581546 475174
rect 581782 474938 581866 475174
rect 582102 474938 582134 475174
rect 581514 474854 582134 474938
rect 581514 474618 581546 474854
rect 581782 474618 581866 474854
rect 582102 474618 582134 474854
rect 581514 439174 582134 474618
rect 581514 438938 581546 439174
rect 581782 438938 581866 439174
rect 582102 438938 582134 439174
rect 581514 438854 582134 438938
rect 581514 438618 581546 438854
rect 581782 438618 581866 438854
rect 582102 438618 582134 438854
rect 581514 403174 582134 438618
rect 581514 402938 581546 403174
rect 581782 402938 581866 403174
rect 582102 402938 582134 403174
rect 581514 402854 582134 402938
rect 581514 402618 581546 402854
rect 581782 402618 581866 402854
rect 582102 402618 582134 402854
rect 581514 367174 582134 402618
rect 581514 366938 581546 367174
rect 581782 366938 581866 367174
rect 582102 366938 582134 367174
rect 581514 366854 582134 366938
rect 581514 366618 581546 366854
rect 581782 366618 581866 366854
rect 582102 366618 582134 366854
rect 581514 331174 582134 366618
rect 581514 330938 581546 331174
rect 581782 330938 581866 331174
rect 582102 330938 582134 331174
rect 581514 330854 582134 330938
rect 581514 330618 581546 330854
rect 581782 330618 581866 330854
rect 582102 330618 582134 330854
rect 581514 295174 582134 330618
rect 581514 294938 581546 295174
rect 581782 294938 581866 295174
rect 582102 294938 582134 295174
rect 581514 294854 582134 294938
rect 581514 294618 581546 294854
rect 581782 294618 581866 294854
rect 582102 294618 582134 294854
rect 581514 259174 582134 294618
rect 581514 258938 581546 259174
rect 581782 258938 581866 259174
rect 582102 258938 582134 259174
rect 581514 258854 582134 258938
rect 581514 258618 581546 258854
rect 581782 258618 581866 258854
rect 582102 258618 582134 258854
rect 581514 223174 582134 258618
rect 581514 222938 581546 223174
rect 581782 222938 581866 223174
rect 582102 222938 582134 223174
rect 581514 222854 582134 222938
rect 581514 222618 581546 222854
rect 581782 222618 581866 222854
rect 582102 222618 582134 222854
rect 581514 187174 582134 222618
rect 581514 186938 581546 187174
rect 581782 186938 581866 187174
rect 582102 186938 582134 187174
rect 581514 186854 582134 186938
rect 581514 186618 581546 186854
rect 581782 186618 581866 186854
rect 582102 186618 582134 186854
rect 581514 151174 582134 186618
rect 581514 150938 581546 151174
rect 581782 150938 581866 151174
rect 582102 150938 582134 151174
rect 581514 150854 582134 150938
rect 581514 150618 581546 150854
rect 581782 150618 581866 150854
rect 582102 150618 582134 150854
rect 581514 115174 582134 150618
rect 581514 114938 581546 115174
rect 581782 114938 581866 115174
rect 582102 114938 582134 115174
rect 581514 114854 582134 114938
rect 581514 114618 581546 114854
rect 581782 114618 581866 114854
rect 582102 114618 582134 114854
rect 581514 79174 582134 114618
rect 581514 78938 581546 79174
rect 581782 78938 581866 79174
rect 582102 78938 582134 79174
rect 581514 78854 582134 78938
rect 581514 78618 581546 78854
rect 581782 78618 581866 78854
rect 582102 78618 582134 78854
rect 581514 43174 582134 78618
rect 581514 42938 581546 43174
rect 581782 42938 581866 43174
rect 582102 42938 582134 43174
rect 581514 42854 582134 42938
rect 581514 42618 581546 42854
rect 581782 42618 581866 42854
rect 582102 42618 582134 42854
rect 581514 7174 582134 42618
rect 581514 6938 581546 7174
rect 581782 6938 581866 7174
rect 582102 6938 582134 7174
rect 581514 6854 582134 6938
rect 581514 6618 581546 6854
rect 581782 6618 581866 6854
rect 582102 6618 582134 6854
rect 581514 -1306 582134 6618
rect 585310 704838 585930 704870
rect 585310 704602 585342 704838
rect 585578 704602 585662 704838
rect 585898 704602 585930 704838
rect 585310 704518 585930 704602
rect 585310 704282 585342 704518
rect 585578 704282 585662 704518
rect 585898 704282 585930 704518
rect 585310 687454 585930 704282
rect 585310 687218 585342 687454
rect 585578 687218 585662 687454
rect 585898 687218 585930 687454
rect 585310 687134 585930 687218
rect 585310 686898 585342 687134
rect 585578 686898 585662 687134
rect 585898 686898 585930 687134
rect 585310 651454 585930 686898
rect 585310 651218 585342 651454
rect 585578 651218 585662 651454
rect 585898 651218 585930 651454
rect 585310 651134 585930 651218
rect 585310 650898 585342 651134
rect 585578 650898 585662 651134
rect 585898 650898 585930 651134
rect 585310 615454 585930 650898
rect 585310 615218 585342 615454
rect 585578 615218 585662 615454
rect 585898 615218 585930 615454
rect 585310 615134 585930 615218
rect 585310 614898 585342 615134
rect 585578 614898 585662 615134
rect 585898 614898 585930 615134
rect 585310 579454 585930 614898
rect 585310 579218 585342 579454
rect 585578 579218 585662 579454
rect 585898 579218 585930 579454
rect 585310 579134 585930 579218
rect 585310 578898 585342 579134
rect 585578 578898 585662 579134
rect 585898 578898 585930 579134
rect 585310 543454 585930 578898
rect 585310 543218 585342 543454
rect 585578 543218 585662 543454
rect 585898 543218 585930 543454
rect 585310 543134 585930 543218
rect 585310 542898 585342 543134
rect 585578 542898 585662 543134
rect 585898 542898 585930 543134
rect 585310 507454 585930 542898
rect 585310 507218 585342 507454
rect 585578 507218 585662 507454
rect 585898 507218 585930 507454
rect 585310 507134 585930 507218
rect 585310 506898 585342 507134
rect 585578 506898 585662 507134
rect 585898 506898 585930 507134
rect 585310 471454 585930 506898
rect 585310 471218 585342 471454
rect 585578 471218 585662 471454
rect 585898 471218 585930 471454
rect 585310 471134 585930 471218
rect 585310 470898 585342 471134
rect 585578 470898 585662 471134
rect 585898 470898 585930 471134
rect 585310 435454 585930 470898
rect 585310 435218 585342 435454
rect 585578 435218 585662 435454
rect 585898 435218 585930 435454
rect 585310 435134 585930 435218
rect 585310 434898 585342 435134
rect 585578 434898 585662 435134
rect 585898 434898 585930 435134
rect 585310 399454 585930 434898
rect 585310 399218 585342 399454
rect 585578 399218 585662 399454
rect 585898 399218 585930 399454
rect 585310 399134 585930 399218
rect 585310 398898 585342 399134
rect 585578 398898 585662 399134
rect 585898 398898 585930 399134
rect 585310 363454 585930 398898
rect 585310 363218 585342 363454
rect 585578 363218 585662 363454
rect 585898 363218 585930 363454
rect 585310 363134 585930 363218
rect 585310 362898 585342 363134
rect 585578 362898 585662 363134
rect 585898 362898 585930 363134
rect 585310 327454 585930 362898
rect 585310 327218 585342 327454
rect 585578 327218 585662 327454
rect 585898 327218 585930 327454
rect 585310 327134 585930 327218
rect 585310 326898 585342 327134
rect 585578 326898 585662 327134
rect 585898 326898 585930 327134
rect 585310 291454 585930 326898
rect 585310 291218 585342 291454
rect 585578 291218 585662 291454
rect 585898 291218 585930 291454
rect 585310 291134 585930 291218
rect 585310 290898 585342 291134
rect 585578 290898 585662 291134
rect 585898 290898 585930 291134
rect 585310 255454 585930 290898
rect 585310 255218 585342 255454
rect 585578 255218 585662 255454
rect 585898 255218 585930 255454
rect 585310 255134 585930 255218
rect 585310 254898 585342 255134
rect 585578 254898 585662 255134
rect 585898 254898 585930 255134
rect 585310 219454 585930 254898
rect 585310 219218 585342 219454
rect 585578 219218 585662 219454
rect 585898 219218 585930 219454
rect 585310 219134 585930 219218
rect 585310 218898 585342 219134
rect 585578 218898 585662 219134
rect 585898 218898 585930 219134
rect 585310 183454 585930 218898
rect 585310 183218 585342 183454
rect 585578 183218 585662 183454
rect 585898 183218 585930 183454
rect 585310 183134 585930 183218
rect 585310 182898 585342 183134
rect 585578 182898 585662 183134
rect 585898 182898 585930 183134
rect 585310 147454 585930 182898
rect 585310 147218 585342 147454
rect 585578 147218 585662 147454
rect 585898 147218 585930 147454
rect 585310 147134 585930 147218
rect 585310 146898 585342 147134
rect 585578 146898 585662 147134
rect 585898 146898 585930 147134
rect 585310 111454 585930 146898
rect 585310 111218 585342 111454
rect 585578 111218 585662 111454
rect 585898 111218 585930 111454
rect 585310 111134 585930 111218
rect 585310 110898 585342 111134
rect 585578 110898 585662 111134
rect 585898 110898 585930 111134
rect 585310 75454 585930 110898
rect 585310 75218 585342 75454
rect 585578 75218 585662 75454
rect 585898 75218 585930 75454
rect 585310 75134 585930 75218
rect 585310 74898 585342 75134
rect 585578 74898 585662 75134
rect 585898 74898 585930 75134
rect 585310 39454 585930 74898
rect 585310 39218 585342 39454
rect 585578 39218 585662 39454
rect 585898 39218 585930 39454
rect 585310 39134 585930 39218
rect 585310 38898 585342 39134
rect 585578 38898 585662 39134
rect 585898 38898 585930 39134
rect 585310 3454 585930 38898
rect 585310 3218 585342 3454
rect 585578 3218 585662 3454
rect 585898 3218 585930 3454
rect 585310 3134 585930 3218
rect 585310 2898 585342 3134
rect 585578 2898 585662 3134
rect 585898 2898 585930 3134
rect 585310 -346 585930 2898
rect 585310 -582 585342 -346
rect 585578 -582 585662 -346
rect 585898 -582 585930 -346
rect 585310 -666 585930 -582
rect 585310 -902 585342 -666
rect 585578 -902 585662 -666
rect 585898 -902 585930 -666
rect 585310 -934 585930 -902
rect 586270 691174 586890 705242
rect 586270 690938 586302 691174
rect 586538 690938 586622 691174
rect 586858 690938 586890 691174
rect 586270 690854 586890 690938
rect 586270 690618 586302 690854
rect 586538 690618 586622 690854
rect 586858 690618 586890 690854
rect 586270 655174 586890 690618
rect 586270 654938 586302 655174
rect 586538 654938 586622 655174
rect 586858 654938 586890 655174
rect 586270 654854 586890 654938
rect 586270 654618 586302 654854
rect 586538 654618 586622 654854
rect 586858 654618 586890 654854
rect 586270 619174 586890 654618
rect 586270 618938 586302 619174
rect 586538 618938 586622 619174
rect 586858 618938 586890 619174
rect 586270 618854 586890 618938
rect 586270 618618 586302 618854
rect 586538 618618 586622 618854
rect 586858 618618 586890 618854
rect 586270 583174 586890 618618
rect 586270 582938 586302 583174
rect 586538 582938 586622 583174
rect 586858 582938 586890 583174
rect 586270 582854 586890 582938
rect 586270 582618 586302 582854
rect 586538 582618 586622 582854
rect 586858 582618 586890 582854
rect 586270 547174 586890 582618
rect 586270 546938 586302 547174
rect 586538 546938 586622 547174
rect 586858 546938 586890 547174
rect 586270 546854 586890 546938
rect 586270 546618 586302 546854
rect 586538 546618 586622 546854
rect 586858 546618 586890 546854
rect 586270 511174 586890 546618
rect 586270 510938 586302 511174
rect 586538 510938 586622 511174
rect 586858 510938 586890 511174
rect 586270 510854 586890 510938
rect 586270 510618 586302 510854
rect 586538 510618 586622 510854
rect 586858 510618 586890 510854
rect 586270 475174 586890 510618
rect 586270 474938 586302 475174
rect 586538 474938 586622 475174
rect 586858 474938 586890 475174
rect 586270 474854 586890 474938
rect 586270 474618 586302 474854
rect 586538 474618 586622 474854
rect 586858 474618 586890 474854
rect 586270 439174 586890 474618
rect 586270 438938 586302 439174
rect 586538 438938 586622 439174
rect 586858 438938 586890 439174
rect 586270 438854 586890 438938
rect 586270 438618 586302 438854
rect 586538 438618 586622 438854
rect 586858 438618 586890 438854
rect 586270 403174 586890 438618
rect 586270 402938 586302 403174
rect 586538 402938 586622 403174
rect 586858 402938 586890 403174
rect 586270 402854 586890 402938
rect 586270 402618 586302 402854
rect 586538 402618 586622 402854
rect 586858 402618 586890 402854
rect 586270 367174 586890 402618
rect 586270 366938 586302 367174
rect 586538 366938 586622 367174
rect 586858 366938 586890 367174
rect 586270 366854 586890 366938
rect 586270 366618 586302 366854
rect 586538 366618 586622 366854
rect 586858 366618 586890 366854
rect 586270 331174 586890 366618
rect 586270 330938 586302 331174
rect 586538 330938 586622 331174
rect 586858 330938 586890 331174
rect 586270 330854 586890 330938
rect 586270 330618 586302 330854
rect 586538 330618 586622 330854
rect 586858 330618 586890 330854
rect 586270 295174 586890 330618
rect 586270 294938 586302 295174
rect 586538 294938 586622 295174
rect 586858 294938 586890 295174
rect 586270 294854 586890 294938
rect 586270 294618 586302 294854
rect 586538 294618 586622 294854
rect 586858 294618 586890 294854
rect 586270 259174 586890 294618
rect 586270 258938 586302 259174
rect 586538 258938 586622 259174
rect 586858 258938 586890 259174
rect 586270 258854 586890 258938
rect 586270 258618 586302 258854
rect 586538 258618 586622 258854
rect 586858 258618 586890 258854
rect 586270 223174 586890 258618
rect 586270 222938 586302 223174
rect 586538 222938 586622 223174
rect 586858 222938 586890 223174
rect 586270 222854 586890 222938
rect 586270 222618 586302 222854
rect 586538 222618 586622 222854
rect 586858 222618 586890 222854
rect 586270 187174 586890 222618
rect 586270 186938 586302 187174
rect 586538 186938 586622 187174
rect 586858 186938 586890 187174
rect 586270 186854 586890 186938
rect 586270 186618 586302 186854
rect 586538 186618 586622 186854
rect 586858 186618 586890 186854
rect 586270 151174 586890 186618
rect 586270 150938 586302 151174
rect 586538 150938 586622 151174
rect 586858 150938 586890 151174
rect 586270 150854 586890 150938
rect 586270 150618 586302 150854
rect 586538 150618 586622 150854
rect 586858 150618 586890 150854
rect 586270 115174 586890 150618
rect 586270 114938 586302 115174
rect 586538 114938 586622 115174
rect 586858 114938 586890 115174
rect 586270 114854 586890 114938
rect 586270 114618 586302 114854
rect 586538 114618 586622 114854
rect 586858 114618 586890 114854
rect 586270 79174 586890 114618
rect 586270 78938 586302 79174
rect 586538 78938 586622 79174
rect 586858 78938 586890 79174
rect 586270 78854 586890 78938
rect 586270 78618 586302 78854
rect 586538 78618 586622 78854
rect 586858 78618 586890 78854
rect 586270 43174 586890 78618
rect 586270 42938 586302 43174
rect 586538 42938 586622 43174
rect 586858 42938 586890 43174
rect 586270 42854 586890 42938
rect 586270 42618 586302 42854
rect 586538 42618 586622 42854
rect 586858 42618 586890 42854
rect 586270 7174 586890 42618
rect 586270 6938 586302 7174
rect 586538 6938 586622 7174
rect 586858 6938 586890 7174
rect 586270 6854 586890 6938
rect 586270 6618 586302 6854
rect 586538 6618 586622 6854
rect 586858 6618 586890 6854
rect 581514 -1542 581546 -1306
rect 581782 -1542 581866 -1306
rect 582102 -1542 582134 -1306
rect 581514 -1626 582134 -1542
rect 581514 -1862 581546 -1626
rect 581782 -1862 581866 -1626
rect 582102 -1862 582134 -1626
rect 581514 -7654 582134 -1862
rect 586270 -1306 586890 6618
rect 586270 -1542 586302 -1306
rect 586538 -1542 586622 -1306
rect 586858 -1542 586890 -1306
rect 586270 -1626 586890 -1542
rect 586270 -1862 586302 -1626
rect 586538 -1862 586622 -1626
rect 586858 -1862 586890 -1626
rect 586270 -1894 586890 -1862
rect 587230 694894 587850 706202
rect 587230 694658 587262 694894
rect 587498 694658 587582 694894
rect 587818 694658 587850 694894
rect 587230 694574 587850 694658
rect 587230 694338 587262 694574
rect 587498 694338 587582 694574
rect 587818 694338 587850 694574
rect 587230 658894 587850 694338
rect 587230 658658 587262 658894
rect 587498 658658 587582 658894
rect 587818 658658 587850 658894
rect 587230 658574 587850 658658
rect 587230 658338 587262 658574
rect 587498 658338 587582 658574
rect 587818 658338 587850 658574
rect 587230 622894 587850 658338
rect 587230 622658 587262 622894
rect 587498 622658 587582 622894
rect 587818 622658 587850 622894
rect 587230 622574 587850 622658
rect 587230 622338 587262 622574
rect 587498 622338 587582 622574
rect 587818 622338 587850 622574
rect 587230 586894 587850 622338
rect 587230 586658 587262 586894
rect 587498 586658 587582 586894
rect 587818 586658 587850 586894
rect 587230 586574 587850 586658
rect 587230 586338 587262 586574
rect 587498 586338 587582 586574
rect 587818 586338 587850 586574
rect 587230 550894 587850 586338
rect 587230 550658 587262 550894
rect 587498 550658 587582 550894
rect 587818 550658 587850 550894
rect 587230 550574 587850 550658
rect 587230 550338 587262 550574
rect 587498 550338 587582 550574
rect 587818 550338 587850 550574
rect 587230 514894 587850 550338
rect 587230 514658 587262 514894
rect 587498 514658 587582 514894
rect 587818 514658 587850 514894
rect 587230 514574 587850 514658
rect 587230 514338 587262 514574
rect 587498 514338 587582 514574
rect 587818 514338 587850 514574
rect 587230 478894 587850 514338
rect 587230 478658 587262 478894
rect 587498 478658 587582 478894
rect 587818 478658 587850 478894
rect 587230 478574 587850 478658
rect 587230 478338 587262 478574
rect 587498 478338 587582 478574
rect 587818 478338 587850 478574
rect 587230 442894 587850 478338
rect 587230 442658 587262 442894
rect 587498 442658 587582 442894
rect 587818 442658 587850 442894
rect 587230 442574 587850 442658
rect 587230 442338 587262 442574
rect 587498 442338 587582 442574
rect 587818 442338 587850 442574
rect 587230 406894 587850 442338
rect 587230 406658 587262 406894
rect 587498 406658 587582 406894
rect 587818 406658 587850 406894
rect 587230 406574 587850 406658
rect 587230 406338 587262 406574
rect 587498 406338 587582 406574
rect 587818 406338 587850 406574
rect 587230 370894 587850 406338
rect 587230 370658 587262 370894
rect 587498 370658 587582 370894
rect 587818 370658 587850 370894
rect 587230 370574 587850 370658
rect 587230 370338 587262 370574
rect 587498 370338 587582 370574
rect 587818 370338 587850 370574
rect 587230 334894 587850 370338
rect 587230 334658 587262 334894
rect 587498 334658 587582 334894
rect 587818 334658 587850 334894
rect 587230 334574 587850 334658
rect 587230 334338 587262 334574
rect 587498 334338 587582 334574
rect 587818 334338 587850 334574
rect 587230 298894 587850 334338
rect 587230 298658 587262 298894
rect 587498 298658 587582 298894
rect 587818 298658 587850 298894
rect 587230 298574 587850 298658
rect 587230 298338 587262 298574
rect 587498 298338 587582 298574
rect 587818 298338 587850 298574
rect 587230 262894 587850 298338
rect 587230 262658 587262 262894
rect 587498 262658 587582 262894
rect 587818 262658 587850 262894
rect 587230 262574 587850 262658
rect 587230 262338 587262 262574
rect 587498 262338 587582 262574
rect 587818 262338 587850 262574
rect 587230 226894 587850 262338
rect 587230 226658 587262 226894
rect 587498 226658 587582 226894
rect 587818 226658 587850 226894
rect 587230 226574 587850 226658
rect 587230 226338 587262 226574
rect 587498 226338 587582 226574
rect 587818 226338 587850 226574
rect 587230 190894 587850 226338
rect 587230 190658 587262 190894
rect 587498 190658 587582 190894
rect 587818 190658 587850 190894
rect 587230 190574 587850 190658
rect 587230 190338 587262 190574
rect 587498 190338 587582 190574
rect 587818 190338 587850 190574
rect 587230 154894 587850 190338
rect 587230 154658 587262 154894
rect 587498 154658 587582 154894
rect 587818 154658 587850 154894
rect 587230 154574 587850 154658
rect 587230 154338 587262 154574
rect 587498 154338 587582 154574
rect 587818 154338 587850 154574
rect 587230 118894 587850 154338
rect 587230 118658 587262 118894
rect 587498 118658 587582 118894
rect 587818 118658 587850 118894
rect 587230 118574 587850 118658
rect 587230 118338 587262 118574
rect 587498 118338 587582 118574
rect 587818 118338 587850 118574
rect 587230 82894 587850 118338
rect 587230 82658 587262 82894
rect 587498 82658 587582 82894
rect 587818 82658 587850 82894
rect 587230 82574 587850 82658
rect 587230 82338 587262 82574
rect 587498 82338 587582 82574
rect 587818 82338 587850 82574
rect 587230 46894 587850 82338
rect 587230 46658 587262 46894
rect 587498 46658 587582 46894
rect 587818 46658 587850 46894
rect 587230 46574 587850 46658
rect 587230 46338 587262 46574
rect 587498 46338 587582 46574
rect 587818 46338 587850 46574
rect 587230 10894 587850 46338
rect 587230 10658 587262 10894
rect 587498 10658 587582 10894
rect 587818 10658 587850 10894
rect 587230 10574 587850 10658
rect 587230 10338 587262 10574
rect 587498 10338 587582 10574
rect 587818 10338 587850 10574
rect 587230 -2266 587850 10338
rect 587230 -2502 587262 -2266
rect 587498 -2502 587582 -2266
rect 587818 -2502 587850 -2266
rect 587230 -2586 587850 -2502
rect 587230 -2822 587262 -2586
rect 587498 -2822 587582 -2586
rect 587818 -2822 587850 -2586
rect 587230 -2854 587850 -2822
rect 588190 698614 588810 707162
rect 588190 698378 588222 698614
rect 588458 698378 588542 698614
rect 588778 698378 588810 698614
rect 588190 698294 588810 698378
rect 588190 698058 588222 698294
rect 588458 698058 588542 698294
rect 588778 698058 588810 698294
rect 588190 662614 588810 698058
rect 588190 662378 588222 662614
rect 588458 662378 588542 662614
rect 588778 662378 588810 662614
rect 588190 662294 588810 662378
rect 588190 662058 588222 662294
rect 588458 662058 588542 662294
rect 588778 662058 588810 662294
rect 588190 626614 588810 662058
rect 588190 626378 588222 626614
rect 588458 626378 588542 626614
rect 588778 626378 588810 626614
rect 588190 626294 588810 626378
rect 588190 626058 588222 626294
rect 588458 626058 588542 626294
rect 588778 626058 588810 626294
rect 588190 590614 588810 626058
rect 588190 590378 588222 590614
rect 588458 590378 588542 590614
rect 588778 590378 588810 590614
rect 588190 590294 588810 590378
rect 588190 590058 588222 590294
rect 588458 590058 588542 590294
rect 588778 590058 588810 590294
rect 588190 554614 588810 590058
rect 588190 554378 588222 554614
rect 588458 554378 588542 554614
rect 588778 554378 588810 554614
rect 588190 554294 588810 554378
rect 588190 554058 588222 554294
rect 588458 554058 588542 554294
rect 588778 554058 588810 554294
rect 588190 518614 588810 554058
rect 588190 518378 588222 518614
rect 588458 518378 588542 518614
rect 588778 518378 588810 518614
rect 588190 518294 588810 518378
rect 588190 518058 588222 518294
rect 588458 518058 588542 518294
rect 588778 518058 588810 518294
rect 588190 482614 588810 518058
rect 588190 482378 588222 482614
rect 588458 482378 588542 482614
rect 588778 482378 588810 482614
rect 588190 482294 588810 482378
rect 588190 482058 588222 482294
rect 588458 482058 588542 482294
rect 588778 482058 588810 482294
rect 588190 446614 588810 482058
rect 588190 446378 588222 446614
rect 588458 446378 588542 446614
rect 588778 446378 588810 446614
rect 588190 446294 588810 446378
rect 588190 446058 588222 446294
rect 588458 446058 588542 446294
rect 588778 446058 588810 446294
rect 588190 410614 588810 446058
rect 588190 410378 588222 410614
rect 588458 410378 588542 410614
rect 588778 410378 588810 410614
rect 588190 410294 588810 410378
rect 588190 410058 588222 410294
rect 588458 410058 588542 410294
rect 588778 410058 588810 410294
rect 588190 374614 588810 410058
rect 588190 374378 588222 374614
rect 588458 374378 588542 374614
rect 588778 374378 588810 374614
rect 588190 374294 588810 374378
rect 588190 374058 588222 374294
rect 588458 374058 588542 374294
rect 588778 374058 588810 374294
rect 588190 338614 588810 374058
rect 588190 338378 588222 338614
rect 588458 338378 588542 338614
rect 588778 338378 588810 338614
rect 588190 338294 588810 338378
rect 588190 338058 588222 338294
rect 588458 338058 588542 338294
rect 588778 338058 588810 338294
rect 588190 302614 588810 338058
rect 588190 302378 588222 302614
rect 588458 302378 588542 302614
rect 588778 302378 588810 302614
rect 588190 302294 588810 302378
rect 588190 302058 588222 302294
rect 588458 302058 588542 302294
rect 588778 302058 588810 302294
rect 588190 266614 588810 302058
rect 588190 266378 588222 266614
rect 588458 266378 588542 266614
rect 588778 266378 588810 266614
rect 588190 266294 588810 266378
rect 588190 266058 588222 266294
rect 588458 266058 588542 266294
rect 588778 266058 588810 266294
rect 588190 230614 588810 266058
rect 588190 230378 588222 230614
rect 588458 230378 588542 230614
rect 588778 230378 588810 230614
rect 588190 230294 588810 230378
rect 588190 230058 588222 230294
rect 588458 230058 588542 230294
rect 588778 230058 588810 230294
rect 588190 194614 588810 230058
rect 588190 194378 588222 194614
rect 588458 194378 588542 194614
rect 588778 194378 588810 194614
rect 588190 194294 588810 194378
rect 588190 194058 588222 194294
rect 588458 194058 588542 194294
rect 588778 194058 588810 194294
rect 588190 158614 588810 194058
rect 588190 158378 588222 158614
rect 588458 158378 588542 158614
rect 588778 158378 588810 158614
rect 588190 158294 588810 158378
rect 588190 158058 588222 158294
rect 588458 158058 588542 158294
rect 588778 158058 588810 158294
rect 588190 122614 588810 158058
rect 588190 122378 588222 122614
rect 588458 122378 588542 122614
rect 588778 122378 588810 122614
rect 588190 122294 588810 122378
rect 588190 122058 588222 122294
rect 588458 122058 588542 122294
rect 588778 122058 588810 122294
rect 588190 86614 588810 122058
rect 588190 86378 588222 86614
rect 588458 86378 588542 86614
rect 588778 86378 588810 86614
rect 588190 86294 588810 86378
rect 588190 86058 588222 86294
rect 588458 86058 588542 86294
rect 588778 86058 588810 86294
rect 588190 50614 588810 86058
rect 588190 50378 588222 50614
rect 588458 50378 588542 50614
rect 588778 50378 588810 50614
rect 588190 50294 588810 50378
rect 588190 50058 588222 50294
rect 588458 50058 588542 50294
rect 588778 50058 588810 50294
rect 588190 14614 588810 50058
rect 588190 14378 588222 14614
rect 588458 14378 588542 14614
rect 588778 14378 588810 14614
rect 588190 14294 588810 14378
rect 588190 14058 588222 14294
rect 588458 14058 588542 14294
rect 588778 14058 588810 14294
rect 588190 -3226 588810 14058
rect 588190 -3462 588222 -3226
rect 588458 -3462 588542 -3226
rect 588778 -3462 588810 -3226
rect 588190 -3546 588810 -3462
rect 588190 -3782 588222 -3546
rect 588458 -3782 588542 -3546
rect 588778 -3782 588810 -3546
rect 588190 -3814 588810 -3782
rect 589150 666334 589770 708122
rect 589150 666098 589182 666334
rect 589418 666098 589502 666334
rect 589738 666098 589770 666334
rect 589150 666014 589770 666098
rect 589150 665778 589182 666014
rect 589418 665778 589502 666014
rect 589738 665778 589770 666014
rect 589150 630334 589770 665778
rect 589150 630098 589182 630334
rect 589418 630098 589502 630334
rect 589738 630098 589770 630334
rect 589150 630014 589770 630098
rect 589150 629778 589182 630014
rect 589418 629778 589502 630014
rect 589738 629778 589770 630014
rect 589150 594334 589770 629778
rect 589150 594098 589182 594334
rect 589418 594098 589502 594334
rect 589738 594098 589770 594334
rect 589150 594014 589770 594098
rect 589150 593778 589182 594014
rect 589418 593778 589502 594014
rect 589738 593778 589770 594014
rect 589150 558334 589770 593778
rect 589150 558098 589182 558334
rect 589418 558098 589502 558334
rect 589738 558098 589770 558334
rect 589150 558014 589770 558098
rect 589150 557778 589182 558014
rect 589418 557778 589502 558014
rect 589738 557778 589770 558014
rect 589150 522334 589770 557778
rect 589150 522098 589182 522334
rect 589418 522098 589502 522334
rect 589738 522098 589770 522334
rect 589150 522014 589770 522098
rect 589150 521778 589182 522014
rect 589418 521778 589502 522014
rect 589738 521778 589770 522014
rect 589150 486334 589770 521778
rect 589150 486098 589182 486334
rect 589418 486098 589502 486334
rect 589738 486098 589770 486334
rect 589150 486014 589770 486098
rect 589150 485778 589182 486014
rect 589418 485778 589502 486014
rect 589738 485778 589770 486014
rect 589150 450334 589770 485778
rect 589150 450098 589182 450334
rect 589418 450098 589502 450334
rect 589738 450098 589770 450334
rect 589150 450014 589770 450098
rect 589150 449778 589182 450014
rect 589418 449778 589502 450014
rect 589738 449778 589770 450014
rect 589150 414334 589770 449778
rect 589150 414098 589182 414334
rect 589418 414098 589502 414334
rect 589738 414098 589770 414334
rect 589150 414014 589770 414098
rect 589150 413778 589182 414014
rect 589418 413778 589502 414014
rect 589738 413778 589770 414014
rect 589150 378334 589770 413778
rect 589150 378098 589182 378334
rect 589418 378098 589502 378334
rect 589738 378098 589770 378334
rect 589150 378014 589770 378098
rect 589150 377778 589182 378014
rect 589418 377778 589502 378014
rect 589738 377778 589770 378014
rect 589150 342334 589770 377778
rect 589150 342098 589182 342334
rect 589418 342098 589502 342334
rect 589738 342098 589770 342334
rect 589150 342014 589770 342098
rect 589150 341778 589182 342014
rect 589418 341778 589502 342014
rect 589738 341778 589770 342014
rect 589150 306334 589770 341778
rect 589150 306098 589182 306334
rect 589418 306098 589502 306334
rect 589738 306098 589770 306334
rect 589150 306014 589770 306098
rect 589150 305778 589182 306014
rect 589418 305778 589502 306014
rect 589738 305778 589770 306014
rect 589150 270334 589770 305778
rect 589150 270098 589182 270334
rect 589418 270098 589502 270334
rect 589738 270098 589770 270334
rect 589150 270014 589770 270098
rect 589150 269778 589182 270014
rect 589418 269778 589502 270014
rect 589738 269778 589770 270014
rect 589150 234334 589770 269778
rect 589150 234098 589182 234334
rect 589418 234098 589502 234334
rect 589738 234098 589770 234334
rect 589150 234014 589770 234098
rect 589150 233778 589182 234014
rect 589418 233778 589502 234014
rect 589738 233778 589770 234014
rect 589150 198334 589770 233778
rect 589150 198098 589182 198334
rect 589418 198098 589502 198334
rect 589738 198098 589770 198334
rect 589150 198014 589770 198098
rect 589150 197778 589182 198014
rect 589418 197778 589502 198014
rect 589738 197778 589770 198014
rect 589150 162334 589770 197778
rect 589150 162098 589182 162334
rect 589418 162098 589502 162334
rect 589738 162098 589770 162334
rect 589150 162014 589770 162098
rect 589150 161778 589182 162014
rect 589418 161778 589502 162014
rect 589738 161778 589770 162014
rect 589150 126334 589770 161778
rect 589150 126098 589182 126334
rect 589418 126098 589502 126334
rect 589738 126098 589770 126334
rect 589150 126014 589770 126098
rect 589150 125778 589182 126014
rect 589418 125778 589502 126014
rect 589738 125778 589770 126014
rect 589150 90334 589770 125778
rect 589150 90098 589182 90334
rect 589418 90098 589502 90334
rect 589738 90098 589770 90334
rect 589150 90014 589770 90098
rect 589150 89778 589182 90014
rect 589418 89778 589502 90014
rect 589738 89778 589770 90014
rect 589150 54334 589770 89778
rect 589150 54098 589182 54334
rect 589418 54098 589502 54334
rect 589738 54098 589770 54334
rect 589150 54014 589770 54098
rect 589150 53778 589182 54014
rect 589418 53778 589502 54014
rect 589738 53778 589770 54014
rect 589150 18334 589770 53778
rect 589150 18098 589182 18334
rect 589418 18098 589502 18334
rect 589738 18098 589770 18334
rect 589150 18014 589770 18098
rect 589150 17778 589182 18014
rect 589418 17778 589502 18014
rect 589738 17778 589770 18014
rect 589150 -4186 589770 17778
rect 589150 -4422 589182 -4186
rect 589418 -4422 589502 -4186
rect 589738 -4422 589770 -4186
rect 589150 -4506 589770 -4422
rect 589150 -4742 589182 -4506
rect 589418 -4742 589502 -4506
rect 589738 -4742 589770 -4506
rect 589150 -4774 589770 -4742
rect 590110 670054 590730 709082
rect 590110 669818 590142 670054
rect 590378 669818 590462 670054
rect 590698 669818 590730 670054
rect 590110 669734 590730 669818
rect 590110 669498 590142 669734
rect 590378 669498 590462 669734
rect 590698 669498 590730 669734
rect 590110 634054 590730 669498
rect 590110 633818 590142 634054
rect 590378 633818 590462 634054
rect 590698 633818 590730 634054
rect 590110 633734 590730 633818
rect 590110 633498 590142 633734
rect 590378 633498 590462 633734
rect 590698 633498 590730 633734
rect 590110 598054 590730 633498
rect 590110 597818 590142 598054
rect 590378 597818 590462 598054
rect 590698 597818 590730 598054
rect 590110 597734 590730 597818
rect 590110 597498 590142 597734
rect 590378 597498 590462 597734
rect 590698 597498 590730 597734
rect 590110 562054 590730 597498
rect 590110 561818 590142 562054
rect 590378 561818 590462 562054
rect 590698 561818 590730 562054
rect 590110 561734 590730 561818
rect 590110 561498 590142 561734
rect 590378 561498 590462 561734
rect 590698 561498 590730 561734
rect 590110 526054 590730 561498
rect 590110 525818 590142 526054
rect 590378 525818 590462 526054
rect 590698 525818 590730 526054
rect 590110 525734 590730 525818
rect 590110 525498 590142 525734
rect 590378 525498 590462 525734
rect 590698 525498 590730 525734
rect 590110 490054 590730 525498
rect 590110 489818 590142 490054
rect 590378 489818 590462 490054
rect 590698 489818 590730 490054
rect 590110 489734 590730 489818
rect 590110 489498 590142 489734
rect 590378 489498 590462 489734
rect 590698 489498 590730 489734
rect 590110 454054 590730 489498
rect 590110 453818 590142 454054
rect 590378 453818 590462 454054
rect 590698 453818 590730 454054
rect 590110 453734 590730 453818
rect 590110 453498 590142 453734
rect 590378 453498 590462 453734
rect 590698 453498 590730 453734
rect 590110 418054 590730 453498
rect 590110 417818 590142 418054
rect 590378 417818 590462 418054
rect 590698 417818 590730 418054
rect 590110 417734 590730 417818
rect 590110 417498 590142 417734
rect 590378 417498 590462 417734
rect 590698 417498 590730 417734
rect 590110 382054 590730 417498
rect 590110 381818 590142 382054
rect 590378 381818 590462 382054
rect 590698 381818 590730 382054
rect 590110 381734 590730 381818
rect 590110 381498 590142 381734
rect 590378 381498 590462 381734
rect 590698 381498 590730 381734
rect 590110 346054 590730 381498
rect 590110 345818 590142 346054
rect 590378 345818 590462 346054
rect 590698 345818 590730 346054
rect 590110 345734 590730 345818
rect 590110 345498 590142 345734
rect 590378 345498 590462 345734
rect 590698 345498 590730 345734
rect 590110 310054 590730 345498
rect 590110 309818 590142 310054
rect 590378 309818 590462 310054
rect 590698 309818 590730 310054
rect 590110 309734 590730 309818
rect 590110 309498 590142 309734
rect 590378 309498 590462 309734
rect 590698 309498 590730 309734
rect 590110 274054 590730 309498
rect 590110 273818 590142 274054
rect 590378 273818 590462 274054
rect 590698 273818 590730 274054
rect 590110 273734 590730 273818
rect 590110 273498 590142 273734
rect 590378 273498 590462 273734
rect 590698 273498 590730 273734
rect 590110 238054 590730 273498
rect 590110 237818 590142 238054
rect 590378 237818 590462 238054
rect 590698 237818 590730 238054
rect 590110 237734 590730 237818
rect 590110 237498 590142 237734
rect 590378 237498 590462 237734
rect 590698 237498 590730 237734
rect 590110 202054 590730 237498
rect 590110 201818 590142 202054
rect 590378 201818 590462 202054
rect 590698 201818 590730 202054
rect 590110 201734 590730 201818
rect 590110 201498 590142 201734
rect 590378 201498 590462 201734
rect 590698 201498 590730 201734
rect 590110 166054 590730 201498
rect 590110 165818 590142 166054
rect 590378 165818 590462 166054
rect 590698 165818 590730 166054
rect 590110 165734 590730 165818
rect 590110 165498 590142 165734
rect 590378 165498 590462 165734
rect 590698 165498 590730 165734
rect 590110 130054 590730 165498
rect 590110 129818 590142 130054
rect 590378 129818 590462 130054
rect 590698 129818 590730 130054
rect 590110 129734 590730 129818
rect 590110 129498 590142 129734
rect 590378 129498 590462 129734
rect 590698 129498 590730 129734
rect 590110 94054 590730 129498
rect 590110 93818 590142 94054
rect 590378 93818 590462 94054
rect 590698 93818 590730 94054
rect 590110 93734 590730 93818
rect 590110 93498 590142 93734
rect 590378 93498 590462 93734
rect 590698 93498 590730 93734
rect 590110 58054 590730 93498
rect 590110 57818 590142 58054
rect 590378 57818 590462 58054
rect 590698 57818 590730 58054
rect 590110 57734 590730 57818
rect 590110 57498 590142 57734
rect 590378 57498 590462 57734
rect 590698 57498 590730 57734
rect 590110 22054 590730 57498
rect 590110 21818 590142 22054
rect 590378 21818 590462 22054
rect 590698 21818 590730 22054
rect 590110 21734 590730 21818
rect 590110 21498 590142 21734
rect 590378 21498 590462 21734
rect 590698 21498 590730 21734
rect 590110 -5146 590730 21498
rect 590110 -5382 590142 -5146
rect 590378 -5382 590462 -5146
rect 590698 -5382 590730 -5146
rect 590110 -5466 590730 -5382
rect 590110 -5702 590142 -5466
rect 590378 -5702 590462 -5466
rect 590698 -5702 590730 -5466
rect 590110 -5734 590730 -5702
rect 591070 673774 591690 710042
rect 591070 673538 591102 673774
rect 591338 673538 591422 673774
rect 591658 673538 591690 673774
rect 591070 673454 591690 673538
rect 591070 673218 591102 673454
rect 591338 673218 591422 673454
rect 591658 673218 591690 673454
rect 591070 637774 591690 673218
rect 591070 637538 591102 637774
rect 591338 637538 591422 637774
rect 591658 637538 591690 637774
rect 591070 637454 591690 637538
rect 591070 637218 591102 637454
rect 591338 637218 591422 637454
rect 591658 637218 591690 637454
rect 591070 601774 591690 637218
rect 591070 601538 591102 601774
rect 591338 601538 591422 601774
rect 591658 601538 591690 601774
rect 591070 601454 591690 601538
rect 591070 601218 591102 601454
rect 591338 601218 591422 601454
rect 591658 601218 591690 601454
rect 591070 565774 591690 601218
rect 591070 565538 591102 565774
rect 591338 565538 591422 565774
rect 591658 565538 591690 565774
rect 591070 565454 591690 565538
rect 591070 565218 591102 565454
rect 591338 565218 591422 565454
rect 591658 565218 591690 565454
rect 591070 529774 591690 565218
rect 591070 529538 591102 529774
rect 591338 529538 591422 529774
rect 591658 529538 591690 529774
rect 591070 529454 591690 529538
rect 591070 529218 591102 529454
rect 591338 529218 591422 529454
rect 591658 529218 591690 529454
rect 591070 493774 591690 529218
rect 591070 493538 591102 493774
rect 591338 493538 591422 493774
rect 591658 493538 591690 493774
rect 591070 493454 591690 493538
rect 591070 493218 591102 493454
rect 591338 493218 591422 493454
rect 591658 493218 591690 493454
rect 591070 457774 591690 493218
rect 591070 457538 591102 457774
rect 591338 457538 591422 457774
rect 591658 457538 591690 457774
rect 591070 457454 591690 457538
rect 591070 457218 591102 457454
rect 591338 457218 591422 457454
rect 591658 457218 591690 457454
rect 591070 421774 591690 457218
rect 591070 421538 591102 421774
rect 591338 421538 591422 421774
rect 591658 421538 591690 421774
rect 591070 421454 591690 421538
rect 591070 421218 591102 421454
rect 591338 421218 591422 421454
rect 591658 421218 591690 421454
rect 591070 385774 591690 421218
rect 591070 385538 591102 385774
rect 591338 385538 591422 385774
rect 591658 385538 591690 385774
rect 591070 385454 591690 385538
rect 591070 385218 591102 385454
rect 591338 385218 591422 385454
rect 591658 385218 591690 385454
rect 591070 349774 591690 385218
rect 591070 349538 591102 349774
rect 591338 349538 591422 349774
rect 591658 349538 591690 349774
rect 591070 349454 591690 349538
rect 591070 349218 591102 349454
rect 591338 349218 591422 349454
rect 591658 349218 591690 349454
rect 591070 313774 591690 349218
rect 591070 313538 591102 313774
rect 591338 313538 591422 313774
rect 591658 313538 591690 313774
rect 591070 313454 591690 313538
rect 591070 313218 591102 313454
rect 591338 313218 591422 313454
rect 591658 313218 591690 313454
rect 591070 277774 591690 313218
rect 591070 277538 591102 277774
rect 591338 277538 591422 277774
rect 591658 277538 591690 277774
rect 591070 277454 591690 277538
rect 591070 277218 591102 277454
rect 591338 277218 591422 277454
rect 591658 277218 591690 277454
rect 591070 241774 591690 277218
rect 591070 241538 591102 241774
rect 591338 241538 591422 241774
rect 591658 241538 591690 241774
rect 591070 241454 591690 241538
rect 591070 241218 591102 241454
rect 591338 241218 591422 241454
rect 591658 241218 591690 241454
rect 591070 205774 591690 241218
rect 591070 205538 591102 205774
rect 591338 205538 591422 205774
rect 591658 205538 591690 205774
rect 591070 205454 591690 205538
rect 591070 205218 591102 205454
rect 591338 205218 591422 205454
rect 591658 205218 591690 205454
rect 591070 169774 591690 205218
rect 591070 169538 591102 169774
rect 591338 169538 591422 169774
rect 591658 169538 591690 169774
rect 591070 169454 591690 169538
rect 591070 169218 591102 169454
rect 591338 169218 591422 169454
rect 591658 169218 591690 169454
rect 591070 133774 591690 169218
rect 591070 133538 591102 133774
rect 591338 133538 591422 133774
rect 591658 133538 591690 133774
rect 591070 133454 591690 133538
rect 591070 133218 591102 133454
rect 591338 133218 591422 133454
rect 591658 133218 591690 133454
rect 591070 97774 591690 133218
rect 591070 97538 591102 97774
rect 591338 97538 591422 97774
rect 591658 97538 591690 97774
rect 591070 97454 591690 97538
rect 591070 97218 591102 97454
rect 591338 97218 591422 97454
rect 591658 97218 591690 97454
rect 591070 61774 591690 97218
rect 591070 61538 591102 61774
rect 591338 61538 591422 61774
rect 591658 61538 591690 61774
rect 591070 61454 591690 61538
rect 591070 61218 591102 61454
rect 591338 61218 591422 61454
rect 591658 61218 591690 61454
rect 591070 25774 591690 61218
rect 591070 25538 591102 25774
rect 591338 25538 591422 25774
rect 591658 25538 591690 25774
rect 591070 25454 591690 25538
rect 591070 25218 591102 25454
rect 591338 25218 591422 25454
rect 591658 25218 591690 25454
rect 591070 -6106 591690 25218
rect 591070 -6342 591102 -6106
rect 591338 -6342 591422 -6106
rect 591658 -6342 591690 -6106
rect 591070 -6426 591690 -6342
rect 591070 -6662 591102 -6426
rect 591338 -6662 591422 -6426
rect 591658 -6662 591690 -6426
rect 591070 -6694 591690 -6662
rect 592030 677494 592650 711002
rect 592030 677258 592062 677494
rect 592298 677258 592382 677494
rect 592618 677258 592650 677494
rect 592030 677174 592650 677258
rect 592030 676938 592062 677174
rect 592298 676938 592382 677174
rect 592618 676938 592650 677174
rect 592030 641494 592650 676938
rect 592030 641258 592062 641494
rect 592298 641258 592382 641494
rect 592618 641258 592650 641494
rect 592030 641174 592650 641258
rect 592030 640938 592062 641174
rect 592298 640938 592382 641174
rect 592618 640938 592650 641174
rect 592030 605494 592650 640938
rect 592030 605258 592062 605494
rect 592298 605258 592382 605494
rect 592618 605258 592650 605494
rect 592030 605174 592650 605258
rect 592030 604938 592062 605174
rect 592298 604938 592382 605174
rect 592618 604938 592650 605174
rect 592030 569494 592650 604938
rect 592030 569258 592062 569494
rect 592298 569258 592382 569494
rect 592618 569258 592650 569494
rect 592030 569174 592650 569258
rect 592030 568938 592062 569174
rect 592298 568938 592382 569174
rect 592618 568938 592650 569174
rect 592030 533494 592650 568938
rect 592030 533258 592062 533494
rect 592298 533258 592382 533494
rect 592618 533258 592650 533494
rect 592030 533174 592650 533258
rect 592030 532938 592062 533174
rect 592298 532938 592382 533174
rect 592618 532938 592650 533174
rect 592030 497494 592650 532938
rect 592030 497258 592062 497494
rect 592298 497258 592382 497494
rect 592618 497258 592650 497494
rect 592030 497174 592650 497258
rect 592030 496938 592062 497174
rect 592298 496938 592382 497174
rect 592618 496938 592650 497174
rect 592030 461494 592650 496938
rect 592030 461258 592062 461494
rect 592298 461258 592382 461494
rect 592618 461258 592650 461494
rect 592030 461174 592650 461258
rect 592030 460938 592062 461174
rect 592298 460938 592382 461174
rect 592618 460938 592650 461174
rect 592030 425494 592650 460938
rect 592030 425258 592062 425494
rect 592298 425258 592382 425494
rect 592618 425258 592650 425494
rect 592030 425174 592650 425258
rect 592030 424938 592062 425174
rect 592298 424938 592382 425174
rect 592618 424938 592650 425174
rect 592030 389494 592650 424938
rect 592030 389258 592062 389494
rect 592298 389258 592382 389494
rect 592618 389258 592650 389494
rect 592030 389174 592650 389258
rect 592030 388938 592062 389174
rect 592298 388938 592382 389174
rect 592618 388938 592650 389174
rect 592030 353494 592650 388938
rect 592030 353258 592062 353494
rect 592298 353258 592382 353494
rect 592618 353258 592650 353494
rect 592030 353174 592650 353258
rect 592030 352938 592062 353174
rect 592298 352938 592382 353174
rect 592618 352938 592650 353174
rect 592030 317494 592650 352938
rect 592030 317258 592062 317494
rect 592298 317258 592382 317494
rect 592618 317258 592650 317494
rect 592030 317174 592650 317258
rect 592030 316938 592062 317174
rect 592298 316938 592382 317174
rect 592618 316938 592650 317174
rect 592030 281494 592650 316938
rect 592030 281258 592062 281494
rect 592298 281258 592382 281494
rect 592618 281258 592650 281494
rect 592030 281174 592650 281258
rect 592030 280938 592062 281174
rect 592298 280938 592382 281174
rect 592618 280938 592650 281174
rect 592030 245494 592650 280938
rect 592030 245258 592062 245494
rect 592298 245258 592382 245494
rect 592618 245258 592650 245494
rect 592030 245174 592650 245258
rect 592030 244938 592062 245174
rect 592298 244938 592382 245174
rect 592618 244938 592650 245174
rect 592030 209494 592650 244938
rect 592030 209258 592062 209494
rect 592298 209258 592382 209494
rect 592618 209258 592650 209494
rect 592030 209174 592650 209258
rect 592030 208938 592062 209174
rect 592298 208938 592382 209174
rect 592618 208938 592650 209174
rect 592030 173494 592650 208938
rect 592030 173258 592062 173494
rect 592298 173258 592382 173494
rect 592618 173258 592650 173494
rect 592030 173174 592650 173258
rect 592030 172938 592062 173174
rect 592298 172938 592382 173174
rect 592618 172938 592650 173174
rect 592030 137494 592650 172938
rect 592030 137258 592062 137494
rect 592298 137258 592382 137494
rect 592618 137258 592650 137494
rect 592030 137174 592650 137258
rect 592030 136938 592062 137174
rect 592298 136938 592382 137174
rect 592618 136938 592650 137174
rect 592030 101494 592650 136938
rect 592030 101258 592062 101494
rect 592298 101258 592382 101494
rect 592618 101258 592650 101494
rect 592030 101174 592650 101258
rect 592030 100938 592062 101174
rect 592298 100938 592382 101174
rect 592618 100938 592650 101174
rect 592030 65494 592650 100938
rect 592030 65258 592062 65494
rect 592298 65258 592382 65494
rect 592618 65258 592650 65494
rect 592030 65174 592650 65258
rect 592030 64938 592062 65174
rect 592298 64938 592382 65174
rect 592618 64938 592650 65174
rect 592030 29494 592650 64938
rect 592030 29258 592062 29494
rect 592298 29258 592382 29494
rect 592618 29258 592650 29494
rect 592030 29174 592650 29258
rect 592030 28938 592062 29174
rect 592298 28938 592382 29174
rect 592618 28938 592650 29174
rect 592030 -7066 592650 28938
rect 592030 -7302 592062 -7066
rect 592298 -7302 592382 -7066
rect 592618 -7302 592650 -7066
rect 592030 -7386 592650 -7302
rect 592030 -7622 592062 -7386
rect 592298 -7622 592382 -7386
rect 592618 -7622 592650 -7386
rect 592030 -7654 592650 -7622
<< via4 >>
rect -8694 711322 -8458 711558
rect -8374 711322 -8138 711558
rect -8694 711002 -8458 711238
rect -8374 711002 -8138 711238
rect -8694 677258 -8458 677494
rect -8374 677258 -8138 677494
rect -8694 676938 -8458 677174
rect -8374 676938 -8138 677174
rect -8694 641258 -8458 641494
rect -8374 641258 -8138 641494
rect -8694 640938 -8458 641174
rect -8374 640938 -8138 641174
rect -8694 605258 -8458 605494
rect -8374 605258 -8138 605494
rect -8694 604938 -8458 605174
rect -8374 604938 -8138 605174
rect -8694 569258 -8458 569494
rect -8374 569258 -8138 569494
rect -8694 568938 -8458 569174
rect -8374 568938 -8138 569174
rect -8694 533258 -8458 533494
rect -8374 533258 -8138 533494
rect -8694 532938 -8458 533174
rect -8374 532938 -8138 533174
rect -8694 497258 -8458 497494
rect -8374 497258 -8138 497494
rect -8694 496938 -8458 497174
rect -8374 496938 -8138 497174
rect -8694 461258 -8458 461494
rect -8374 461258 -8138 461494
rect -8694 460938 -8458 461174
rect -8374 460938 -8138 461174
rect -8694 425258 -8458 425494
rect -8374 425258 -8138 425494
rect -8694 424938 -8458 425174
rect -8374 424938 -8138 425174
rect -8694 389258 -8458 389494
rect -8374 389258 -8138 389494
rect -8694 388938 -8458 389174
rect -8374 388938 -8138 389174
rect -8694 353258 -8458 353494
rect -8374 353258 -8138 353494
rect -8694 352938 -8458 353174
rect -8374 352938 -8138 353174
rect -8694 317258 -8458 317494
rect -8374 317258 -8138 317494
rect -8694 316938 -8458 317174
rect -8374 316938 -8138 317174
rect -8694 281258 -8458 281494
rect -8374 281258 -8138 281494
rect -8694 280938 -8458 281174
rect -8374 280938 -8138 281174
rect -8694 245258 -8458 245494
rect -8374 245258 -8138 245494
rect -8694 244938 -8458 245174
rect -8374 244938 -8138 245174
rect -8694 209258 -8458 209494
rect -8374 209258 -8138 209494
rect -8694 208938 -8458 209174
rect -8374 208938 -8138 209174
rect -8694 173258 -8458 173494
rect -8374 173258 -8138 173494
rect -8694 172938 -8458 173174
rect -8374 172938 -8138 173174
rect -8694 137258 -8458 137494
rect -8374 137258 -8138 137494
rect -8694 136938 -8458 137174
rect -8374 136938 -8138 137174
rect -8694 101258 -8458 101494
rect -8374 101258 -8138 101494
rect -8694 100938 -8458 101174
rect -8374 100938 -8138 101174
rect -8694 65258 -8458 65494
rect -8374 65258 -8138 65494
rect -8694 64938 -8458 65174
rect -8374 64938 -8138 65174
rect -8694 29258 -8458 29494
rect -8374 29258 -8138 29494
rect -8694 28938 -8458 29174
rect -8374 28938 -8138 29174
rect -7734 710362 -7498 710598
rect -7414 710362 -7178 710598
rect -7734 710042 -7498 710278
rect -7414 710042 -7178 710278
rect -7734 673538 -7498 673774
rect -7414 673538 -7178 673774
rect -7734 673218 -7498 673454
rect -7414 673218 -7178 673454
rect -7734 637538 -7498 637774
rect -7414 637538 -7178 637774
rect -7734 637218 -7498 637454
rect -7414 637218 -7178 637454
rect -7734 601538 -7498 601774
rect -7414 601538 -7178 601774
rect -7734 601218 -7498 601454
rect -7414 601218 -7178 601454
rect -7734 565538 -7498 565774
rect -7414 565538 -7178 565774
rect -7734 565218 -7498 565454
rect -7414 565218 -7178 565454
rect -7734 529538 -7498 529774
rect -7414 529538 -7178 529774
rect -7734 529218 -7498 529454
rect -7414 529218 -7178 529454
rect -7734 493538 -7498 493774
rect -7414 493538 -7178 493774
rect -7734 493218 -7498 493454
rect -7414 493218 -7178 493454
rect -7734 457538 -7498 457774
rect -7414 457538 -7178 457774
rect -7734 457218 -7498 457454
rect -7414 457218 -7178 457454
rect -7734 421538 -7498 421774
rect -7414 421538 -7178 421774
rect -7734 421218 -7498 421454
rect -7414 421218 -7178 421454
rect -7734 385538 -7498 385774
rect -7414 385538 -7178 385774
rect -7734 385218 -7498 385454
rect -7414 385218 -7178 385454
rect -7734 349538 -7498 349774
rect -7414 349538 -7178 349774
rect -7734 349218 -7498 349454
rect -7414 349218 -7178 349454
rect -7734 313538 -7498 313774
rect -7414 313538 -7178 313774
rect -7734 313218 -7498 313454
rect -7414 313218 -7178 313454
rect -7734 277538 -7498 277774
rect -7414 277538 -7178 277774
rect -7734 277218 -7498 277454
rect -7414 277218 -7178 277454
rect -7734 241538 -7498 241774
rect -7414 241538 -7178 241774
rect -7734 241218 -7498 241454
rect -7414 241218 -7178 241454
rect -7734 205538 -7498 205774
rect -7414 205538 -7178 205774
rect -7734 205218 -7498 205454
rect -7414 205218 -7178 205454
rect -7734 169538 -7498 169774
rect -7414 169538 -7178 169774
rect -7734 169218 -7498 169454
rect -7414 169218 -7178 169454
rect -7734 133538 -7498 133774
rect -7414 133538 -7178 133774
rect -7734 133218 -7498 133454
rect -7414 133218 -7178 133454
rect -7734 97538 -7498 97774
rect -7414 97538 -7178 97774
rect -7734 97218 -7498 97454
rect -7414 97218 -7178 97454
rect -7734 61538 -7498 61774
rect -7414 61538 -7178 61774
rect -7734 61218 -7498 61454
rect -7414 61218 -7178 61454
rect -7734 25538 -7498 25774
rect -7414 25538 -7178 25774
rect -7734 25218 -7498 25454
rect -7414 25218 -7178 25454
rect -6774 709402 -6538 709638
rect -6454 709402 -6218 709638
rect -6774 709082 -6538 709318
rect -6454 709082 -6218 709318
rect -6774 669818 -6538 670054
rect -6454 669818 -6218 670054
rect -6774 669498 -6538 669734
rect -6454 669498 -6218 669734
rect -6774 633818 -6538 634054
rect -6454 633818 -6218 634054
rect -6774 633498 -6538 633734
rect -6454 633498 -6218 633734
rect -6774 597818 -6538 598054
rect -6454 597818 -6218 598054
rect -6774 597498 -6538 597734
rect -6454 597498 -6218 597734
rect -6774 561818 -6538 562054
rect -6454 561818 -6218 562054
rect -6774 561498 -6538 561734
rect -6454 561498 -6218 561734
rect -6774 525818 -6538 526054
rect -6454 525818 -6218 526054
rect -6774 525498 -6538 525734
rect -6454 525498 -6218 525734
rect -6774 489818 -6538 490054
rect -6454 489818 -6218 490054
rect -6774 489498 -6538 489734
rect -6454 489498 -6218 489734
rect -6774 453818 -6538 454054
rect -6454 453818 -6218 454054
rect -6774 453498 -6538 453734
rect -6454 453498 -6218 453734
rect -6774 417818 -6538 418054
rect -6454 417818 -6218 418054
rect -6774 417498 -6538 417734
rect -6454 417498 -6218 417734
rect -6774 381818 -6538 382054
rect -6454 381818 -6218 382054
rect -6774 381498 -6538 381734
rect -6454 381498 -6218 381734
rect -6774 345818 -6538 346054
rect -6454 345818 -6218 346054
rect -6774 345498 -6538 345734
rect -6454 345498 -6218 345734
rect -6774 309818 -6538 310054
rect -6454 309818 -6218 310054
rect -6774 309498 -6538 309734
rect -6454 309498 -6218 309734
rect -6774 273818 -6538 274054
rect -6454 273818 -6218 274054
rect -6774 273498 -6538 273734
rect -6454 273498 -6218 273734
rect -6774 237818 -6538 238054
rect -6454 237818 -6218 238054
rect -6774 237498 -6538 237734
rect -6454 237498 -6218 237734
rect -6774 201818 -6538 202054
rect -6454 201818 -6218 202054
rect -6774 201498 -6538 201734
rect -6454 201498 -6218 201734
rect -6774 165818 -6538 166054
rect -6454 165818 -6218 166054
rect -6774 165498 -6538 165734
rect -6454 165498 -6218 165734
rect -6774 129818 -6538 130054
rect -6454 129818 -6218 130054
rect -6774 129498 -6538 129734
rect -6454 129498 -6218 129734
rect -6774 93818 -6538 94054
rect -6454 93818 -6218 94054
rect -6774 93498 -6538 93734
rect -6454 93498 -6218 93734
rect -6774 57818 -6538 58054
rect -6454 57818 -6218 58054
rect -6774 57498 -6538 57734
rect -6454 57498 -6218 57734
rect -6774 21818 -6538 22054
rect -6454 21818 -6218 22054
rect -6774 21498 -6538 21734
rect -6454 21498 -6218 21734
rect -5814 708442 -5578 708678
rect -5494 708442 -5258 708678
rect -5814 708122 -5578 708358
rect -5494 708122 -5258 708358
rect -5814 666098 -5578 666334
rect -5494 666098 -5258 666334
rect -5814 665778 -5578 666014
rect -5494 665778 -5258 666014
rect -5814 630098 -5578 630334
rect -5494 630098 -5258 630334
rect -5814 629778 -5578 630014
rect -5494 629778 -5258 630014
rect -5814 594098 -5578 594334
rect -5494 594098 -5258 594334
rect -5814 593778 -5578 594014
rect -5494 593778 -5258 594014
rect -5814 558098 -5578 558334
rect -5494 558098 -5258 558334
rect -5814 557778 -5578 558014
rect -5494 557778 -5258 558014
rect -5814 522098 -5578 522334
rect -5494 522098 -5258 522334
rect -5814 521778 -5578 522014
rect -5494 521778 -5258 522014
rect -5814 486098 -5578 486334
rect -5494 486098 -5258 486334
rect -5814 485778 -5578 486014
rect -5494 485778 -5258 486014
rect -5814 450098 -5578 450334
rect -5494 450098 -5258 450334
rect -5814 449778 -5578 450014
rect -5494 449778 -5258 450014
rect -5814 414098 -5578 414334
rect -5494 414098 -5258 414334
rect -5814 413778 -5578 414014
rect -5494 413778 -5258 414014
rect -5814 378098 -5578 378334
rect -5494 378098 -5258 378334
rect -5814 377778 -5578 378014
rect -5494 377778 -5258 378014
rect -5814 342098 -5578 342334
rect -5494 342098 -5258 342334
rect -5814 341778 -5578 342014
rect -5494 341778 -5258 342014
rect -5814 306098 -5578 306334
rect -5494 306098 -5258 306334
rect -5814 305778 -5578 306014
rect -5494 305778 -5258 306014
rect -5814 270098 -5578 270334
rect -5494 270098 -5258 270334
rect -5814 269778 -5578 270014
rect -5494 269778 -5258 270014
rect -5814 234098 -5578 234334
rect -5494 234098 -5258 234334
rect -5814 233778 -5578 234014
rect -5494 233778 -5258 234014
rect -5814 198098 -5578 198334
rect -5494 198098 -5258 198334
rect -5814 197778 -5578 198014
rect -5494 197778 -5258 198014
rect -5814 162098 -5578 162334
rect -5494 162098 -5258 162334
rect -5814 161778 -5578 162014
rect -5494 161778 -5258 162014
rect -5814 126098 -5578 126334
rect -5494 126098 -5258 126334
rect -5814 125778 -5578 126014
rect -5494 125778 -5258 126014
rect -5814 90098 -5578 90334
rect -5494 90098 -5258 90334
rect -5814 89778 -5578 90014
rect -5494 89778 -5258 90014
rect -5814 54098 -5578 54334
rect -5494 54098 -5258 54334
rect -5814 53778 -5578 54014
rect -5494 53778 -5258 54014
rect -5814 18098 -5578 18334
rect -5494 18098 -5258 18334
rect -5814 17778 -5578 18014
rect -5494 17778 -5258 18014
rect -4854 707482 -4618 707718
rect -4534 707482 -4298 707718
rect -4854 707162 -4618 707398
rect -4534 707162 -4298 707398
rect -4854 698378 -4618 698614
rect -4534 698378 -4298 698614
rect -4854 698058 -4618 698294
rect -4534 698058 -4298 698294
rect -4854 662378 -4618 662614
rect -4534 662378 -4298 662614
rect -4854 662058 -4618 662294
rect -4534 662058 -4298 662294
rect -4854 626378 -4618 626614
rect -4534 626378 -4298 626614
rect -4854 626058 -4618 626294
rect -4534 626058 -4298 626294
rect -4854 590378 -4618 590614
rect -4534 590378 -4298 590614
rect -4854 590058 -4618 590294
rect -4534 590058 -4298 590294
rect -4854 554378 -4618 554614
rect -4534 554378 -4298 554614
rect -4854 554058 -4618 554294
rect -4534 554058 -4298 554294
rect -4854 518378 -4618 518614
rect -4534 518378 -4298 518614
rect -4854 518058 -4618 518294
rect -4534 518058 -4298 518294
rect -4854 482378 -4618 482614
rect -4534 482378 -4298 482614
rect -4854 482058 -4618 482294
rect -4534 482058 -4298 482294
rect -4854 446378 -4618 446614
rect -4534 446378 -4298 446614
rect -4854 446058 -4618 446294
rect -4534 446058 -4298 446294
rect -4854 410378 -4618 410614
rect -4534 410378 -4298 410614
rect -4854 410058 -4618 410294
rect -4534 410058 -4298 410294
rect -4854 374378 -4618 374614
rect -4534 374378 -4298 374614
rect -4854 374058 -4618 374294
rect -4534 374058 -4298 374294
rect -4854 338378 -4618 338614
rect -4534 338378 -4298 338614
rect -4854 338058 -4618 338294
rect -4534 338058 -4298 338294
rect -4854 302378 -4618 302614
rect -4534 302378 -4298 302614
rect -4854 302058 -4618 302294
rect -4534 302058 -4298 302294
rect -4854 266378 -4618 266614
rect -4534 266378 -4298 266614
rect -4854 266058 -4618 266294
rect -4534 266058 -4298 266294
rect -4854 230378 -4618 230614
rect -4534 230378 -4298 230614
rect -4854 230058 -4618 230294
rect -4534 230058 -4298 230294
rect -4854 194378 -4618 194614
rect -4534 194378 -4298 194614
rect -4854 194058 -4618 194294
rect -4534 194058 -4298 194294
rect -4854 158378 -4618 158614
rect -4534 158378 -4298 158614
rect -4854 158058 -4618 158294
rect -4534 158058 -4298 158294
rect -4854 122378 -4618 122614
rect -4534 122378 -4298 122614
rect -4854 122058 -4618 122294
rect -4534 122058 -4298 122294
rect -4854 86378 -4618 86614
rect -4534 86378 -4298 86614
rect -4854 86058 -4618 86294
rect -4534 86058 -4298 86294
rect -4854 50378 -4618 50614
rect -4534 50378 -4298 50614
rect -4854 50058 -4618 50294
rect -4534 50058 -4298 50294
rect -4854 14378 -4618 14614
rect -4534 14378 -4298 14614
rect -4854 14058 -4618 14294
rect -4534 14058 -4298 14294
rect -3894 706522 -3658 706758
rect -3574 706522 -3338 706758
rect -3894 706202 -3658 706438
rect -3574 706202 -3338 706438
rect -3894 694658 -3658 694894
rect -3574 694658 -3338 694894
rect -3894 694338 -3658 694574
rect -3574 694338 -3338 694574
rect -3894 658658 -3658 658894
rect -3574 658658 -3338 658894
rect -3894 658338 -3658 658574
rect -3574 658338 -3338 658574
rect -3894 622658 -3658 622894
rect -3574 622658 -3338 622894
rect -3894 622338 -3658 622574
rect -3574 622338 -3338 622574
rect -3894 586658 -3658 586894
rect -3574 586658 -3338 586894
rect -3894 586338 -3658 586574
rect -3574 586338 -3338 586574
rect -3894 550658 -3658 550894
rect -3574 550658 -3338 550894
rect -3894 550338 -3658 550574
rect -3574 550338 -3338 550574
rect -3894 514658 -3658 514894
rect -3574 514658 -3338 514894
rect -3894 514338 -3658 514574
rect -3574 514338 -3338 514574
rect -3894 478658 -3658 478894
rect -3574 478658 -3338 478894
rect -3894 478338 -3658 478574
rect -3574 478338 -3338 478574
rect -3894 442658 -3658 442894
rect -3574 442658 -3338 442894
rect -3894 442338 -3658 442574
rect -3574 442338 -3338 442574
rect -3894 406658 -3658 406894
rect -3574 406658 -3338 406894
rect -3894 406338 -3658 406574
rect -3574 406338 -3338 406574
rect -3894 370658 -3658 370894
rect -3574 370658 -3338 370894
rect -3894 370338 -3658 370574
rect -3574 370338 -3338 370574
rect -3894 334658 -3658 334894
rect -3574 334658 -3338 334894
rect -3894 334338 -3658 334574
rect -3574 334338 -3338 334574
rect -3894 298658 -3658 298894
rect -3574 298658 -3338 298894
rect -3894 298338 -3658 298574
rect -3574 298338 -3338 298574
rect -3894 262658 -3658 262894
rect -3574 262658 -3338 262894
rect -3894 262338 -3658 262574
rect -3574 262338 -3338 262574
rect -3894 226658 -3658 226894
rect -3574 226658 -3338 226894
rect -3894 226338 -3658 226574
rect -3574 226338 -3338 226574
rect -3894 190658 -3658 190894
rect -3574 190658 -3338 190894
rect -3894 190338 -3658 190574
rect -3574 190338 -3338 190574
rect -3894 154658 -3658 154894
rect -3574 154658 -3338 154894
rect -3894 154338 -3658 154574
rect -3574 154338 -3338 154574
rect -3894 118658 -3658 118894
rect -3574 118658 -3338 118894
rect -3894 118338 -3658 118574
rect -3574 118338 -3338 118574
rect -3894 82658 -3658 82894
rect -3574 82658 -3338 82894
rect -3894 82338 -3658 82574
rect -3574 82338 -3338 82574
rect -3894 46658 -3658 46894
rect -3574 46658 -3338 46894
rect -3894 46338 -3658 46574
rect -3574 46338 -3338 46574
rect -3894 10658 -3658 10894
rect -3574 10658 -3338 10894
rect -3894 10338 -3658 10574
rect -3574 10338 -3338 10574
rect -2934 705562 -2698 705798
rect -2614 705562 -2378 705798
rect -2934 705242 -2698 705478
rect -2614 705242 -2378 705478
rect -2934 690938 -2698 691174
rect -2614 690938 -2378 691174
rect -2934 690618 -2698 690854
rect -2614 690618 -2378 690854
rect -2934 654938 -2698 655174
rect -2614 654938 -2378 655174
rect -2934 654618 -2698 654854
rect -2614 654618 -2378 654854
rect -2934 618938 -2698 619174
rect -2614 618938 -2378 619174
rect -2934 618618 -2698 618854
rect -2614 618618 -2378 618854
rect -2934 582938 -2698 583174
rect -2614 582938 -2378 583174
rect -2934 582618 -2698 582854
rect -2614 582618 -2378 582854
rect -2934 546938 -2698 547174
rect -2614 546938 -2378 547174
rect -2934 546618 -2698 546854
rect -2614 546618 -2378 546854
rect -2934 510938 -2698 511174
rect -2614 510938 -2378 511174
rect -2934 510618 -2698 510854
rect -2614 510618 -2378 510854
rect -2934 474938 -2698 475174
rect -2614 474938 -2378 475174
rect -2934 474618 -2698 474854
rect -2614 474618 -2378 474854
rect -2934 438938 -2698 439174
rect -2614 438938 -2378 439174
rect -2934 438618 -2698 438854
rect -2614 438618 -2378 438854
rect -2934 402938 -2698 403174
rect -2614 402938 -2378 403174
rect -2934 402618 -2698 402854
rect -2614 402618 -2378 402854
rect -2934 366938 -2698 367174
rect -2614 366938 -2378 367174
rect -2934 366618 -2698 366854
rect -2614 366618 -2378 366854
rect -2934 330938 -2698 331174
rect -2614 330938 -2378 331174
rect -2934 330618 -2698 330854
rect -2614 330618 -2378 330854
rect -2934 294938 -2698 295174
rect -2614 294938 -2378 295174
rect -2934 294618 -2698 294854
rect -2614 294618 -2378 294854
rect -2934 258938 -2698 259174
rect -2614 258938 -2378 259174
rect -2934 258618 -2698 258854
rect -2614 258618 -2378 258854
rect -2934 222938 -2698 223174
rect -2614 222938 -2378 223174
rect -2934 222618 -2698 222854
rect -2614 222618 -2378 222854
rect -2934 186938 -2698 187174
rect -2614 186938 -2378 187174
rect -2934 186618 -2698 186854
rect -2614 186618 -2378 186854
rect -2934 150938 -2698 151174
rect -2614 150938 -2378 151174
rect -2934 150618 -2698 150854
rect -2614 150618 -2378 150854
rect -2934 114938 -2698 115174
rect -2614 114938 -2378 115174
rect -2934 114618 -2698 114854
rect -2614 114618 -2378 114854
rect -2934 78938 -2698 79174
rect -2614 78938 -2378 79174
rect -2934 78618 -2698 78854
rect -2614 78618 -2378 78854
rect -2934 42938 -2698 43174
rect -2614 42938 -2378 43174
rect -2934 42618 -2698 42854
rect -2614 42618 -2378 42854
rect -2934 6938 -2698 7174
rect -2614 6938 -2378 7174
rect -2934 6618 -2698 6854
rect -2614 6618 -2378 6854
rect -1974 704602 -1738 704838
rect -1654 704602 -1418 704838
rect -1974 704282 -1738 704518
rect -1654 704282 -1418 704518
rect -1974 687218 -1738 687454
rect -1654 687218 -1418 687454
rect -1974 686898 -1738 687134
rect -1654 686898 -1418 687134
rect -1974 651218 -1738 651454
rect -1654 651218 -1418 651454
rect -1974 650898 -1738 651134
rect -1654 650898 -1418 651134
rect -1974 615218 -1738 615454
rect -1654 615218 -1418 615454
rect -1974 614898 -1738 615134
rect -1654 614898 -1418 615134
rect -1974 579218 -1738 579454
rect -1654 579218 -1418 579454
rect -1974 578898 -1738 579134
rect -1654 578898 -1418 579134
rect -1974 543218 -1738 543454
rect -1654 543218 -1418 543454
rect -1974 542898 -1738 543134
rect -1654 542898 -1418 543134
rect -1974 507218 -1738 507454
rect -1654 507218 -1418 507454
rect -1974 506898 -1738 507134
rect -1654 506898 -1418 507134
rect -1974 471218 -1738 471454
rect -1654 471218 -1418 471454
rect -1974 470898 -1738 471134
rect -1654 470898 -1418 471134
rect -1974 435218 -1738 435454
rect -1654 435218 -1418 435454
rect -1974 434898 -1738 435134
rect -1654 434898 -1418 435134
rect -1974 399218 -1738 399454
rect -1654 399218 -1418 399454
rect -1974 398898 -1738 399134
rect -1654 398898 -1418 399134
rect -1974 363218 -1738 363454
rect -1654 363218 -1418 363454
rect -1974 362898 -1738 363134
rect -1654 362898 -1418 363134
rect -1974 327218 -1738 327454
rect -1654 327218 -1418 327454
rect -1974 326898 -1738 327134
rect -1654 326898 -1418 327134
rect -1974 291218 -1738 291454
rect -1654 291218 -1418 291454
rect -1974 290898 -1738 291134
rect -1654 290898 -1418 291134
rect -1974 255218 -1738 255454
rect -1654 255218 -1418 255454
rect -1974 254898 -1738 255134
rect -1654 254898 -1418 255134
rect -1974 219218 -1738 219454
rect -1654 219218 -1418 219454
rect -1974 218898 -1738 219134
rect -1654 218898 -1418 219134
rect -1974 183218 -1738 183454
rect -1654 183218 -1418 183454
rect -1974 182898 -1738 183134
rect -1654 182898 -1418 183134
rect -1974 147218 -1738 147454
rect -1654 147218 -1418 147454
rect -1974 146898 -1738 147134
rect -1654 146898 -1418 147134
rect -1974 111218 -1738 111454
rect -1654 111218 -1418 111454
rect -1974 110898 -1738 111134
rect -1654 110898 -1418 111134
rect -1974 75218 -1738 75454
rect -1654 75218 -1418 75454
rect -1974 74898 -1738 75134
rect -1654 74898 -1418 75134
rect -1974 39218 -1738 39454
rect -1654 39218 -1418 39454
rect -1974 38898 -1738 39134
rect -1654 38898 -1418 39134
rect -1974 3218 -1738 3454
rect -1654 3218 -1418 3454
rect -1974 2898 -1738 3134
rect -1654 2898 -1418 3134
rect -1974 -582 -1738 -346
rect -1654 -582 -1418 -346
rect -1974 -902 -1738 -666
rect -1654 -902 -1418 -666
rect 1826 704602 2062 704838
rect 2146 704602 2382 704838
rect 1826 704282 2062 704518
rect 2146 704282 2382 704518
rect 1826 687218 2062 687454
rect 2146 687218 2382 687454
rect 1826 686898 2062 687134
rect 2146 686898 2382 687134
rect 1826 651218 2062 651454
rect 2146 651218 2382 651454
rect 1826 650898 2062 651134
rect 2146 650898 2382 651134
rect 1826 615218 2062 615454
rect 2146 615218 2382 615454
rect 1826 614898 2062 615134
rect 2146 614898 2382 615134
rect 1826 579218 2062 579454
rect 2146 579218 2382 579454
rect 1826 578898 2062 579134
rect 2146 578898 2382 579134
rect 1826 543218 2062 543454
rect 2146 543218 2382 543454
rect 1826 542898 2062 543134
rect 2146 542898 2382 543134
rect 1826 507218 2062 507454
rect 2146 507218 2382 507454
rect 1826 506898 2062 507134
rect 2146 506898 2382 507134
rect 1826 471218 2062 471454
rect 2146 471218 2382 471454
rect 1826 470898 2062 471134
rect 2146 470898 2382 471134
rect 1826 435218 2062 435454
rect 2146 435218 2382 435454
rect 1826 434898 2062 435134
rect 2146 434898 2382 435134
rect 1826 399218 2062 399454
rect 2146 399218 2382 399454
rect 1826 398898 2062 399134
rect 2146 398898 2382 399134
rect 1826 363218 2062 363454
rect 2146 363218 2382 363454
rect 1826 362898 2062 363134
rect 2146 362898 2382 363134
rect 1826 327218 2062 327454
rect 2146 327218 2382 327454
rect 1826 326898 2062 327134
rect 2146 326898 2382 327134
rect 1826 291218 2062 291454
rect 2146 291218 2382 291454
rect 1826 290898 2062 291134
rect 2146 290898 2382 291134
rect 1826 255218 2062 255454
rect 2146 255218 2382 255454
rect 1826 254898 2062 255134
rect 2146 254898 2382 255134
rect 1826 219218 2062 219454
rect 2146 219218 2382 219454
rect 1826 218898 2062 219134
rect 2146 218898 2382 219134
rect 1826 183218 2062 183454
rect 2146 183218 2382 183454
rect 1826 182898 2062 183134
rect 2146 182898 2382 183134
rect 1826 147218 2062 147454
rect 2146 147218 2382 147454
rect 1826 146898 2062 147134
rect 2146 146898 2382 147134
rect 1826 111218 2062 111454
rect 2146 111218 2382 111454
rect 1826 110898 2062 111134
rect 2146 110898 2382 111134
rect 1826 75218 2062 75454
rect 2146 75218 2382 75454
rect 1826 74898 2062 75134
rect 2146 74898 2382 75134
rect 1826 39218 2062 39454
rect 2146 39218 2382 39454
rect 1826 38898 2062 39134
rect 2146 38898 2382 39134
rect 1826 3218 2062 3454
rect 2146 3218 2382 3454
rect 1826 2898 2062 3134
rect 2146 2898 2382 3134
rect 1826 -582 2062 -346
rect 2146 -582 2382 -346
rect 1826 -902 2062 -666
rect 2146 -902 2382 -666
rect -2934 -1542 -2698 -1306
rect -2614 -1542 -2378 -1306
rect -2934 -1862 -2698 -1626
rect -2614 -1862 -2378 -1626
rect -3894 -2502 -3658 -2266
rect -3574 -2502 -3338 -2266
rect -3894 -2822 -3658 -2586
rect -3574 -2822 -3338 -2586
rect -4854 -3462 -4618 -3226
rect -4534 -3462 -4298 -3226
rect -4854 -3782 -4618 -3546
rect -4534 -3782 -4298 -3546
rect -5814 -4422 -5578 -4186
rect -5494 -4422 -5258 -4186
rect -5814 -4742 -5578 -4506
rect -5494 -4742 -5258 -4506
rect -6774 -5382 -6538 -5146
rect -6454 -5382 -6218 -5146
rect -6774 -5702 -6538 -5466
rect -6454 -5702 -6218 -5466
rect -7734 -6342 -7498 -6106
rect -7414 -6342 -7178 -6106
rect -7734 -6662 -7498 -6426
rect -7414 -6662 -7178 -6426
rect -8694 -7302 -8458 -7066
rect -8374 -7302 -8138 -7066
rect -8694 -7622 -8458 -7386
rect -8374 -7622 -8138 -7386
rect 5546 705562 5782 705798
rect 5866 705562 6102 705798
rect 5546 705242 5782 705478
rect 5866 705242 6102 705478
rect 5546 690938 5782 691174
rect 5866 690938 6102 691174
rect 5546 690618 5782 690854
rect 5866 690618 6102 690854
rect 5546 654938 5782 655174
rect 5866 654938 6102 655174
rect 5546 654618 5782 654854
rect 5866 654618 6102 654854
rect 5546 618938 5782 619174
rect 5866 618938 6102 619174
rect 5546 618618 5782 618854
rect 5866 618618 6102 618854
rect 5546 582938 5782 583174
rect 5866 582938 6102 583174
rect 5546 582618 5782 582854
rect 5866 582618 6102 582854
rect 5546 546938 5782 547174
rect 5866 546938 6102 547174
rect 5546 546618 5782 546854
rect 5866 546618 6102 546854
rect 5546 510938 5782 511174
rect 5866 510938 6102 511174
rect 5546 510618 5782 510854
rect 5866 510618 6102 510854
rect 5546 474938 5782 475174
rect 5866 474938 6102 475174
rect 5546 474618 5782 474854
rect 5866 474618 6102 474854
rect 5546 438938 5782 439174
rect 5866 438938 6102 439174
rect 5546 438618 5782 438854
rect 5866 438618 6102 438854
rect 5546 402938 5782 403174
rect 5866 402938 6102 403174
rect 5546 402618 5782 402854
rect 5866 402618 6102 402854
rect 5546 366938 5782 367174
rect 5866 366938 6102 367174
rect 5546 366618 5782 366854
rect 5866 366618 6102 366854
rect 5546 330938 5782 331174
rect 5866 330938 6102 331174
rect 5546 330618 5782 330854
rect 5866 330618 6102 330854
rect 5546 294938 5782 295174
rect 5866 294938 6102 295174
rect 5546 294618 5782 294854
rect 5866 294618 6102 294854
rect 5546 258938 5782 259174
rect 5866 258938 6102 259174
rect 5546 258618 5782 258854
rect 5866 258618 6102 258854
rect 5546 222938 5782 223174
rect 5866 222938 6102 223174
rect 5546 222618 5782 222854
rect 5866 222618 6102 222854
rect 5546 186938 5782 187174
rect 5866 186938 6102 187174
rect 5546 186618 5782 186854
rect 5866 186618 6102 186854
rect 5546 150938 5782 151174
rect 5866 150938 6102 151174
rect 5546 150618 5782 150854
rect 5866 150618 6102 150854
rect 5546 114938 5782 115174
rect 5866 114938 6102 115174
rect 5546 114618 5782 114854
rect 5866 114618 6102 114854
rect 5546 78938 5782 79174
rect 5866 78938 6102 79174
rect 5546 78618 5782 78854
rect 5866 78618 6102 78854
rect 5546 42938 5782 43174
rect 5866 42938 6102 43174
rect 5546 42618 5782 42854
rect 5866 42618 6102 42854
rect 5546 6938 5782 7174
rect 5866 6938 6102 7174
rect 5546 6618 5782 6854
rect 5866 6618 6102 6854
rect 5546 -1542 5782 -1306
rect 5866 -1542 6102 -1306
rect 5546 -1862 5782 -1626
rect 5866 -1862 6102 -1626
rect 9266 706522 9502 706758
rect 9586 706522 9822 706758
rect 9266 706202 9502 706438
rect 9586 706202 9822 706438
rect 9266 694658 9502 694894
rect 9586 694658 9822 694894
rect 9266 694338 9502 694574
rect 9586 694338 9822 694574
rect 9266 658658 9502 658894
rect 9586 658658 9822 658894
rect 9266 658338 9502 658574
rect 9586 658338 9822 658574
rect 9266 622658 9502 622894
rect 9586 622658 9822 622894
rect 9266 622338 9502 622574
rect 9586 622338 9822 622574
rect 9266 586658 9502 586894
rect 9586 586658 9822 586894
rect 9266 586338 9502 586574
rect 9586 586338 9822 586574
rect 9266 550658 9502 550894
rect 9586 550658 9822 550894
rect 9266 550338 9502 550574
rect 9586 550338 9822 550574
rect 9266 514658 9502 514894
rect 9586 514658 9822 514894
rect 9266 514338 9502 514574
rect 9586 514338 9822 514574
rect 9266 478658 9502 478894
rect 9586 478658 9822 478894
rect 9266 478338 9502 478574
rect 9586 478338 9822 478574
rect 9266 442658 9502 442894
rect 9586 442658 9822 442894
rect 9266 442338 9502 442574
rect 9586 442338 9822 442574
rect 9266 406658 9502 406894
rect 9586 406658 9822 406894
rect 9266 406338 9502 406574
rect 9586 406338 9822 406574
rect 9266 370658 9502 370894
rect 9586 370658 9822 370894
rect 9266 370338 9502 370574
rect 9586 370338 9822 370574
rect 9266 334658 9502 334894
rect 9586 334658 9822 334894
rect 9266 334338 9502 334574
rect 9586 334338 9822 334574
rect 9266 298658 9502 298894
rect 9586 298658 9822 298894
rect 9266 298338 9502 298574
rect 9586 298338 9822 298574
rect 9266 262658 9502 262894
rect 9586 262658 9822 262894
rect 9266 262338 9502 262574
rect 9586 262338 9822 262574
rect 9266 226658 9502 226894
rect 9586 226658 9822 226894
rect 9266 226338 9502 226574
rect 9586 226338 9822 226574
rect 9266 190658 9502 190894
rect 9586 190658 9822 190894
rect 9266 190338 9502 190574
rect 9586 190338 9822 190574
rect 9266 154658 9502 154894
rect 9586 154658 9822 154894
rect 9266 154338 9502 154574
rect 9586 154338 9822 154574
rect 9266 118658 9502 118894
rect 9586 118658 9822 118894
rect 9266 118338 9502 118574
rect 9586 118338 9822 118574
rect 9266 82658 9502 82894
rect 9586 82658 9822 82894
rect 9266 82338 9502 82574
rect 9586 82338 9822 82574
rect 9266 46658 9502 46894
rect 9586 46658 9822 46894
rect 9266 46338 9502 46574
rect 9586 46338 9822 46574
rect 9266 10658 9502 10894
rect 9586 10658 9822 10894
rect 9266 10338 9502 10574
rect 9586 10338 9822 10574
rect 9266 -2502 9502 -2266
rect 9586 -2502 9822 -2266
rect 9266 -2822 9502 -2586
rect 9586 -2822 9822 -2586
rect 12986 707482 13222 707718
rect 13306 707482 13542 707718
rect 12986 707162 13222 707398
rect 13306 707162 13542 707398
rect 12986 698378 13222 698614
rect 13306 698378 13542 698614
rect 12986 698058 13222 698294
rect 13306 698058 13542 698294
rect 12986 662378 13222 662614
rect 13306 662378 13542 662614
rect 12986 662058 13222 662294
rect 13306 662058 13542 662294
rect 12986 626378 13222 626614
rect 13306 626378 13542 626614
rect 12986 626058 13222 626294
rect 13306 626058 13542 626294
rect 12986 590378 13222 590614
rect 13306 590378 13542 590614
rect 12986 590058 13222 590294
rect 13306 590058 13542 590294
rect 12986 554378 13222 554614
rect 13306 554378 13542 554614
rect 12986 554058 13222 554294
rect 13306 554058 13542 554294
rect 12986 518378 13222 518614
rect 13306 518378 13542 518614
rect 12986 518058 13222 518294
rect 13306 518058 13542 518294
rect 12986 482378 13222 482614
rect 13306 482378 13542 482614
rect 12986 482058 13222 482294
rect 13306 482058 13542 482294
rect 12986 446378 13222 446614
rect 13306 446378 13542 446614
rect 12986 446058 13222 446294
rect 13306 446058 13542 446294
rect 12986 410378 13222 410614
rect 13306 410378 13542 410614
rect 12986 410058 13222 410294
rect 13306 410058 13542 410294
rect 12986 374378 13222 374614
rect 13306 374378 13542 374614
rect 12986 374058 13222 374294
rect 13306 374058 13542 374294
rect 12986 338378 13222 338614
rect 13306 338378 13542 338614
rect 12986 338058 13222 338294
rect 13306 338058 13542 338294
rect 12986 302378 13222 302614
rect 13306 302378 13542 302614
rect 12986 302058 13222 302294
rect 13306 302058 13542 302294
rect 12986 266378 13222 266614
rect 13306 266378 13542 266614
rect 12986 266058 13222 266294
rect 13306 266058 13542 266294
rect 12986 230378 13222 230614
rect 13306 230378 13542 230614
rect 12986 230058 13222 230294
rect 13306 230058 13542 230294
rect 12986 194378 13222 194614
rect 13306 194378 13542 194614
rect 12986 194058 13222 194294
rect 13306 194058 13542 194294
rect 12986 158378 13222 158614
rect 13306 158378 13542 158614
rect 12986 158058 13222 158294
rect 13306 158058 13542 158294
rect 12986 122378 13222 122614
rect 13306 122378 13542 122614
rect 12986 122058 13222 122294
rect 13306 122058 13542 122294
rect 12986 86378 13222 86614
rect 13306 86378 13542 86614
rect 12986 86058 13222 86294
rect 13306 86058 13542 86294
rect 12986 50378 13222 50614
rect 13306 50378 13542 50614
rect 12986 50058 13222 50294
rect 13306 50058 13542 50294
rect 12986 14378 13222 14614
rect 13306 14378 13542 14614
rect 12986 14058 13222 14294
rect 13306 14058 13542 14294
rect 12986 -3462 13222 -3226
rect 13306 -3462 13542 -3226
rect 12986 -3782 13222 -3546
rect 13306 -3782 13542 -3546
rect 16706 708442 16942 708678
rect 17026 708442 17262 708678
rect 16706 708122 16942 708358
rect 17026 708122 17262 708358
rect 16706 666098 16942 666334
rect 17026 666098 17262 666334
rect 16706 665778 16942 666014
rect 17026 665778 17262 666014
rect 16706 630098 16942 630334
rect 17026 630098 17262 630334
rect 16706 629778 16942 630014
rect 17026 629778 17262 630014
rect 16706 594098 16942 594334
rect 17026 594098 17262 594334
rect 16706 593778 16942 594014
rect 17026 593778 17262 594014
rect 16706 558098 16942 558334
rect 17026 558098 17262 558334
rect 16706 557778 16942 558014
rect 17026 557778 17262 558014
rect 16706 522098 16942 522334
rect 17026 522098 17262 522334
rect 16706 521778 16942 522014
rect 17026 521778 17262 522014
rect 16706 486098 16942 486334
rect 17026 486098 17262 486334
rect 16706 485778 16942 486014
rect 17026 485778 17262 486014
rect 16706 450098 16942 450334
rect 17026 450098 17262 450334
rect 16706 449778 16942 450014
rect 17026 449778 17262 450014
rect 16706 414098 16942 414334
rect 17026 414098 17262 414334
rect 16706 413778 16942 414014
rect 17026 413778 17262 414014
rect 16706 378098 16942 378334
rect 17026 378098 17262 378334
rect 16706 377778 16942 378014
rect 17026 377778 17262 378014
rect 16706 342098 16942 342334
rect 17026 342098 17262 342334
rect 16706 341778 16942 342014
rect 17026 341778 17262 342014
rect 16706 306098 16942 306334
rect 17026 306098 17262 306334
rect 16706 305778 16942 306014
rect 17026 305778 17262 306014
rect 16706 270098 16942 270334
rect 17026 270098 17262 270334
rect 16706 269778 16942 270014
rect 17026 269778 17262 270014
rect 16706 234098 16942 234334
rect 17026 234098 17262 234334
rect 16706 233778 16942 234014
rect 17026 233778 17262 234014
rect 16706 198098 16942 198334
rect 17026 198098 17262 198334
rect 16706 197778 16942 198014
rect 17026 197778 17262 198014
rect 16706 162098 16942 162334
rect 17026 162098 17262 162334
rect 16706 161778 16942 162014
rect 17026 161778 17262 162014
rect 16706 126098 16942 126334
rect 17026 126098 17262 126334
rect 16706 125778 16942 126014
rect 17026 125778 17262 126014
rect 16706 90098 16942 90334
rect 17026 90098 17262 90334
rect 16706 89778 16942 90014
rect 17026 89778 17262 90014
rect 16706 54098 16942 54334
rect 17026 54098 17262 54334
rect 16706 53778 16942 54014
rect 17026 53778 17262 54014
rect 16706 18098 16942 18334
rect 17026 18098 17262 18334
rect 16706 17778 16942 18014
rect 17026 17778 17262 18014
rect 16706 -4422 16942 -4186
rect 17026 -4422 17262 -4186
rect 16706 -4742 16942 -4506
rect 17026 -4742 17262 -4506
rect 20426 709402 20662 709638
rect 20746 709402 20982 709638
rect 20426 709082 20662 709318
rect 20746 709082 20982 709318
rect 20426 669818 20662 670054
rect 20746 669818 20982 670054
rect 20426 669498 20662 669734
rect 20746 669498 20982 669734
rect 20426 633818 20662 634054
rect 20746 633818 20982 634054
rect 20426 633498 20662 633734
rect 20746 633498 20982 633734
rect 20426 597818 20662 598054
rect 20746 597818 20982 598054
rect 20426 597498 20662 597734
rect 20746 597498 20982 597734
rect 20426 561818 20662 562054
rect 20746 561818 20982 562054
rect 20426 561498 20662 561734
rect 20746 561498 20982 561734
rect 20426 525818 20662 526054
rect 20746 525818 20982 526054
rect 20426 525498 20662 525734
rect 20746 525498 20982 525734
rect 20426 489818 20662 490054
rect 20746 489818 20982 490054
rect 20426 489498 20662 489734
rect 20746 489498 20982 489734
rect 20426 453818 20662 454054
rect 20746 453818 20982 454054
rect 20426 453498 20662 453734
rect 20746 453498 20982 453734
rect 20426 417818 20662 418054
rect 20746 417818 20982 418054
rect 20426 417498 20662 417734
rect 20746 417498 20982 417734
rect 20426 381818 20662 382054
rect 20746 381818 20982 382054
rect 20426 381498 20662 381734
rect 20746 381498 20982 381734
rect 20426 345818 20662 346054
rect 20746 345818 20982 346054
rect 20426 345498 20662 345734
rect 20746 345498 20982 345734
rect 20426 309818 20662 310054
rect 20746 309818 20982 310054
rect 20426 309498 20662 309734
rect 20746 309498 20982 309734
rect 20426 273818 20662 274054
rect 20746 273818 20982 274054
rect 20426 273498 20662 273734
rect 20746 273498 20982 273734
rect 20426 237818 20662 238054
rect 20746 237818 20982 238054
rect 20426 237498 20662 237734
rect 20746 237498 20982 237734
rect 20426 201818 20662 202054
rect 20746 201818 20982 202054
rect 20426 201498 20662 201734
rect 20746 201498 20982 201734
rect 20426 165818 20662 166054
rect 20746 165818 20982 166054
rect 20426 165498 20662 165734
rect 20746 165498 20982 165734
rect 20426 129818 20662 130054
rect 20746 129818 20982 130054
rect 20426 129498 20662 129734
rect 20746 129498 20982 129734
rect 20426 93818 20662 94054
rect 20746 93818 20982 94054
rect 20426 93498 20662 93734
rect 20746 93498 20982 93734
rect 20426 57818 20662 58054
rect 20746 57818 20982 58054
rect 20426 57498 20662 57734
rect 20746 57498 20982 57734
rect 20426 21818 20662 22054
rect 20746 21818 20982 22054
rect 20426 21498 20662 21734
rect 20746 21498 20982 21734
rect 20426 -5382 20662 -5146
rect 20746 -5382 20982 -5146
rect 20426 -5702 20662 -5466
rect 20746 -5702 20982 -5466
rect 24146 710362 24382 710598
rect 24466 710362 24702 710598
rect 24146 710042 24382 710278
rect 24466 710042 24702 710278
rect 24146 673538 24382 673774
rect 24466 673538 24702 673774
rect 24146 673218 24382 673454
rect 24466 673218 24702 673454
rect 24146 637538 24382 637774
rect 24466 637538 24702 637774
rect 24146 637218 24382 637454
rect 24466 637218 24702 637454
rect 24146 601538 24382 601774
rect 24466 601538 24702 601774
rect 24146 601218 24382 601454
rect 24466 601218 24702 601454
rect 24146 565538 24382 565774
rect 24466 565538 24702 565774
rect 24146 565218 24382 565454
rect 24466 565218 24702 565454
rect 24146 529538 24382 529774
rect 24466 529538 24702 529774
rect 24146 529218 24382 529454
rect 24466 529218 24702 529454
rect 24146 493538 24382 493774
rect 24466 493538 24702 493774
rect 24146 493218 24382 493454
rect 24466 493218 24702 493454
rect 24146 457538 24382 457774
rect 24466 457538 24702 457774
rect 24146 457218 24382 457454
rect 24466 457218 24702 457454
rect 24146 421538 24382 421774
rect 24466 421538 24702 421774
rect 24146 421218 24382 421454
rect 24466 421218 24702 421454
rect 24146 385538 24382 385774
rect 24466 385538 24702 385774
rect 24146 385218 24382 385454
rect 24466 385218 24702 385454
rect 24146 349538 24382 349774
rect 24466 349538 24702 349774
rect 24146 349218 24382 349454
rect 24466 349218 24702 349454
rect 24146 313538 24382 313774
rect 24466 313538 24702 313774
rect 24146 313218 24382 313454
rect 24466 313218 24702 313454
rect 24146 277538 24382 277774
rect 24466 277538 24702 277774
rect 24146 277218 24382 277454
rect 24466 277218 24702 277454
rect 24146 241538 24382 241774
rect 24466 241538 24702 241774
rect 24146 241218 24382 241454
rect 24466 241218 24702 241454
rect 24146 205538 24382 205774
rect 24466 205538 24702 205774
rect 24146 205218 24382 205454
rect 24466 205218 24702 205454
rect 24146 169538 24382 169774
rect 24466 169538 24702 169774
rect 24146 169218 24382 169454
rect 24466 169218 24702 169454
rect 27866 711322 28102 711558
rect 28186 711322 28422 711558
rect 27866 711002 28102 711238
rect 28186 711002 28422 711238
rect 27866 677258 28102 677494
rect 28186 677258 28422 677494
rect 27866 676938 28102 677174
rect 28186 676938 28422 677174
rect 27866 641258 28102 641494
rect 28186 641258 28422 641494
rect 27866 640938 28102 641174
rect 28186 640938 28422 641174
rect 27866 605258 28102 605494
rect 28186 605258 28422 605494
rect 27866 604938 28102 605174
rect 28186 604938 28422 605174
rect 37826 704602 38062 704838
rect 38146 704602 38382 704838
rect 37826 704282 38062 704518
rect 38146 704282 38382 704518
rect 37826 687218 38062 687454
rect 38146 687218 38382 687454
rect 37826 686898 38062 687134
rect 38146 686898 38382 687134
rect 37826 651218 38062 651454
rect 38146 651218 38382 651454
rect 37826 650898 38062 651134
rect 38146 650898 38382 651134
rect 37826 615218 38062 615454
rect 38146 615218 38382 615454
rect 37826 614898 38062 615134
rect 38146 614898 38382 615134
rect 34250 579218 34486 579454
rect 34250 578898 34486 579134
rect 37826 579218 38062 579454
rect 38146 579218 38382 579454
rect 37826 578898 38062 579134
rect 38146 578898 38382 579134
rect 27866 569258 28102 569494
rect 28186 569258 28422 569494
rect 27866 568938 28102 569174
rect 28186 568938 28422 569174
rect 34250 543218 34486 543454
rect 34250 542898 34486 543134
rect 37826 543218 38062 543454
rect 38146 543218 38382 543454
rect 37826 542898 38062 543134
rect 38146 542898 38382 543134
rect 27866 533258 28102 533494
rect 28186 533258 28422 533494
rect 27866 532938 28102 533174
rect 28186 532938 28422 533174
rect 34250 507218 34486 507454
rect 34250 506898 34486 507134
rect 37826 507218 38062 507454
rect 38146 507218 38382 507454
rect 37826 506898 38062 507134
rect 38146 506898 38382 507134
rect 27866 497258 28102 497494
rect 28186 497258 28422 497494
rect 27866 496938 28102 497174
rect 28186 496938 28422 497174
rect 34250 471218 34486 471454
rect 34250 470898 34486 471134
rect 37826 471218 38062 471454
rect 38146 471218 38382 471454
rect 37826 470898 38062 471134
rect 38146 470898 38382 471134
rect 27866 461258 28102 461494
rect 28186 461258 28422 461494
rect 27866 460938 28102 461174
rect 28186 460938 28422 461174
rect 27866 425258 28102 425494
rect 28186 425258 28422 425494
rect 27866 424938 28102 425174
rect 28186 424938 28422 425174
rect 27866 389258 28102 389494
rect 28186 389258 28422 389494
rect 27866 388938 28102 389174
rect 28186 388938 28422 389174
rect 27866 353258 28102 353494
rect 28186 353258 28422 353494
rect 27866 352938 28102 353174
rect 28186 352938 28422 353174
rect 27866 317258 28102 317494
rect 28186 317258 28422 317494
rect 27866 316938 28102 317174
rect 28186 316938 28422 317174
rect 37826 435218 38062 435454
rect 38146 435218 38382 435454
rect 37826 434898 38062 435134
rect 38146 434898 38382 435134
rect 37826 399218 38062 399454
rect 38146 399218 38382 399454
rect 37826 398898 38062 399134
rect 38146 398898 38382 399134
rect 37826 363218 38062 363454
rect 38146 363218 38382 363454
rect 37826 362898 38062 363134
rect 38146 362898 38382 363134
rect 37826 327218 38062 327454
rect 38146 327218 38382 327454
rect 37826 326898 38062 327134
rect 38146 326898 38382 327134
rect 34250 291218 34486 291454
rect 34250 290898 34486 291134
rect 37826 291218 38062 291454
rect 38146 291218 38382 291454
rect 37826 290898 38062 291134
rect 38146 290898 38382 291134
rect 27866 281258 28102 281494
rect 28186 281258 28422 281494
rect 27866 280938 28102 281174
rect 28186 280938 28422 281174
rect 34250 255218 34486 255454
rect 34250 254898 34486 255134
rect 37826 255218 38062 255454
rect 38146 255218 38382 255454
rect 37826 254898 38062 255134
rect 38146 254898 38382 255134
rect 27866 245258 28102 245494
rect 28186 245258 28422 245494
rect 27866 244938 28102 245174
rect 28186 244938 28422 245174
rect 34250 219218 34486 219454
rect 34250 218898 34486 219134
rect 37826 219218 38062 219454
rect 38146 219218 38382 219454
rect 37826 218898 38062 219134
rect 38146 218898 38382 219134
rect 27866 209258 28102 209494
rect 28186 209258 28422 209494
rect 27866 208938 28102 209174
rect 28186 208938 28422 209174
rect 34250 183218 34486 183454
rect 34250 182898 34486 183134
rect 37826 183218 38062 183454
rect 38146 183218 38382 183454
rect 37826 182898 38062 183134
rect 38146 182898 38382 183134
rect 27866 173258 28102 173494
rect 28186 173258 28422 173494
rect 27866 172938 28102 173174
rect 28186 172938 28422 173174
rect 27866 137258 28102 137494
rect 28186 137258 28422 137494
rect 27866 136938 28102 137174
rect 28186 136938 28422 137174
rect 37826 147218 38062 147454
rect 38146 147218 38382 147454
rect 37826 146898 38062 147134
rect 38146 146898 38382 147134
rect 24146 133538 24382 133774
rect 24466 133538 24702 133774
rect 24146 133218 24382 133454
rect 24466 133218 24702 133454
rect 41546 705562 41782 705798
rect 41866 705562 42102 705798
rect 41546 705242 41782 705478
rect 41866 705242 42102 705478
rect 41546 690938 41782 691174
rect 41866 690938 42102 691174
rect 41546 690618 41782 690854
rect 41866 690618 42102 690854
rect 41546 654938 41782 655174
rect 41866 654938 42102 655174
rect 41546 654618 41782 654854
rect 41866 654618 42102 654854
rect 41546 618938 41782 619174
rect 41866 618938 42102 619174
rect 41546 618618 41782 618854
rect 41866 618618 42102 618854
rect 41546 582938 41782 583174
rect 41866 582938 42102 583174
rect 41546 582618 41782 582854
rect 41866 582618 42102 582854
rect 41546 546938 41782 547174
rect 41866 546938 42102 547174
rect 41546 546618 41782 546854
rect 41866 546618 42102 546854
rect 41546 510938 41782 511174
rect 41866 510938 42102 511174
rect 41546 510618 41782 510854
rect 41866 510618 42102 510854
rect 41546 474938 41782 475174
rect 41866 474938 42102 475174
rect 41546 474618 41782 474854
rect 41866 474618 42102 474854
rect 41546 438938 41782 439174
rect 41866 438938 42102 439174
rect 41546 438618 41782 438854
rect 41866 438618 42102 438854
rect 41546 402938 41782 403174
rect 41866 402938 42102 403174
rect 41546 402618 41782 402854
rect 41866 402618 42102 402854
rect 41546 366938 41782 367174
rect 41866 366938 42102 367174
rect 41546 366618 41782 366854
rect 41866 366618 42102 366854
rect 41546 330938 41782 331174
rect 41866 330938 42102 331174
rect 41546 330618 41782 330854
rect 41866 330618 42102 330854
rect 41546 294938 41782 295174
rect 41866 294938 42102 295174
rect 41546 294618 41782 294854
rect 41866 294618 42102 294854
rect 41546 258938 41782 259174
rect 41866 258938 42102 259174
rect 41546 258618 41782 258854
rect 41866 258618 42102 258854
rect 41546 222938 41782 223174
rect 41866 222938 42102 223174
rect 41546 222618 41782 222854
rect 41866 222618 42102 222854
rect 41546 186938 41782 187174
rect 41866 186938 42102 187174
rect 41546 186618 41782 186854
rect 41866 186618 42102 186854
rect 41546 150938 41782 151174
rect 41866 150938 42102 151174
rect 41546 150618 41782 150854
rect 41866 150618 42102 150854
rect 45266 706522 45502 706758
rect 45586 706522 45822 706758
rect 45266 706202 45502 706438
rect 45586 706202 45822 706438
rect 45266 694658 45502 694894
rect 45586 694658 45822 694894
rect 45266 694338 45502 694574
rect 45586 694338 45822 694574
rect 45266 658658 45502 658894
rect 45586 658658 45822 658894
rect 45266 658338 45502 658574
rect 45586 658338 45822 658574
rect 45266 622658 45502 622894
rect 45586 622658 45822 622894
rect 45266 622338 45502 622574
rect 45586 622338 45822 622574
rect 48986 707482 49222 707718
rect 49306 707482 49542 707718
rect 48986 707162 49222 707398
rect 49306 707162 49542 707398
rect 48986 698378 49222 698614
rect 49306 698378 49542 698614
rect 48986 698058 49222 698294
rect 49306 698058 49542 698294
rect 48986 662378 49222 662614
rect 49306 662378 49542 662614
rect 48986 662058 49222 662294
rect 49306 662058 49542 662294
rect 48986 626378 49222 626614
rect 49306 626378 49542 626614
rect 48986 626058 49222 626294
rect 49306 626058 49542 626294
rect 52706 708442 52942 708678
rect 53026 708442 53262 708678
rect 52706 708122 52942 708358
rect 53026 708122 53262 708358
rect 52706 666098 52942 666334
rect 53026 666098 53262 666334
rect 52706 665778 52942 666014
rect 53026 665778 53262 666014
rect 52706 630098 52942 630334
rect 53026 630098 53262 630334
rect 52706 629778 52942 630014
rect 53026 629778 53262 630014
rect 45266 586658 45502 586894
rect 45586 586658 45822 586894
rect 45266 586338 45502 586574
rect 45586 586338 45822 586574
rect 52706 594098 52942 594334
rect 53026 594098 53262 594334
rect 52706 593778 52942 594014
rect 53026 593778 53262 594014
rect 49610 582938 49846 583174
rect 49610 582618 49846 582854
rect 45266 550658 45502 550894
rect 45586 550658 45822 550894
rect 45266 550338 45502 550574
rect 45586 550338 45822 550574
rect 52706 558098 52942 558334
rect 53026 558098 53262 558334
rect 52706 557778 52942 558014
rect 53026 557778 53262 558014
rect 49610 546938 49846 547174
rect 49610 546618 49846 546854
rect 45266 514658 45502 514894
rect 45586 514658 45822 514894
rect 45266 514338 45502 514574
rect 45586 514338 45822 514574
rect 52706 522098 52942 522334
rect 53026 522098 53262 522334
rect 52706 521778 52942 522014
rect 53026 521778 53262 522014
rect 49610 510938 49846 511174
rect 49610 510618 49846 510854
rect 45266 478658 45502 478894
rect 45586 478658 45822 478894
rect 45266 478338 45502 478574
rect 45586 478338 45822 478574
rect 52706 486098 52942 486334
rect 53026 486098 53262 486334
rect 52706 485778 52942 486014
rect 53026 485778 53262 486014
rect 49610 474938 49846 475174
rect 49610 474618 49846 474854
rect 45266 442658 45502 442894
rect 45586 442658 45822 442894
rect 45266 442338 45502 442574
rect 45586 442338 45822 442574
rect 52706 450098 52942 450334
rect 53026 450098 53262 450334
rect 52706 449778 52942 450014
rect 53026 449778 53262 450014
rect 45266 406658 45502 406894
rect 45586 406658 45822 406894
rect 45266 406338 45502 406574
rect 45586 406338 45822 406574
rect 45266 370658 45502 370894
rect 45586 370658 45822 370894
rect 45266 370338 45502 370574
rect 45586 370338 45822 370574
rect 45266 334658 45502 334894
rect 45586 334658 45822 334894
rect 45266 334338 45502 334574
rect 45586 334338 45822 334574
rect 48986 410378 49222 410614
rect 49306 410378 49542 410614
rect 48986 410058 49222 410294
rect 49306 410058 49542 410294
rect 48986 374378 49222 374614
rect 49306 374378 49542 374614
rect 48986 374058 49222 374294
rect 49306 374058 49542 374294
rect 48986 338378 49222 338614
rect 49306 338378 49542 338614
rect 48986 338058 49222 338294
rect 49306 338058 49542 338294
rect 52706 414098 52942 414334
rect 53026 414098 53262 414334
rect 52706 413778 52942 414014
rect 53026 413778 53262 414014
rect 52706 378098 52942 378334
rect 53026 378098 53262 378334
rect 52706 377778 52942 378014
rect 53026 377778 53262 378014
rect 52706 342098 52942 342334
rect 53026 342098 53262 342334
rect 52706 341778 52942 342014
rect 53026 341778 53262 342014
rect 45266 298658 45502 298894
rect 45586 298658 45822 298894
rect 45266 298338 45502 298574
rect 45586 298338 45822 298574
rect 52706 306098 52942 306334
rect 53026 306098 53262 306334
rect 52706 305778 52942 306014
rect 53026 305778 53262 306014
rect 49610 294938 49846 295174
rect 49610 294618 49846 294854
rect 45266 262658 45502 262894
rect 45586 262658 45822 262894
rect 45266 262338 45502 262574
rect 45586 262338 45822 262574
rect 52706 270098 52942 270334
rect 53026 270098 53262 270334
rect 52706 269778 52942 270014
rect 53026 269778 53262 270014
rect 49610 258938 49846 259174
rect 49610 258618 49846 258854
rect 45266 226658 45502 226894
rect 45586 226658 45822 226894
rect 45266 226338 45502 226574
rect 45586 226338 45822 226574
rect 52706 234098 52942 234334
rect 53026 234098 53262 234334
rect 52706 233778 52942 234014
rect 53026 233778 53262 234014
rect 49610 222938 49846 223174
rect 49610 222618 49846 222854
rect 45266 190658 45502 190894
rect 45586 190658 45822 190894
rect 45266 190338 45502 190574
rect 45586 190338 45822 190574
rect 52706 198098 52942 198334
rect 53026 198098 53262 198334
rect 52706 197778 52942 198014
rect 53026 197778 53262 198014
rect 49610 186938 49846 187174
rect 49610 186618 49846 186854
rect 45266 154658 45502 154894
rect 45586 154658 45822 154894
rect 45266 154338 45502 154574
rect 45586 154338 45822 154574
rect 52706 162098 52942 162334
rect 53026 162098 53262 162334
rect 52706 161778 52942 162014
rect 53026 161778 53262 162014
rect 56426 709402 56662 709638
rect 56746 709402 56982 709638
rect 56426 709082 56662 709318
rect 56746 709082 56982 709318
rect 56426 669818 56662 670054
rect 56746 669818 56982 670054
rect 56426 669498 56662 669734
rect 56746 669498 56982 669734
rect 56426 633818 56662 634054
rect 56746 633818 56982 634054
rect 56426 633498 56662 633734
rect 56746 633498 56982 633734
rect 56426 597818 56662 598054
rect 56746 597818 56982 598054
rect 56426 597498 56662 597734
rect 56746 597498 56982 597734
rect 56426 561818 56662 562054
rect 56746 561818 56982 562054
rect 56426 561498 56662 561734
rect 56746 561498 56982 561734
rect 56426 525818 56662 526054
rect 56746 525818 56982 526054
rect 56426 525498 56662 525734
rect 56746 525498 56982 525734
rect 56426 489818 56662 490054
rect 56746 489818 56982 490054
rect 56426 489498 56662 489734
rect 56746 489498 56982 489734
rect 56426 453818 56662 454054
rect 56746 453818 56982 454054
rect 56426 453498 56662 453734
rect 56746 453498 56982 453734
rect 56426 417818 56662 418054
rect 56746 417818 56982 418054
rect 56426 417498 56662 417734
rect 56746 417498 56982 417734
rect 56426 381818 56662 382054
rect 56746 381818 56982 382054
rect 56426 381498 56662 381734
rect 56746 381498 56982 381734
rect 56426 345818 56662 346054
rect 56746 345818 56982 346054
rect 56426 345498 56662 345734
rect 56746 345498 56982 345734
rect 56426 309818 56662 310054
rect 56746 309818 56982 310054
rect 56426 309498 56662 309734
rect 56746 309498 56982 309734
rect 56426 273818 56662 274054
rect 56746 273818 56982 274054
rect 56426 273498 56662 273734
rect 56746 273498 56982 273734
rect 56426 237818 56662 238054
rect 56746 237818 56982 238054
rect 56426 237498 56662 237734
rect 56746 237498 56982 237734
rect 56426 201818 56662 202054
rect 56746 201818 56982 202054
rect 56426 201498 56662 201734
rect 56746 201498 56982 201734
rect 56426 165818 56662 166054
rect 56746 165818 56982 166054
rect 56426 165498 56662 165734
rect 56746 165498 56982 165734
rect 60146 710362 60382 710598
rect 60466 710362 60702 710598
rect 60146 710042 60382 710278
rect 60466 710042 60702 710278
rect 60146 673538 60382 673774
rect 60466 673538 60702 673774
rect 60146 673218 60382 673454
rect 60466 673218 60702 673454
rect 60146 637538 60382 637774
rect 60466 637538 60702 637774
rect 60146 637218 60382 637454
rect 60466 637218 60702 637454
rect 60146 601538 60382 601774
rect 60466 601538 60702 601774
rect 60146 601218 60382 601454
rect 60466 601218 60702 601454
rect 63866 711322 64102 711558
rect 64186 711322 64422 711558
rect 63866 711002 64102 711238
rect 64186 711002 64422 711238
rect 63866 677258 64102 677494
rect 64186 677258 64422 677494
rect 63866 676938 64102 677174
rect 64186 676938 64422 677174
rect 63866 641258 64102 641494
rect 64186 641258 64422 641494
rect 63866 640938 64102 641174
rect 64186 640938 64422 641174
rect 63866 605258 64102 605494
rect 64186 605258 64422 605494
rect 63866 604938 64102 605174
rect 64186 604938 64422 605174
rect 73826 704602 74062 704838
rect 74146 704602 74382 704838
rect 73826 704282 74062 704518
rect 74146 704282 74382 704518
rect 73826 687218 74062 687454
rect 74146 687218 74382 687454
rect 73826 686898 74062 687134
rect 74146 686898 74382 687134
rect 73826 651218 74062 651454
rect 74146 651218 74382 651454
rect 73826 650898 74062 651134
rect 74146 650898 74382 651134
rect 73826 615218 74062 615454
rect 74146 615218 74382 615454
rect 73826 614898 74062 615134
rect 74146 614898 74382 615134
rect 77546 705562 77782 705798
rect 77866 705562 78102 705798
rect 77546 705242 77782 705478
rect 77866 705242 78102 705478
rect 77546 690938 77782 691174
rect 77866 690938 78102 691174
rect 77546 690618 77782 690854
rect 77866 690618 78102 690854
rect 77546 654938 77782 655174
rect 77866 654938 78102 655174
rect 77546 654618 77782 654854
rect 77866 654618 78102 654854
rect 77546 618938 77782 619174
rect 77866 618938 78102 619174
rect 77546 618618 77782 618854
rect 77866 618618 78102 618854
rect 81266 706522 81502 706758
rect 81586 706522 81822 706758
rect 81266 706202 81502 706438
rect 81586 706202 81822 706438
rect 81266 694658 81502 694894
rect 81586 694658 81822 694894
rect 81266 694338 81502 694574
rect 81586 694338 81822 694574
rect 81266 658658 81502 658894
rect 81586 658658 81822 658894
rect 81266 658338 81502 658574
rect 81586 658338 81822 658574
rect 81266 622658 81502 622894
rect 81586 622658 81822 622894
rect 81266 622338 81502 622574
rect 81586 622338 81822 622574
rect 84986 707482 85222 707718
rect 85306 707482 85542 707718
rect 84986 707162 85222 707398
rect 85306 707162 85542 707398
rect 84986 698378 85222 698614
rect 85306 698378 85542 698614
rect 84986 698058 85222 698294
rect 85306 698058 85542 698294
rect 84986 662378 85222 662614
rect 85306 662378 85542 662614
rect 84986 662058 85222 662294
rect 85306 662058 85542 662294
rect 84986 626378 85222 626614
rect 85306 626378 85542 626614
rect 84986 626058 85222 626294
rect 85306 626058 85542 626294
rect 88706 708442 88942 708678
rect 89026 708442 89262 708678
rect 88706 708122 88942 708358
rect 89026 708122 89262 708358
rect 88706 666098 88942 666334
rect 89026 666098 89262 666334
rect 88706 665778 88942 666014
rect 89026 665778 89262 666014
rect 88706 630098 88942 630334
rect 89026 630098 89262 630334
rect 88706 629778 88942 630014
rect 89026 629778 89262 630014
rect 92426 709402 92662 709638
rect 92746 709402 92982 709638
rect 92426 709082 92662 709318
rect 92746 709082 92982 709318
rect 92426 669818 92662 670054
rect 92746 669818 92982 670054
rect 92426 669498 92662 669734
rect 92746 669498 92982 669734
rect 92426 633818 92662 634054
rect 92746 633818 92982 634054
rect 92426 633498 92662 633734
rect 92746 633498 92982 633734
rect 92426 597818 92662 598054
rect 92746 597818 92982 598054
rect 92426 597498 92662 597734
rect 92746 597498 92982 597734
rect 96146 710362 96382 710598
rect 96466 710362 96702 710598
rect 96146 710042 96382 710278
rect 96466 710042 96702 710278
rect 96146 673538 96382 673774
rect 96466 673538 96702 673774
rect 96146 673218 96382 673454
rect 96466 673218 96702 673454
rect 96146 637538 96382 637774
rect 96466 637538 96702 637774
rect 96146 637218 96382 637454
rect 96466 637218 96702 637454
rect 96146 601538 96382 601774
rect 96466 601538 96702 601774
rect 96146 601218 96382 601454
rect 96466 601218 96702 601454
rect 99866 711322 100102 711558
rect 100186 711322 100422 711558
rect 99866 711002 100102 711238
rect 100186 711002 100422 711238
rect 99866 677258 100102 677494
rect 100186 677258 100422 677494
rect 99866 676938 100102 677174
rect 100186 676938 100422 677174
rect 99866 641258 100102 641494
rect 100186 641258 100422 641494
rect 99866 640938 100102 641174
rect 100186 640938 100422 641174
rect 99866 605258 100102 605494
rect 100186 605258 100422 605494
rect 99866 604938 100102 605174
rect 100186 604938 100422 605174
rect 109826 704602 110062 704838
rect 110146 704602 110382 704838
rect 109826 704282 110062 704518
rect 110146 704282 110382 704518
rect 109826 687218 110062 687454
rect 110146 687218 110382 687454
rect 109826 686898 110062 687134
rect 110146 686898 110382 687134
rect 109826 651218 110062 651454
rect 110146 651218 110382 651454
rect 109826 650898 110062 651134
rect 110146 650898 110382 651134
rect 109826 615218 110062 615454
rect 110146 615218 110382 615454
rect 109826 614898 110062 615134
rect 110146 614898 110382 615134
rect 80330 582938 80566 583174
rect 80330 582618 80566 582854
rect 64970 579218 65206 579454
rect 64970 578898 65206 579134
rect 95690 579218 95926 579454
rect 95690 578898 95926 579134
rect 109826 579218 110062 579454
rect 110146 579218 110382 579454
rect 109826 578898 110062 579134
rect 110146 578898 110382 579134
rect 60146 565538 60382 565774
rect 60466 565538 60702 565774
rect 60146 565218 60382 565454
rect 60466 565218 60702 565454
rect 80330 546938 80566 547174
rect 80330 546618 80566 546854
rect 64970 543218 65206 543454
rect 64970 542898 65206 543134
rect 95690 543218 95926 543454
rect 95690 542898 95926 543134
rect 109826 543218 110062 543454
rect 110146 543218 110382 543454
rect 109826 542898 110062 543134
rect 110146 542898 110382 543134
rect 60146 529538 60382 529774
rect 60466 529538 60702 529774
rect 60146 529218 60382 529454
rect 60466 529218 60702 529454
rect 80330 510938 80566 511174
rect 80330 510618 80566 510854
rect 64970 507218 65206 507454
rect 64970 506898 65206 507134
rect 95690 507218 95926 507454
rect 95690 506898 95926 507134
rect 109826 507218 110062 507454
rect 110146 507218 110382 507454
rect 109826 506898 110062 507134
rect 110146 506898 110382 507134
rect 60146 493538 60382 493774
rect 60466 493538 60702 493774
rect 60146 493218 60382 493454
rect 60466 493218 60702 493454
rect 80330 474938 80566 475174
rect 80330 474618 80566 474854
rect 64970 471218 65206 471454
rect 64970 470898 65206 471134
rect 95690 471218 95926 471454
rect 95690 470898 95926 471134
rect 109826 471218 110062 471454
rect 110146 471218 110382 471454
rect 109826 470898 110062 471134
rect 110146 470898 110382 471134
rect 60146 457538 60382 457774
rect 60466 457538 60702 457774
rect 60146 457218 60382 457454
rect 60466 457218 60702 457454
rect 60146 421538 60382 421774
rect 60466 421538 60702 421774
rect 60146 421218 60382 421454
rect 60466 421218 60702 421454
rect 60146 385538 60382 385774
rect 60466 385538 60702 385774
rect 60146 385218 60382 385454
rect 60466 385218 60702 385454
rect 60146 349538 60382 349774
rect 60466 349538 60702 349774
rect 60146 349218 60382 349454
rect 60466 349218 60702 349454
rect 63866 425258 64102 425494
rect 64186 425258 64422 425494
rect 63866 424938 64102 425174
rect 64186 424938 64422 425174
rect 63866 389258 64102 389494
rect 64186 389258 64422 389494
rect 63866 388938 64102 389174
rect 64186 388938 64422 389174
rect 63866 353258 64102 353494
rect 64186 353258 64422 353494
rect 63866 352938 64102 353174
rect 64186 352938 64422 353174
rect 73826 435218 74062 435454
rect 74146 435218 74382 435454
rect 73826 434898 74062 435134
rect 74146 434898 74382 435134
rect 73826 399218 74062 399454
rect 74146 399218 74382 399454
rect 73826 398898 74062 399134
rect 74146 398898 74382 399134
rect 73826 363218 74062 363454
rect 74146 363218 74382 363454
rect 73826 362898 74062 363134
rect 74146 362898 74382 363134
rect 73826 327218 74062 327454
rect 74146 327218 74382 327454
rect 73826 326898 74062 327134
rect 74146 326898 74382 327134
rect 77546 438938 77782 439174
rect 77866 438938 78102 439174
rect 77546 438618 77782 438854
rect 77866 438618 78102 438854
rect 77546 402938 77782 403174
rect 77866 402938 78102 403174
rect 77546 402618 77782 402854
rect 77866 402618 78102 402854
rect 77546 366938 77782 367174
rect 77866 366938 78102 367174
rect 77546 366618 77782 366854
rect 77866 366618 78102 366854
rect 77546 330938 77782 331174
rect 77866 330938 78102 331174
rect 77546 330618 77782 330854
rect 77866 330618 78102 330854
rect 81266 442658 81502 442894
rect 81586 442658 81822 442894
rect 81266 442338 81502 442574
rect 81586 442338 81822 442574
rect 81266 406658 81502 406894
rect 81586 406658 81822 406894
rect 81266 406338 81502 406574
rect 81586 406338 81822 406574
rect 81266 370658 81502 370894
rect 81586 370658 81822 370894
rect 81266 370338 81502 370574
rect 81586 370338 81822 370574
rect 81266 334658 81502 334894
rect 81586 334658 81822 334894
rect 81266 334338 81502 334574
rect 81586 334338 81822 334574
rect 84986 446378 85222 446614
rect 85306 446378 85542 446614
rect 84986 446058 85222 446294
rect 85306 446058 85542 446294
rect 84986 410378 85222 410614
rect 85306 410378 85542 410614
rect 84986 410058 85222 410294
rect 85306 410058 85542 410294
rect 84986 374378 85222 374614
rect 85306 374378 85542 374614
rect 84986 374058 85222 374294
rect 85306 374058 85542 374294
rect 84986 338378 85222 338614
rect 85306 338378 85542 338614
rect 84986 338058 85222 338294
rect 85306 338058 85542 338294
rect 88706 414098 88942 414334
rect 89026 414098 89262 414334
rect 88706 413778 88942 414014
rect 89026 413778 89262 414014
rect 88706 378098 88942 378334
rect 89026 378098 89262 378334
rect 88706 377778 88942 378014
rect 89026 377778 89262 378014
rect 88706 342098 88942 342334
rect 89026 342098 89262 342334
rect 88706 341778 88942 342014
rect 89026 341778 89262 342014
rect 92426 417818 92662 418054
rect 92746 417818 92982 418054
rect 92426 417498 92662 417734
rect 92746 417498 92982 417734
rect 92426 381818 92662 382054
rect 92746 381818 92982 382054
rect 92426 381498 92662 381734
rect 92746 381498 92982 381734
rect 92426 345818 92662 346054
rect 92746 345818 92982 346054
rect 92426 345498 92662 345734
rect 92746 345498 92982 345734
rect 96146 421538 96382 421774
rect 96466 421538 96702 421774
rect 96146 421218 96382 421454
rect 96466 421218 96702 421454
rect 96146 385538 96382 385774
rect 96466 385538 96702 385774
rect 96146 385218 96382 385454
rect 96466 385218 96702 385454
rect 96146 349538 96382 349774
rect 96466 349538 96702 349774
rect 96146 349218 96382 349454
rect 96466 349218 96702 349454
rect 99866 425258 100102 425494
rect 100186 425258 100422 425494
rect 99866 424938 100102 425174
rect 100186 424938 100422 425174
rect 99866 389258 100102 389494
rect 100186 389258 100422 389494
rect 99866 388938 100102 389174
rect 100186 388938 100422 389174
rect 99866 353258 100102 353494
rect 100186 353258 100422 353494
rect 99866 352938 100102 353174
rect 100186 352938 100422 353174
rect 109826 435218 110062 435454
rect 110146 435218 110382 435454
rect 109826 434898 110062 435134
rect 110146 434898 110382 435134
rect 109826 399218 110062 399454
rect 110146 399218 110382 399454
rect 109826 398898 110062 399134
rect 110146 398898 110382 399134
rect 109826 363218 110062 363454
rect 110146 363218 110382 363454
rect 109826 362898 110062 363134
rect 110146 362898 110382 363134
rect 109826 327218 110062 327454
rect 110146 327218 110382 327454
rect 109826 326898 110062 327134
rect 110146 326898 110382 327134
rect 60146 313538 60382 313774
rect 60466 313538 60702 313774
rect 60146 313218 60382 313454
rect 60466 313218 60702 313454
rect 80330 294938 80566 295174
rect 80330 294618 80566 294854
rect 64970 291218 65206 291454
rect 64970 290898 65206 291134
rect 95690 291218 95926 291454
rect 95690 290898 95926 291134
rect 109826 291218 110062 291454
rect 110146 291218 110382 291454
rect 109826 290898 110062 291134
rect 110146 290898 110382 291134
rect 60146 277538 60382 277774
rect 60466 277538 60702 277774
rect 60146 277218 60382 277454
rect 60466 277218 60702 277454
rect 80330 258938 80566 259174
rect 80330 258618 80566 258854
rect 64970 255218 65206 255454
rect 64970 254898 65206 255134
rect 95690 255218 95926 255454
rect 95690 254898 95926 255134
rect 109826 255218 110062 255454
rect 110146 255218 110382 255454
rect 109826 254898 110062 255134
rect 110146 254898 110382 255134
rect 60146 241538 60382 241774
rect 60466 241538 60702 241774
rect 60146 241218 60382 241454
rect 60466 241218 60702 241454
rect 80330 222938 80566 223174
rect 80330 222618 80566 222854
rect 64970 219218 65206 219454
rect 64970 218898 65206 219134
rect 95690 219218 95926 219454
rect 95690 218898 95926 219134
rect 109826 219218 110062 219454
rect 110146 219218 110382 219454
rect 109826 218898 110062 219134
rect 110146 218898 110382 219134
rect 60146 205538 60382 205774
rect 60466 205538 60702 205774
rect 60146 205218 60382 205454
rect 60466 205218 60702 205454
rect 80330 186938 80566 187174
rect 80330 186618 80566 186854
rect 64970 183218 65206 183454
rect 64970 182898 65206 183134
rect 95690 183218 95926 183454
rect 95690 182898 95926 183134
rect 109826 183218 110062 183454
rect 110146 183218 110382 183454
rect 109826 182898 110062 183134
rect 110146 182898 110382 183134
rect 60146 169538 60382 169774
rect 60466 169538 60702 169774
rect 60146 169218 60382 169454
rect 60466 169218 60702 169454
rect 60146 133538 60382 133774
rect 60466 133538 60702 133774
rect 60146 133218 60382 133454
rect 60466 133218 60702 133454
rect 88706 162098 88942 162334
rect 89026 162098 89262 162334
rect 88706 161778 88942 162014
rect 89026 161778 89262 162014
rect 92426 165818 92662 166054
rect 92746 165818 92982 166054
rect 92426 165498 92662 165734
rect 92746 165498 92982 165734
rect 96146 133538 96382 133774
rect 96466 133538 96702 133774
rect 96146 133218 96382 133454
rect 96466 133218 96702 133454
rect 109826 147218 110062 147454
rect 110146 147218 110382 147454
rect 109826 146898 110062 147134
rect 110146 146898 110382 147134
rect 113546 705562 113782 705798
rect 113866 705562 114102 705798
rect 113546 705242 113782 705478
rect 113866 705242 114102 705478
rect 113546 690938 113782 691174
rect 113866 690938 114102 691174
rect 113546 690618 113782 690854
rect 113866 690618 114102 690854
rect 113546 654938 113782 655174
rect 113866 654938 114102 655174
rect 113546 654618 113782 654854
rect 113866 654618 114102 654854
rect 113546 618938 113782 619174
rect 113866 618938 114102 619174
rect 113546 618618 113782 618854
rect 113866 618618 114102 618854
rect 113546 582938 113782 583174
rect 113866 582938 114102 583174
rect 113546 582618 113782 582854
rect 113866 582618 114102 582854
rect 113546 546938 113782 547174
rect 113866 546938 114102 547174
rect 113546 546618 113782 546854
rect 113866 546618 114102 546854
rect 113546 510938 113782 511174
rect 113866 510938 114102 511174
rect 113546 510618 113782 510854
rect 113866 510618 114102 510854
rect 113546 474938 113782 475174
rect 113866 474938 114102 475174
rect 113546 474618 113782 474854
rect 113866 474618 114102 474854
rect 113546 438938 113782 439174
rect 113866 438938 114102 439174
rect 113546 438618 113782 438854
rect 113866 438618 114102 438854
rect 113546 402938 113782 403174
rect 113866 402938 114102 403174
rect 113546 402618 113782 402854
rect 113866 402618 114102 402854
rect 113546 366938 113782 367174
rect 113866 366938 114102 367174
rect 113546 366618 113782 366854
rect 113866 366618 114102 366854
rect 113546 330938 113782 331174
rect 113866 330938 114102 331174
rect 113546 330618 113782 330854
rect 113866 330618 114102 330854
rect 113546 294938 113782 295174
rect 113866 294938 114102 295174
rect 113546 294618 113782 294854
rect 113866 294618 114102 294854
rect 113546 258938 113782 259174
rect 113866 258938 114102 259174
rect 113546 258618 113782 258854
rect 113866 258618 114102 258854
rect 113546 222938 113782 223174
rect 113866 222938 114102 223174
rect 113546 222618 113782 222854
rect 113866 222618 114102 222854
rect 113546 186938 113782 187174
rect 113866 186938 114102 187174
rect 113546 186618 113782 186854
rect 113866 186618 114102 186854
rect 113546 150938 113782 151174
rect 113866 150938 114102 151174
rect 113546 150618 113782 150854
rect 113866 150618 114102 150854
rect 117266 706522 117502 706758
rect 117586 706522 117822 706758
rect 117266 706202 117502 706438
rect 117586 706202 117822 706438
rect 117266 694658 117502 694894
rect 117586 694658 117822 694894
rect 117266 694338 117502 694574
rect 117586 694338 117822 694574
rect 117266 658658 117502 658894
rect 117586 658658 117822 658894
rect 117266 658338 117502 658574
rect 117586 658338 117822 658574
rect 117266 622658 117502 622894
rect 117586 622658 117822 622894
rect 117266 622338 117502 622574
rect 117586 622338 117822 622574
rect 117266 586658 117502 586894
rect 117586 586658 117822 586894
rect 117266 586338 117502 586574
rect 117586 586338 117822 586574
rect 117266 550658 117502 550894
rect 117586 550658 117822 550894
rect 117266 550338 117502 550574
rect 117586 550338 117822 550574
rect 117266 514658 117502 514894
rect 117586 514658 117822 514894
rect 117266 514338 117502 514574
rect 117586 514338 117822 514574
rect 117266 478658 117502 478894
rect 117586 478658 117822 478894
rect 117266 478338 117502 478574
rect 117586 478338 117822 478574
rect 117266 442658 117502 442894
rect 117586 442658 117822 442894
rect 117266 442338 117502 442574
rect 117586 442338 117822 442574
rect 117266 406658 117502 406894
rect 117586 406658 117822 406894
rect 117266 406338 117502 406574
rect 117586 406338 117822 406574
rect 117266 370658 117502 370894
rect 117586 370658 117822 370894
rect 117266 370338 117502 370574
rect 117586 370338 117822 370574
rect 117266 334658 117502 334894
rect 117586 334658 117822 334894
rect 117266 334338 117502 334574
rect 117586 334338 117822 334574
rect 117266 298658 117502 298894
rect 117586 298658 117822 298894
rect 117266 298338 117502 298574
rect 117586 298338 117822 298574
rect 117266 262658 117502 262894
rect 117586 262658 117822 262894
rect 117266 262338 117502 262574
rect 117586 262338 117822 262574
rect 117266 226658 117502 226894
rect 117586 226658 117822 226894
rect 117266 226338 117502 226574
rect 117586 226338 117822 226574
rect 117266 190658 117502 190894
rect 117586 190658 117822 190894
rect 117266 190338 117502 190574
rect 117586 190338 117822 190574
rect 117266 154658 117502 154894
rect 117586 154658 117822 154894
rect 117266 154338 117502 154574
rect 117586 154338 117822 154574
rect 120986 707482 121222 707718
rect 121306 707482 121542 707718
rect 120986 707162 121222 707398
rect 121306 707162 121542 707398
rect 120986 698378 121222 698614
rect 121306 698378 121542 698614
rect 120986 698058 121222 698294
rect 121306 698058 121542 698294
rect 120986 662378 121222 662614
rect 121306 662378 121542 662614
rect 120986 662058 121222 662294
rect 121306 662058 121542 662294
rect 120986 626378 121222 626614
rect 121306 626378 121542 626614
rect 120986 626058 121222 626294
rect 121306 626058 121542 626294
rect 120986 590378 121222 590614
rect 121306 590378 121542 590614
rect 120986 590058 121222 590294
rect 121306 590058 121542 590294
rect 120986 554378 121222 554614
rect 121306 554378 121542 554614
rect 120986 554058 121222 554294
rect 121306 554058 121542 554294
rect 120986 518378 121222 518614
rect 121306 518378 121542 518614
rect 120986 518058 121222 518294
rect 121306 518058 121542 518294
rect 120986 482378 121222 482614
rect 121306 482378 121542 482614
rect 120986 482058 121222 482294
rect 121306 482058 121542 482294
rect 120986 446378 121222 446614
rect 121306 446378 121542 446614
rect 120986 446058 121222 446294
rect 121306 446058 121542 446294
rect 120986 410378 121222 410614
rect 121306 410378 121542 410614
rect 120986 410058 121222 410294
rect 121306 410058 121542 410294
rect 120986 374378 121222 374614
rect 121306 374378 121542 374614
rect 120986 374058 121222 374294
rect 121306 374058 121542 374294
rect 120986 338378 121222 338614
rect 121306 338378 121542 338614
rect 120986 338058 121222 338294
rect 121306 338058 121542 338294
rect 120986 302378 121222 302614
rect 121306 302378 121542 302614
rect 120986 302058 121222 302294
rect 121306 302058 121542 302294
rect 120986 266378 121222 266614
rect 121306 266378 121542 266614
rect 120986 266058 121222 266294
rect 121306 266058 121542 266294
rect 120986 230378 121222 230614
rect 121306 230378 121542 230614
rect 120986 230058 121222 230294
rect 121306 230058 121542 230294
rect 120986 194378 121222 194614
rect 121306 194378 121542 194614
rect 120986 194058 121222 194294
rect 121306 194058 121542 194294
rect 120986 158378 121222 158614
rect 121306 158378 121542 158614
rect 120986 158058 121222 158294
rect 121306 158058 121542 158294
rect 124706 708442 124942 708678
rect 125026 708442 125262 708678
rect 124706 708122 124942 708358
rect 125026 708122 125262 708358
rect 124706 666098 124942 666334
rect 125026 666098 125262 666334
rect 124706 665778 124942 666014
rect 125026 665778 125262 666014
rect 124706 630098 124942 630334
rect 125026 630098 125262 630334
rect 124706 629778 124942 630014
rect 125026 629778 125262 630014
rect 124706 594098 124942 594334
rect 125026 594098 125262 594334
rect 124706 593778 124942 594014
rect 125026 593778 125262 594014
rect 124706 558098 124942 558334
rect 125026 558098 125262 558334
rect 124706 557778 124942 558014
rect 125026 557778 125262 558014
rect 124706 522098 124942 522334
rect 125026 522098 125262 522334
rect 124706 521778 124942 522014
rect 125026 521778 125262 522014
rect 124706 486098 124942 486334
rect 125026 486098 125262 486334
rect 124706 485778 124942 486014
rect 125026 485778 125262 486014
rect 124706 450098 124942 450334
rect 125026 450098 125262 450334
rect 124706 449778 124942 450014
rect 125026 449778 125262 450014
rect 124706 414098 124942 414334
rect 125026 414098 125262 414334
rect 124706 413778 124942 414014
rect 125026 413778 125262 414014
rect 124706 378098 124942 378334
rect 125026 378098 125262 378334
rect 124706 377778 124942 378014
rect 125026 377778 125262 378014
rect 124706 342098 124942 342334
rect 125026 342098 125262 342334
rect 124706 341778 124942 342014
rect 125026 341778 125262 342014
rect 124706 306098 124942 306334
rect 125026 306098 125262 306334
rect 124706 305778 124942 306014
rect 125026 305778 125262 306014
rect 124706 270098 124942 270334
rect 125026 270098 125262 270334
rect 124706 269778 124942 270014
rect 125026 269778 125262 270014
rect 124706 234098 124942 234334
rect 125026 234098 125262 234334
rect 124706 233778 124942 234014
rect 125026 233778 125262 234014
rect 124706 198098 124942 198334
rect 125026 198098 125262 198334
rect 124706 197778 124942 198014
rect 125026 197778 125262 198014
rect 124706 162098 124942 162334
rect 125026 162098 125262 162334
rect 124706 161778 124942 162014
rect 125026 161778 125262 162014
rect 128426 709402 128662 709638
rect 128746 709402 128982 709638
rect 128426 709082 128662 709318
rect 128746 709082 128982 709318
rect 128426 669818 128662 670054
rect 128746 669818 128982 670054
rect 128426 669498 128662 669734
rect 128746 669498 128982 669734
rect 128426 633818 128662 634054
rect 128746 633818 128982 634054
rect 128426 633498 128662 633734
rect 128746 633498 128982 633734
rect 128426 597818 128662 598054
rect 128746 597818 128982 598054
rect 128426 597498 128662 597734
rect 128746 597498 128982 597734
rect 128426 561818 128662 562054
rect 128746 561818 128982 562054
rect 128426 561498 128662 561734
rect 128746 561498 128982 561734
rect 128426 525818 128662 526054
rect 128746 525818 128982 526054
rect 128426 525498 128662 525734
rect 128746 525498 128982 525734
rect 128426 489818 128662 490054
rect 128746 489818 128982 490054
rect 128426 489498 128662 489734
rect 128746 489498 128982 489734
rect 128426 453818 128662 454054
rect 128746 453818 128982 454054
rect 128426 453498 128662 453734
rect 128746 453498 128982 453734
rect 128426 417818 128662 418054
rect 128746 417818 128982 418054
rect 128426 417498 128662 417734
rect 128746 417498 128982 417734
rect 128426 381818 128662 382054
rect 128746 381818 128982 382054
rect 128426 381498 128662 381734
rect 128746 381498 128982 381734
rect 128426 345818 128662 346054
rect 128746 345818 128982 346054
rect 128426 345498 128662 345734
rect 128746 345498 128982 345734
rect 128426 309818 128662 310054
rect 128746 309818 128982 310054
rect 128426 309498 128662 309734
rect 128746 309498 128982 309734
rect 128426 273818 128662 274054
rect 128746 273818 128982 274054
rect 128426 273498 128662 273734
rect 128746 273498 128982 273734
rect 128426 237818 128662 238054
rect 128746 237818 128982 238054
rect 128426 237498 128662 237734
rect 128746 237498 128982 237734
rect 128426 201818 128662 202054
rect 128746 201818 128982 202054
rect 128426 201498 128662 201734
rect 128746 201498 128982 201734
rect 128426 165818 128662 166054
rect 128746 165818 128982 166054
rect 128426 165498 128662 165734
rect 128746 165498 128982 165734
rect 132146 710362 132382 710598
rect 132466 710362 132702 710598
rect 132146 710042 132382 710278
rect 132466 710042 132702 710278
rect 132146 673538 132382 673774
rect 132466 673538 132702 673774
rect 132146 673218 132382 673454
rect 132466 673218 132702 673454
rect 132146 637538 132382 637774
rect 132466 637538 132702 637774
rect 132146 637218 132382 637454
rect 132466 637218 132702 637454
rect 132146 601538 132382 601774
rect 132466 601538 132702 601774
rect 132146 601218 132382 601454
rect 132466 601218 132702 601454
rect 132146 565538 132382 565774
rect 132466 565538 132702 565774
rect 132146 565218 132382 565454
rect 132466 565218 132702 565454
rect 132146 529538 132382 529774
rect 132466 529538 132702 529774
rect 132146 529218 132382 529454
rect 132466 529218 132702 529454
rect 132146 493538 132382 493774
rect 132466 493538 132702 493774
rect 132146 493218 132382 493454
rect 132466 493218 132702 493454
rect 132146 457538 132382 457774
rect 132466 457538 132702 457774
rect 132146 457218 132382 457454
rect 132466 457218 132702 457454
rect 132146 421538 132382 421774
rect 132466 421538 132702 421774
rect 132146 421218 132382 421454
rect 132466 421218 132702 421454
rect 132146 385538 132382 385774
rect 132466 385538 132702 385774
rect 132146 385218 132382 385454
rect 132466 385218 132702 385454
rect 132146 349538 132382 349774
rect 132466 349538 132702 349774
rect 132146 349218 132382 349454
rect 132466 349218 132702 349454
rect 132146 313538 132382 313774
rect 132466 313538 132702 313774
rect 132146 313218 132382 313454
rect 132466 313218 132702 313454
rect 132146 277538 132382 277774
rect 132466 277538 132702 277774
rect 132146 277218 132382 277454
rect 132466 277218 132702 277454
rect 132146 241538 132382 241774
rect 132466 241538 132702 241774
rect 132146 241218 132382 241454
rect 132466 241218 132702 241454
rect 132146 205538 132382 205774
rect 132466 205538 132702 205774
rect 132146 205218 132382 205454
rect 132466 205218 132702 205454
rect 132146 169538 132382 169774
rect 132466 169538 132702 169774
rect 132146 169218 132382 169454
rect 132466 169218 132702 169454
rect 132146 133538 132382 133774
rect 132466 133538 132702 133774
rect 132146 133218 132382 133454
rect 132466 133218 132702 133454
rect 135866 711322 136102 711558
rect 136186 711322 136422 711558
rect 135866 711002 136102 711238
rect 136186 711002 136422 711238
rect 135866 677258 136102 677494
rect 136186 677258 136422 677494
rect 135866 676938 136102 677174
rect 136186 676938 136422 677174
rect 135866 641258 136102 641494
rect 136186 641258 136422 641494
rect 135866 640938 136102 641174
rect 136186 640938 136422 641174
rect 135866 605258 136102 605494
rect 136186 605258 136422 605494
rect 135866 604938 136102 605174
rect 136186 604938 136422 605174
rect 135866 569258 136102 569494
rect 136186 569258 136422 569494
rect 135866 568938 136102 569174
rect 136186 568938 136422 569174
rect 135866 533258 136102 533494
rect 136186 533258 136422 533494
rect 135866 532938 136102 533174
rect 136186 532938 136422 533174
rect 135866 497258 136102 497494
rect 136186 497258 136422 497494
rect 135866 496938 136102 497174
rect 136186 496938 136422 497174
rect 135866 461258 136102 461494
rect 136186 461258 136422 461494
rect 135866 460938 136102 461174
rect 136186 460938 136422 461174
rect 135866 425258 136102 425494
rect 136186 425258 136422 425494
rect 135866 424938 136102 425174
rect 136186 424938 136422 425174
rect 135866 389258 136102 389494
rect 136186 389258 136422 389494
rect 135866 388938 136102 389174
rect 136186 388938 136422 389174
rect 135866 353258 136102 353494
rect 136186 353258 136422 353494
rect 135866 352938 136102 353174
rect 136186 352938 136422 353174
rect 135866 317258 136102 317494
rect 136186 317258 136422 317494
rect 135866 316938 136102 317174
rect 136186 316938 136422 317174
rect 135866 281258 136102 281494
rect 136186 281258 136422 281494
rect 135866 280938 136102 281174
rect 136186 280938 136422 281174
rect 135866 245258 136102 245494
rect 136186 245258 136422 245494
rect 135866 244938 136102 245174
rect 136186 244938 136422 245174
rect 135866 209258 136102 209494
rect 136186 209258 136422 209494
rect 135866 208938 136102 209174
rect 136186 208938 136422 209174
rect 135866 173258 136102 173494
rect 136186 173258 136422 173494
rect 135866 172938 136102 173174
rect 136186 172938 136422 173174
rect 135866 137258 136102 137494
rect 136186 137258 136422 137494
rect 135866 136938 136102 137174
rect 136186 136938 136422 137174
rect 43610 114938 43846 115174
rect 43610 114618 43846 114854
rect 74330 114938 74566 115174
rect 74330 114618 74566 114854
rect 105050 114938 105286 115174
rect 105050 114618 105286 114854
rect 28250 111218 28486 111454
rect 28250 110898 28486 111134
rect 58970 111218 59206 111454
rect 58970 110898 59206 111134
rect 89690 111218 89926 111454
rect 89690 110898 89926 111134
rect 120410 111218 120646 111454
rect 120410 110898 120646 111134
rect 24146 97538 24382 97774
rect 24466 97538 24702 97774
rect 24146 97218 24382 97454
rect 24466 97218 24702 97454
rect 135866 101258 136102 101494
rect 136186 101258 136422 101494
rect 135866 100938 136102 101174
rect 136186 100938 136422 101174
rect 43610 78938 43846 79174
rect 43610 78618 43846 78854
rect 74330 78938 74566 79174
rect 74330 78618 74566 78854
rect 105050 78938 105286 79174
rect 105050 78618 105286 78854
rect 28250 75218 28486 75454
rect 28250 74898 28486 75134
rect 58970 75218 59206 75454
rect 58970 74898 59206 75134
rect 89690 75218 89926 75454
rect 89690 74898 89926 75134
rect 120410 75218 120646 75454
rect 120410 74898 120646 75134
rect 24146 61538 24382 61774
rect 24466 61538 24702 61774
rect 24146 61218 24382 61454
rect 24466 61218 24702 61454
rect 135866 65258 136102 65494
rect 136186 65258 136422 65494
rect 135866 64938 136102 65174
rect 136186 64938 136422 65174
rect 43610 42938 43846 43174
rect 43610 42618 43846 42854
rect 74330 42938 74566 43174
rect 74330 42618 74566 42854
rect 105050 42938 105286 43174
rect 105050 42618 105286 42854
rect 28250 39218 28486 39454
rect 28250 38898 28486 39134
rect 58970 39218 59206 39454
rect 58970 38898 59206 39134
rect 89690 39218 89926 39454
rect 89690 38898 89926 39134
rect 120410 39218 120646 39454
rect 120410 38898 120646 39134
rect 24146 25538 24382 25774
rect 24466 25538 24702 25774
rect 24146 25218 24382 25454
rect 24466 25218 24702 25454
rect 135866 29258 136102 29494
rect 136186 29258 136422 29494
rect 135866 28938 136102 29174
rect 136186 28938 136422 29174
rect 24146 -6342 24382 -6106
rect 24466 -6342 24702 -6106
rect 24146 -6662 24382 -6426
rect 24466 -6662 24702 -6426
rect 37826 3218 38062 3454
rect 38146 3218 38382 3454
rect 37826 2898 38062 3134
rect 38146 2898 38382 3134
rect 37826 -582 38062 -346
rect 38146 -582 38382 -346
rect 37826 -902 38062 -666
rect 38146 -902 38382 -666
rect 41546 6938 41782 7174
rect 41866 6938 42102 7174
rect 41546 6618 41782 6854
rect 41866 6618 42102 6854
rect 41546 -1542 41782 -1306
rect 41866 -1542 42102 -1306
rect 41546 -1862 41782 -1626
rect 41866 -1862 42102 -1626
rect 45266 10658 45502 10894
rect 45586 10658 45822 10894
rect 45266 10338 45502 10574
rect 45586 10338 45822 10574
rect 45266 -2502 45502 -2266
rect 45586 -2502 45822 -2266
rect 45266 -2822 45502 -2586
rect 45586 -2822 45822 -2586
rect 48986 14378 49222 14614
rect 49306 14378 49542 14614
rect 48986 14058 49222 14294
rect 49306 14058 49542 14294
rect 48986 -3462 49222 -3226
rect 49306 -3462 49542 -3226
rect 48986 -3782 49222 -3546
rect 49306 -3782 49542 -3546
rect 52706 18098 52942 18334
rect 53026 18098 53262 18334
rect 52706 17778 52942 18014
rect 53026 17778 53262 18014
rect 52706 -4422 52942 -4186
rect 53026 -4422 53262 -4186
rect 52706 -4742 52942 -4506
rect 53026 -4742 53262 -4506
rect 56426 21818 56662 22054
rect 56746 21818 56982 22054
rect 56426 21498 56662 21734
rect 56746 21498 56982 21734
rect 56426 -5382 56662 -5146
rect 56746 -5382 56982 -5146
rect 56426 -5702 56662 -5466
rect 56746 -5702 56982 -5466
rect 73826 3218 74062 3454
rect 74146 3218 74382 3454
rect 73826 2898 74062 3134
rect 74146 2898 74382 3134
rect 73826 -582 74062 -346
rect 74146 -582 74382 -346
rect 73826 -902 74062 -666
rect 74146 -902 74382 -666
rect 77546 6938 77782 7174
rect 77866 6938 78102 7174
rect 77546 6618 77782 6854
rect 77866 6618 78102 6854
rect 77546 -1542 77782 -1306
rect 77866 -1542 78102 -1306
rect 77546 -1862 77782 -1626
rect 77866 -1862 78102 -1626
rect 81266 10658 81502 10894
rect 81586 10658 81822 10894
rect 81266 10338 81502 10574
rect 81586 10338 81822 10574
rect 81266 -2502 81502 -2266
rect 81586 -2502 81822 -2266
rect 81266 -2822 81502 -2586
rect 81586 -2822 81822 -2586
rect 84986 14378 85222 14614
rect 85306 14378 85542 14614
rect 84986 14058 85222 14294
rect 85306 14058 85542 14294
rect 84986 -3462 85222 -3226
rect 85306 -3462 85542 -3226
rect 84986 -3782 85222 -3546
rect 85306 -3782 85542 -3546
rect 88706 18098 88942 18334
rect 89026 18098 89262 18334
rect 88706 17778 88942 18014
rect 89026 17778 89262 18014
rect 88706 -4422 88942 -4186
rect 89026 -4422 89262 -4186
rect 88706 -4742 88942 -4506
rect 89026 -4742 89262 -4506
rect 92426 21818 92662 22054
rect 92746 21818 92982 22054
rect 92426 21498 92662 21734
rect 92746 21498 92982 21734
rect 92426 -5382 92662 -5146
rect 92746 -5382 92982 -5146
rect 92426 -5702 92662 -5466
rect 92746 -5702 92982 -5466
rect 109826 3218 110062 3454
rect 110146 3218 110382 3454
rect 109826 2898 110062 3134
rect 110146 2898 110382 3134
rect 109826 -582 110062 -346
rect 110146 -582 110382 -346
rect 109826 -902 110062 -666
rect 110146 -902 110382 -666
rect 113546 6938 113782 7174
rect 113866 6938 114102 7174
rect 113546 6618 113782 6854
rect 113866 6618 114102 6854
rect 113546 -1542 113782 -1306
rect 113866 -1542 114102 -1306
rect 113546 -1862 113782 -1626
rect 113866 -1862 114102 -1626
rect 117266 10658 117502 10894
rect 117586 10658 117822 10894
rect 117266 10338 117502 10574
rect 117586 10338 117822 10574
rect 117266 -2502 117502 -2266
rect 117586 -2502 117822 -2266
rect 117266 -2822 117502 -2586
rect 117586 -2822 117822 -2586
rect 120986 14378 121222 14614
rect 121306 14378 121542 14614
rect 120986 14058 121222 14294
rect 121306 14058 121542 14294
rect 120986 -3462 121222 -3226
rect 121306 -3462 121542 -3226
rect 120986 -3782 121222 -3546
rect 121306 -3782 121542 -3546
rect 124706 18098 124942 18334
rect 125026 18098 125262 18334
rect 124706 17778 124942 18014
rect 125026 17778 125262 18014
rect 124706 -4422 124942 -4186
rect 125026 -4422 125262 -4186
rect 124706 -4742 124942 -4506
rect 125026 -4742 125262 -4506
rect 128426 21818 128662 22054
rect 128746 21818 128982 22054
rect 128426 21498 128662 21734
rect 128746 21498 128982 21734
rect 128426 -5382 128662 -5146
rect 128746 -5382 128982 -5146
rect 128426 -5702 128662 -5466
rect 128746 -5702 128982 -5466
rect 135866 -7302 136102 -7066
rect 136186 -7302 136422 -7066
rect 135866 -7622 136102 -7386
rect 136186 -7622 136422 -7386
rect 145826 704602 146062 704838
rect 146146 704602 146382 704838
rect 145826 704282 146062 704518
rect 146146 704282 146382 704518
rect 145826 687218 146062 687454
rect 146146 687218 146382 687454
rect 145826 686898 146062 687134
rect 146146 686898 146382 687134
rect 145826 651218 146062 651454
rect 146146 651218 146382 651454
rect 145826 650898 146062 651134
rect 146146 650898 146382 651134
rect 145826 615218 146062 615454
rect 146146 615218 146382 615454
rect 145826 614898 146062 615134
rect 146146 614898 146382 615134
rect 145826 579218 146062 579454
rect 146146 579218 146382 579454
rect 145826 578898 146062 579134
rect 146146 578898 146382 579134
rect 145826 543218 146062 543454
rect 146146 543218 146382 543454
rect 145826 542898 146062 543134
rect 146146 542898 146382 543134
rect 145826 507218 146062 507454
rect 146146 507218 146382 507454
rect 145826 506898 146062 507134
rect 146146 506898 146382 507134
rect 145826 471218 146062 471454
rect 146146 471218 146382 471454
rect 145826 470898 146062 471134
rect 146146 470898 146382 471134
rect 145826 435218 146062 435454
rect 146146 435218 146382 435454
rect 145826 434898 146062 435134
rect 146146 434898 146382 435134
rect 145826 399218 146062 399454
rect 146146 399218 146382 399454
rect 145826 398898 146062 399134
rect 146146 398898 146382 399134
rect 145826 363218 146062 363454
rect 146146 363218 146382 363454
rect 145826 362898 146062 363134
rect 146146 362898 146382 363134
rect 145826 327218 146062 327454
rect 146146 327218 146382 327454
rect 145826 326898 146062 327134
rect 146146 326898 146382 327134
rect 145826 291218 146062 291454
rect 146146 291218 146382 291454
rect 145826 290898 146062 291134
rect 146146 290898 146382 291134
rect 145826 255218 146062 255454
rect 146146 255218 146382 255454
rect 145826 254898 146062 255134
rect 146146 254898 146382 255134
rect 145826 219218 146062 219454
rect 146146 219218 146382 219454
rect 145826 218898 146062 219134
rect 146146 218898 146382 219134
rect 145826 183218 146062 183454
rect 146146 183218 146382 183454
rect 145826 182898 146062 183134
rect 146146 182898 146382 183134
rect 145826 147218 146062 147454
rect 146146 147218 146382 147454
rect 145826 146898 146062 147134
rect 146146 146898 146382 147134
rect 145826 111218 146062 111454
rect 146146 111218 146382 111454
rect 145826 110898 146062 111134
rect 146146 110898 146382 111134
rect 145826 75218 146062 75454
rect 146146 75218 146382 75454
rect 145826 74898 146062 75134
rect 146146 74898 146382 75134
rect 145826 39218 146062 39454
rect 146146 39218 146382 39454
rect 145826 38898 146062 39134
rect 146146 38898 146382 39134
rect 145826 3218 146062 3454
rect 146146 3218 146382 3454
rect 145826 2898 146062 3134
rect 146146 2898 146382 3134
rect 145826 -582 146062 -346
rect 146146 -582 146382 -346
rect 145826 -902 146062 -666
rect 146146 -902 146382 -666
rect 149546 705562 149782 705798
rect 149866 705562 150102 705798
rect 149546 705242 149782 705478
rect 149866 705242 150102 705478
rect 149546 690938 149782 691174
rect 149866 690938 150102 691174
rect 149546 690618 149782 690854
rect 149866 690618 150102 690854
rect 149546 654938 149782 655174
rect 149866 654938 150102 655174
rect 149546 654618 149782 654854
rect 149866 654618 150102 654854
rect 149546 618938 149782 619174
rect 149866 618938 150102 619174
rect 149546 618618 149782 618854
rect 149866 618618 150102 618854
rect 149546 582938 149782 583174
rect 149866 582938 150102 583174
rect 149546 582618 149782 582854
rect 149866 582618 150102 582854
rect 149546 546938 149782 547174
rect 149866 546938 150102 547174
rect 149546 546618 149782 546854
rect 149866 546618 150102 546854
rect 149546 510938 149782 511174
rect 149866 510938 150102 511174
rect 149546 510618 149782 510854
rect 149866 510618 150102 510854
rect 149546 474938 149782 475174
rect 149866 474938 150102 475174
rect 149546 474618 149782 474854
rect 149866 474618 150102 474854
rect 149546 438938 149782 439174
rect 149866 438938 150102 439174
rect 149546 438618 149782 438854
rect 149866 438618 150102 438854
rect 149546 402938 149782 403174
rect 149866 402938 150102 403174
rect 149546 402618 149782 402854
rect 149866 402618 150102 402854
rect 149546 366938 149782 367174
rect 149866 366938 150102 367174
rect 149546 366618 149782 366854
rect 149866 366618 150102 366854
rect 149546 330938 149782 331174
rect 149866 330938 150102 331174
rect 149546 330618 149782 330854
rect 149866 330618 150102 330854
rect 149546 294938 149782 295174
rect 149866 294938 150102 295174
rect 149546 294618 149782 294854
rect 149866 294618 150102 294854
rect 149546 258938 149782 259174
rect 149866 258938 150102 259174
rect 149546 258618 149782 258854
rect 149866 258618 150102 258854
rect 149546 222938 149782 223174
rect 149866 222938 150102 223174
rect 149546 222618 149782 222854
rect 149866 222618 150102 222854
rect 149546 186938 149782 187174
rect 149866 186938 150102 187174
rect 149546 186618 149782 186854
rect 149866 186618 150102 186854
rect 149546 150938 149782 151174
rect 149866 150938 150102 151174
rect 149546 150618 149782 150854
rect 149866 150618 150102 150854
rect 149546 114938 149782 115174
rect 149866 114938 150102 115174
rect 149546 114618 149782 114854
rect 149866 114618 150102 114854
rect 149546 78938 149782 79174
rect 149866 78938 150102 79174
rect 149546 78618 149782 78854
rect 149866 78618 150102 78854
rect 149546 42938 149782 43174
rect 149866 42938 150102 43174
rect 149546 42618 149782 42854
rect 149866 42618 150102 42854
rect 149546 6938 149782 7174
rect 149866 6938 150102 7174
rect 149546 6618 149782 6854
rect 149866 6618 150102 6854
rect 149546 -1542 149782 -1306
rect 149866 -1542 150102 -1306
rect 149546 -1862 149782 -1626
rect 149866 -1862 150102 -1626
rect 153266 706522 153502 706758
rect 153586 706522 153822 706758
rect 153266 706202 153502 706438
rect 153586 706202 153822 706438
rect 153266 694658 153502 694894
rect 153586 694658 153822 694894
rect 153266 694338 153502 694574
rect 153586 694338 153822 694574
rect 153266 658658 153502 658894
rect 153586 658658 153822 658894
rect 153266 658338 153502 658574
rect 153586 658338 153822 658574
rect 153266 622658 153502 622894
rect 153586 622658 153822 622894
rect 153266 622338 153502 622574
rect 153586 622338 153822 622574
rect 153266 586658 153502 586894
rect 153586 586658 153822 586894
rect 153266 586338 153502 586574
rect 153586 586338 153822 586574
rect 153266 550658 153502 550894
rect 153586 550658 153822 550894
rect 153266 550338 153502 550574
rect 153586 550338 153822 550574
rect 153266 514658 153502 514894
rect 153586 514658 153822 514894
rect 153266 514338 153502 514574
rect 153586 514338 153822 514574
rect 153266 478658 153502 478894
rect 153586 478658 153822 478894
rect 153266 478338 153502 478574
rect 153586 478338 153822 478574
rect 153266 442658 153502 442894
rect 153586 442658 153822 442894
rect 153266 442338 153502 442574
rect 153586 442338 153822 442574
rect 156986 707482 157222 707718
rect 157306 707482 157542 707718
rect 156986 707162 157222 707398
rect 157306 707162 157542 707398
rect 156986 698378 157222 698614
rect 157306 698378 157542 698614
rect 156986 698058 157222 698294
rect 157306 698058 157542 698294
rect 156986 662378 157222 662614
rect 157306 662378 157542 662614
rect 156986 662058 157222 662294
rect 157306 662058 157542 662294
rect 156986 626378 157222 626614
rect 157306 626378 157542 626614
rect 156986 626058 157222 626294
rect 157306 626058 157542 626294
rect 156986 590378 157222 590614
rect 157306 590378 157542 590614
rect 156986 590058 157222 590294
rect 157306 590058 157542 590294
rect 156986 554378 157222 554614
rect 157306 554378 157542 554614
rect 156986 554058 157222 554294
rect 157306 554058 157542 554294
rect 156986 518378 157222 518614
rect 157306 518378 157542 518614
rect 156986 518058 157222 518294
rect 157306 518058 157542 518294
rect 156986 482378 157222 482614
rect 157306 482378 157542 482614
rect 156986 482058 157222 482294
rect 157306 482058 157542 482294
rect 156986 446378 157222 446614
rect 157306 446378 157542 446614
rect 156986 446058 157222 446294
rect 157306 446058 157542 446294
rect 160706 708442 160942 708678
rect 161026 708442 161262 708678
rect 160706 708122 160942 708358
rect 161026 708122 161262 708358
rect 160706 666098 160942 666334
rect 161026 666098 161262 666334
rect 160706 665778 160942 666014
rect 161026 665778 161262 666014
rect 160706 630098 160942 630334
rect 161026 630098 161262 630334
rect 160706 629778 160942 630014
rect 161026 629778 161262 630014
rect 160706 594098 160942 594334
rect 161026 594098 161262 594334
rect 160706 593778 160942 594014
rect 161026 593778 161262 594014
rect 160706 558098 160942 558334
rect 161026 558098 161262 558334
rect 160706 557778 160942 558014
rect 161026 557778 161262 558014
rect 160706 522098 160942 522334
rect 161026 522098 161262 522334
rect 160706 521778 160942 522014
rect 161026 521778 161262 522014
rect 160706 486098 160942 486334
rect 161026 486098 161262 486334
rect 160706 485778 160942 486014
rect 161026 485778 161262 486014
rect 160706 450098 160942 450334
rect 161026 450098 161262 450334
rect 160706 449778 160942 450014
rect 161026 449778 161262 450014
rect 164426 709402 164662 709638
rect 164746 709402 164982 709638
rect 164426 709082 164662 709318
rect 164746 709082 164982 709318
rect 164426 669818 164662 670054
rect 164746 669818 164982 670054
rect 164426 669498 164662 669734
rect 164746 669498 164982 669734
rect 164426 633818 164662 634054
rect 164746 633818 164982 634054
rect 164426 633498 164662 633734
rect 164746 633498 164982 633734
rect 164426 597818 164662 598054
rect 164746 597818 164982 598054
rect 164426 597498 164662 597734
rect 164746 597498 164982 597734
rect 164426 561818 164662 562054
rect 164746 561818 164982 562054
rect 164426 561498 164662 561734
rect 164746 561498 164982 561734
rect 164426 525818 164662 526054
rect 164746 525818 164982 526054
rect 164426 525498 164662 525734
rect 164746 525498 164982 525734
rect 164426 489818 164662 490054
rect 164746 489818 164982 490054
rect 164426 489498 164662 489734
rect 164746 489498 164982 489734
rect 164426 453818 164662 454054
rect 164746 453818 164982 454054
rect 164426 453498 164662 453734
rect 164746 453498 164982 453734
rect 168146 710362 168382 710598
rect 168466 710362 168702 710598
rect 168146 710042 168382 710278
rect 168466 710042 168702 710278
rect 168146 673538 168382 673774
rect 168466 673538 168702 673774
rect 168146 673218 168382 673454
rect 168466 673218 168702 673454
rect 168146 637538 168382 637774
rect 168466 637538 168702 637774
rect 168146 637218 168382 637454
rect 168466 637218 168702 637454
rect 168146 601538 168382 601774
rect 168466 601538 168702 601774
rect 168146 601218 168382 601454
rect 168466 601218 168702 601454
rect 168146 565538 168382 565774
rect 168466 565538 168702 565774
rect 168146 565218 168382 565454
rect 168466 565218 168702 565454
rect 168146 529538 168382 529774
rect 168466 529538 168702 529774
rect 168146 529218 168382 529454
rect 168466 529218 168702 529454
rect 168146 493538 168382 493774
rect 168466 493538 168702 493774
rect 168146 493218 168382 493454
rect 168466 493218 168702 493454
rect 168146 457538 168382 457774
rect 168466 457538 168702 457774
rect 168146 457218 168382 457454
rect 168466 457218 168702 457454
rect 171866 711322 172102 711558
rect 172186 711322 172422 711558
rect 171866 711002 172102 711238
rect 172186 711002 172422 711238
rect 171866 677258 172102 677494
rect 172186 677258 172422 677494
rect 171866 676938 172102 677174
rect 172186 676938 172422 677174
rect 171866 641258 172102 641494
rect 172186 641258 172422 641494
rect 171866 640938 172102 641174
rect 172186 640938 172422 641174
rect 171866 605258 172102 605494
rect 172186 605258 172422 605494
rect 171866 604938 172102 605174
rect 172186 604938 172422 605174
rect 171866 569258 172102 569494
rect 172186 569258 172422 569494
rect 171866 568938 172102 569174
rect 172186 568938 172422 569174
rect 171866 533258 172102 533494
rect 172186 533258 172422 533494
rect 171866 532938 172102 533174
rect 172186 532938 172422 533174
rect 171866 497258 172102 497494
rect 172186 497258 172422 497494
rect 171866 496938 172102 497174
rect 172186 496938 172422 497174
rect 171866 461258 172102 461494
rect 172186 461258 172422 461494
rect 171866 460938 172102 461174
rect 172186 460938 172422 461174
rect 171866 425258 172102 425494
rect 172186 425258 172422 425494
rect 171866 424938 172102 425174
rect 172186 424938 172422 425174
rect 181826 704602 182062 704838
rect 182146 704602 182382 704838
rect 181826 704282 182062 704518
rect 182146 704282 182382 704518
rect 181826 687218 182062 687454
rect 182146 687218 182382 687454
rect 181826 686898 182062 687134
rect 182146 686898 182382 687134
rect 181826 651218 182062 651454
rect 182146 651218 182382 651454
rect 181826 650898 182062 651134
rect 182146 650898 182382 651134
rect 181826 615218 182062 615454
rect 182146 615218 182382 615454
rect 181826 614898 182062 615134
rect 182146 614898 182382 615134
rect 181826 579218 182062 579454
rect 182146 579218 182382 579454
rect 181826 578898 182062 579134
rect 182146 578898 182382 579134
rect 181826 543218 182062 543454
rect 182146 543218 182382 543454
rect 181826 542898 182062 543134
rect 182146 542898 182382 543134
rect 181826 507218 182062 507454
rect 182146 507218 182382 507454
rect 181826 506898 182062 507134
rect 182146 506898 182382 507134
rect 181826 471218 182062 471454
rect 182146 471218 182382 471454
rect 181826 470898 182062 471134
rect 182146 470898 182382 471134
rect 181826 435218 182062 435454
rect 182146 435218 182382 435454
rect 181826 434898 182062 435134
rect 182146 434898 182382 435134
rect 185546 705562 185782 705798
rect 185866 705562 186102 705798
rect 185546 705242 185782 705478
rect 185866 705242 186102 705478
rect 185546 690938 185782 691174
rect 185866 690938 186102 691174
rect 185546 690618 185782 690854
rect 185866 690618 186102 690854
rect 185546 654938 185782 655174
rect 185866 654938 186102 655174
rect 185546 654618 185782 654854
rect 185866 654618 186102 654854
rect 185546 618938 185782 619174
rect 185866 618938 186102 619174
rect 185546 618618 185782 618854
rect 185866 618618 186102 618854
rect 185546 582938 185782 583174
rect 185866 582938 186102 583174
rect 185546 582618 185782 582854
rect 185866 582618 186102 582854
rect 185546 546938 185782 547174
rect 185866 546938 186102 547174
rect 185546 546618 185782 546854
rect 185866 546618 186102 546854
rect 185546 510938 185782 511174
rect 185866 510938 186102 511174
rect 185546 510618 185782 510854
rect 185866 510618 186102 510854
rect 185546 474938 185782 475174
rect 185866 474938 186102 475174
rect 185546 474618 185782 474854
rect 185866 474618 186102 474854
rect 185546 438938 185782 439174
rect 185866 438938 186102 439174
rect 185546 438618 185782 438854
rect 185866 438618 186102 438854
rect 189266 706522 189502 706758
rect 189586 706522 189822 706758
rect 189266 706202 189502 706438
rect 189586 706202 189822 706438
rect 189266 694658 189502 694894
rect 189586 694658 189822 694894
rect 189266 694338 189502 694574
rect 189586 694338 189822 694574
rect 189266 658658 189502 658894
rect 189586 658658 189822 658894
rect 189266 658338 189502 658574
rect 189586 658338 189822 658574
rect 189266 622658 189502 622894
rect 189586 622658 189822 622894
rect 189266 622338 189502 622574
rect 189586 622338 189822 622574
rect 189266 586658 189502 586894
rect 189586 586658 189822 586894
rect 189266 586338 189502 586574
rect 189586 586338 189822 586574
rect 189266 550658 189502 550894
rect 189586 550658 189822 550894
rect 189266 550338 189502 550574
rect 189586 550338 189822 550574
rect 189266 514658 189502 514894
rect 189586 514658 189822 514894
rect 189266 514338 189502 514574
rect 189586 514338 189822 514574
rect 189266 478658 189502 478894
rect 189586 478658 189822 478894
rect 189266 478338 189502 478574
rect 189586 478338 189822 478574
rect 189266 442658 189502 442894
rect 189586 442658 189822 442894
rect 189266 442338 189502 442574
rect 189586 442338 189822 442574
rect 192986 707482 193222 707718
rect 193306 707482 193542 707718
rect 192986 707162 193222 707398
rect 193306 707162 193542 707398
rect 192986 698378 193222 698614
rect 193306 698378 193542 698614
rect 192986 698058 193222 698294
rect 193306 698058 193542 698294
rect 192986 662378 193222 662614
rect 193306 662378 193542 662614
rect 192986 662058 193222 662294
rect 193306 662058 193542 662294
rect 192986 626378 193222 626614
rect 193306 626378 193542 626614
rect 192986 626058 193222 626294
rect 193306 626058 193542 626294
rect 192986 590378 193222 590614
rect 193306 590378 193542 590614
rect 192986 590058 193222 590294
rect 193306 590058 193542 590294
rect 192986 554378 193222 554614
rect 193306 554378 193542 554614
rect 192986 554058 193222 554294
rect 193306 554058 193542 554294
rect 192986 518378 193222 518614
rect 193306 518378 193542 518614
rect 192986 518058 193222 518294
rect 193306 518058 193542 518294
rect 192986 482378 193222 482614
rect 193306 482378 193542 482614
rect 192986 482058 193222 482294
rect 193306 482058 193542 482294
rect 192986 446378 193222 446614
rect 193306 446378 193542 446614
rect 192986 446058 193222 446294
rect 193306 446058 193542 446294
rect 196706 708442 196942 708678
rect 197026 708442 197262 708678
rect 196706 708122 196942 708358
rect 197026 708122 197262 708358
rect 196706 666098 196942 666334
rect 197026 666098 197262 666334
rect 196706 665778 196942 666014
rect 197026 665778 197262 666014
rect 196706 630098 196942 630334
rect 197026 630098 197262 630334
rect 196706 629778 196942 630014
rect 197026 629778 197262 630014
rect 196706 594098 196942 594334
rect 197026 594098 197262 594334
rect 196706 593778 196942 594014
rect 197026 593778 197262 594014
rect 196706 558098 196942 558334
rect 197026 558098 197262 558334
rect 196706 557778 196942 558014
rect 197026 557778 197262 558014
rect 196706 522098 196942 522334
rect 197026 522098 197262 522334
rect 196706 521778 196942 522014
rect 197026 521778 197262 522014
rect 196706 486098 196942 486334
rect 197026 486098 197262 486334
rect 196706 485778 196942 486014
rect 197026 485778 197262 486014
rect 196706 450098 196942 450334
rect 197026 450098 197262 450334
rect 196706 449778 196942 450014
rect 197026 449778 197262 450014
rect 200426 709402 200662 709638
rect 200746 709402 200982 709638
rect 200426 709082 200662 709318
rect 200746 709082 200982 709318
rect 200426 669818 200662 670054
rect 200746 669818 200982 670054
rect 200426 669498 200662 669734
rect 200746 669498 200982 669734
rect 200426 633818 200662 634054
rect 200746 633818 200982 634054
rect 200426 633498 200662 633734
rect 200746 633498 200982 633734
rect 200426 597818 200662 598054
rect 200746 597818 200982 598054
rect 200426 597498 200662 597734
rect 200746 597498 200982 597734
rect 200426 561818 200662 562054
rect 200746 561818 200982 562054
rect 200426 561498 200662 561734
rect 200746 561498 200982 561734
rect 200426 525818 200662 526054
rect 200746 525818 200982 526054
rect 200426 525498 200662 525734
rect 200746 525498 200982 525734
rect 200426 489818 200662 490054
rect 200746 489818 200982 490054
rect 200426 489498 200662 489734
rect 200746 489498 200982 489734
rect 200426 453818 200662 454054
rect 200746 453818 200982 454054
rect 200426 453498 200662 453734
rect 200746 453498 200982 453734
rect 204146 710362 204382 710598
rect 204466 710362 204702 710598
rect 204146 710042 204382 710278
rect 204466 710042 204702 710278
rect 204146 673538 204382 673774
rect 204466 673538 204702 673774
rect 204146 673218 204382 673454
rect 204466 673218 204702 673454
rect 204146 637538 204382 637774
rect 204466 637538 204702 637774
rect 204146 637218 204382 637454
rect 204466 637218 204702 637454
rect 204146 601538 204382 601774
rect 204466 601538 204702 601774
rect 204146 601218 204382 601454
rect 204466 601218 204702 601454
rect 204146 565538 204382 565774
rect 204466 565538 204702 565774
rect 204146 565218 204382 565454
rect 204466 565218 204702 565454
rect 204146 529538 204382 529774
rect 204466 529538 204702 529774
rect 204146 529218 204382 529454
rect 204466 529218 204702 529454
rect 204146 493538 204382 493774
rect 204466 493538 204702 493774
rect 204146 493218 204382 493454
rect 204466 493218 204702 493454
rect 204146 457538 204382 457774
rect 204466 457538 204702 457774
rect 204146 457218 204382 457454
rect 204466 457218 204702 457454
rect 207866 711322 208102 711558
rect 208186 711322 208422 711558
rect 207866 711002 208102 711238
rect 208186 711002 208422 711238
rect 207866 677258 208102 677494
rect 208186 677258 208422 677494
rect 207866 676938 208102 677174
rect 208186 676938 208422 677174
rect 207866 641258 208102 641494
rect 208186 641258 208422 641494
rect 207866 640938 208102 641174
rect 208186 640938 208422 641174
rect 207866 605258 208102 605494
rect 208186 605258 208422 605494
rect 207866 604938 208102 605174
rect 208186 604938 208422 605174
rect 207866 569258 208102 569494
rect 208186 569258 208422 569494
rect 207866 568938 208102 569174
rect 208186 568938 208422 569174
rect 207866 533258 208102 533494
rect 208186 533258 208422 533494
rect 207866 532938 208102 533174
rect 208186 532938 208422 533174
rect 207866 497258 208102 497494
rect 208186 497258 208422 497494
rect 207866 496938 208102 497174
rect 208186 496938 208422 497174
rect 207866 461258 208102 461494
rect 208186 461258 208422 461494
rect 207866 460938 208102 461174
rect 208186 460938 208422 461174
rect 217826 704602 218062 704838
rect 218146 704602 218382 704838
rect 217826 704282 218062 704518
rect 218146 704282 218382 704518
rect 217826 687218 218062 687454
rect 218146 687218 218382 687454
rect 217826 686898 218062 687134
rect 218146 686898 218382 687134
rect 217826 651218 218062 651454
rect 218146 651218 218382 651454
rect 217826 650898 218062 651134
rect 218146 650898 218382 651134
rect 217826 615218 218062 615454
rect 218146 615218 218382 615454
rect 217826 614898 218062 615134
rect 218146 614898 218382 615134
rect 217826 579218 218062 579454
rect 218146 579218 218382 579454
rect 217826 578898 218062 579134
rect 218146 578898 218382 579134
rect 217826 543218 218062 543454
rect 218146 543218 218382 543454
rect 217826 542898 218062 543134
rect 218146 542898 218382 543134
rect 217826 507218 218062 507454
rect 218146 507218 218382 507454
rect 217826 506898 218062 507134
rect 218146 506898 218382 507134
rect 217826 471218 218062 471454
rect 218146 471218 218382 471454
rect 217826 470898 218062 471134
rect 218146 470898 218382 471134
rect 217826 435218 218062 435454
rect 218146 435218 218382 435454
rect 217826 434898 218062 435134
rect 218146 434898 218382 435134
rect 153266 406658 153502 406894
rect 153586 406658 153822 406894
rect 153266 406338 153502 406574
rect 153586 406338 153822 406574
rect 177610 402938 177846 403174
rect 177610 402618 177846 402854
rect 208330 402938 208566 403174
rect 208330 402618 208566 402854
rect 162250 399218 162486 399454
rect 162250 398898 162486 399134
rect 192970 399218 193206 399454
rect 192970 398898 193206 399134
rect 217826 399218 218062 399454
rect 218146 399218 218382 399454
rect 217826 398898 218062 399134
rect 218146 398898 218382 399134
rect 153266 370658 153502 370894
rect 153586 370658 153822 370894
rect 153266 370338 153502 370574
rect 153586 370338 153822 370574
rect 177610 366938 177846 367174
rect 177610 366618 177846 366854
rect 208330 366938 208566 367174
rect 208330 366618 208566 366854
rect 162250 363218 162486 363454
rect 162250 362898 162486 363134
rect 192970 363218 193206 363454
rect 192970 362898 193206 363134
rect 217826 363218 218062 363454
rect 218146 363218 218382 363454
rect 217826 362898 218062 363134
rect 218146 362898 218382 363134
rect 153266 334658 153502 334894
rect 153586 334658 153822 334894
rect 153266 334338 153502 334574
rect 153586 334338 153822 334574
rect 177610 330938 177846 331174
rect 177610 330618 177846 330854
rect 208330 330938 208566 331174
rect 208330 330618 208566 330854
rect 162250 327218 162486 327454
rect 162250 326898 162486 327134
rect 192970 327218 193206 327454
rect 192970 326898 193206 327134
rect 217826 327218 218062 327454
rect 218146 327218 218382 327454
rect 217826 326898 218062 327134
rect 218146 326898 218382 327134
rect 153266 298658 153502 298894
rect 153586 298658 153822 298894
rect 153266 298338 153502 298574
rect 153586 298338 153822 298574
rect 177610 294938 177846 295174
rect 177610 294618 177846 294854
rect 208330 294938 208566 295174
rect 208330 294618 208566 294854
rect 153266 262658 153502 262894
rect 153586 262658 153822 262894
rect 153266 262338 153502 262574
rect 153586 262338 153822 262574
rect 153266 226658 153502 226894
rect 153586 226658 153822 226894
rect 153266 226338 153502 226574
rect 153586 226338 153822 226574
rect 153266 190658 153502 190894
rect 153586 190658 153822 190894
rect 153266 190338 153502 190574
rect 153586 190338 153822 190574
rect 162250 291218 162486 291454
rect 162250 290898 162486 291134
rect 192970 291218 193206 291454
rect 192970 290898 193206 291134
rect 217826 291218 218062 291454
rect 218146 291218 218382 291454
rect 217826 290898 218062 291134
rect 218146 290898 218382 291134
rect 156986 266378 157222 266614
rect 157306 266378 157542 266614
rect 156986 266058 157222 266294
rect 157306 266058 157542 266294
rect 156986 230378 157222 230614
rect 157306 230378 157542 230614
rect 156986 230058 157222 230294
rect 157306 230058 157542 230294
rect 156986 194378 157222 194614
rect 157306 194378 157542 194614
rect 156986 194058 157222 194294
rect 157306 194058 157542 194294
rect 153266 154658 153502 154894
rect 153586 154658 153822 154894
rect 153266 154338 153502 154574
rect 153586 154338 153822 154574
rect 153266 118658 153502 118894
rect 153586 118658 153822 118894
rect 153266 118338 153502 118574
rect 153586 118338 153822 118574
rect 153266 82658 153502 82894
rect 153586 82658 153822 82894
rect 153266 82338 153502 82574
rect 153586 82338 153822 82574
rect 153266 46658 153502 46894
rect 153586 46658 153822 46894
rect 153266 46338 153502 46574
rect 153586 46338 153822 46574
rect 153266 10658 153502 10894
rect 153586 10658 153822 10894
rect 153266 10338 153502 10574
rect 153586 10338 153822 10574
rect 153266 -2502 153502 -2266
rect 153586 -2502 153822 -2266
rect 153266 -2822 153502 -2586
rect 153586 -2822 153822 -2586
rect 156986 158378 157222 158614
rect 157306 158378 157542 158614
rect 156986 158058 157222 158294
rect 157306 158058 157542 158294
rect 160706 234098 160942 234334
rect 161026 234098 161262 234334
rect 160706 233778 160942 234014
rect 161026 233778 161262 234014
rect 160706 198098 160942 198334
rect 161026 198098 161262 198334
rect 160706 197778 160942 198014
rect 161026 197778 161262 198014
rect 160706 162098 160942 162334
rect 161026 162098 161262 162334
rect 160706 161778 160942 162014
rect 161026 161778 161262 162014
rect 164426 237818 164662 238054
rect 164746 237818 164982 238054
rect 164426 237498 164662 237734
rect 164746 237498 164982 237734
rect 164426 201818 164662 202054
rect 164746 201818 164982 202054
rect 164426 201498 164662 201734
rect 164746 201498 164982 201734
rect 164426 165818 164662 166054
rect 164746 165818 164982 166054
rect 164426 165498 164662 165734
rect 164746 165498 164982 165734
rect 168146 241538 168382 241774
rect 168466 241538 168702 241774
rect 168146 241218 168382 241454
rect 168466 241218 168702 241454
rect 168146 205538 168382 205774
rect 168466 205538 168702 205774
rect 168146 205218 168382 205454
rect 168466 205218 168702 205454
rect 168146 169538 168382 169774
rect 168466 169538 168702 169774
rect 168146 169218 168382 169454
rect 168466 169218 168702 169454
rect 168146 133538 168382 133774
rect 168466 133538 168702 133774
rect 168146 133218 168382 133454
rect 168466 133218 168702 133454
rect 171866 245258 172102 245494
rect 172186 245258 172422 245494
rect 171866 244938 172102 245174
rect 172186 244938 172422 245174
rect 171866 209258 172102 209494
rect 172186 209258 172422 209494
rect 171866 208938 172102 209174
rect 172186 208938 172422 209174
rect 171866 173258 172102 173494
rect 172186 173258 172422 173494
rect 171866 172938 172102 173174
rect 172186 172938 172422 173174
rect 171866 137258 172102 137494
rect 172186 137258 172422 137494
rect 171866 136938 172102 137174
rect 172186 136938 172422 137174
rect 181826 255218 182062 255454
rect 182146 255218 182382 255454
rect 181826 254898 182062 255134
rect 182146 254898 182382 255134
rect 181826 219218 182062 219454
rect 182146 219218 182382 219454
rect 181826 218898 182062 219134
rect 182146 218898 182382 219134
rect 181826 183218 182062 183454
rect 182146 183218 182382 183454
rect 181826 182898 182062 183134
rect 182146 182898 182382 183134
rect 181826 147218 182062 147454
rect 182146 147218 182382 147454
rect 181826 146898 182062 147134
rect 182146 146898 182382 147134
rect 185546 258938 185782 259174
rect 185866 258938 186102 259174
rect 185546 258618 185782 258854
rect 185866 258618 186102 258854
rect 185546 222938 185782 223174
rect 185866 222938 186102 223174
rect 185546 222618 185782 222854
rect 185866 222618 186102 222854
rect 185546 186938 185782 187174
rect 185866 186938 186102 187174
rect 185546 186618 185782 186854
rect 185866 186618 186102 186854
rect 185546 150938 185782 151174
rect 185866 150938 186102 151174
rect 185546 150618 185782 150854
rect 185866 150618 186102 150854
rect 189266 262658 189502 262894
rect 189586 262658 189822 262894
rect 189266 262338 189502 262574
rect 189586 262338 189822 262574
rect 189266 226658 189502 226894
rect 189586 226658 189822 226894
rect 189266 226338 189502 226574
rect 189586 226338 189822 226574
rect 189266 190658 189502 190894
rect 189586 190658 189822 190894
rect 189266 190338 189502 190574
rect 189586 190338 189822 190574
rect 189266 154658 189502 154894
rect 189586 154658 189822 154894
rect 189266 154338 189502 154574
rect 189586 154338 189822 154574
rect 192986 266378 193222 266614
rect 193306 266378 193542 266614
rect 192986 266058 193222 266294
rect 193306 266058 193542 266294
rect 192986 230378 193222 230614
rect 193306 230378 193542 230614
rect 192986 230058 193222 230294
rect 193306 230058 193542 230294
rect 192986 194378 193222 194614
rect 193306 194378 193542 194614
rect 192986 194058 193222 194294
rect 193306 194058 193542 194294
rect 192986 158378 193222 158614
rect 193306 158378 193542 158614
rect 192986 158058 193222 158294
rect 193306 158058 193542 158294
rect 196706 234098 196942 234334
rect 197026 234098 197262 234334
rect 196706 233778 196942 234014
rect 197026 233778 197262 234014
rect 196706 198098 196942 198334
rect 197026 198098 197262 198334
rect 196706 197778 196942 198014
rect 197026 197778 197262 198014
rect 196706 162098 196942 162334
rect 197026 162098 197262 162334
rect 196706 161778 196942 162014
rect 197026 161778 197262 162014
rect 156986 122378 157222 122614
rect 157306 122378 157542 122614
rect 156986 122058 157222 122294
rect 157306 122058 157542 122294
rect 196706 126098 196942 126334
rect 197026 126098 197262 126334
rect 196706 125778 196942 126014
rect 197026 125778 197262 126014
rect 177610 114938 177846 115174
rect 177610 114618 177846 114854
rect 162250 111218 162486 111454
rect 162250 110898 162486 111134
rect 192970 111218 193206 111454
rect 192970 110898 193206 111134
rect 156986 86378 157222 86614
rect 157306 86378 157542 86614
rect 156986 86058 157222 86294
rect 157306 86058 157542 86294
rect 196706 90098 196942 90334
rect 197026 90098 197262 90334
rect 196706 89778 196942 90014
rect 197026 89778 197262 90014
rect 177610 78938 177846 79174
rect 177610 78618 177846 78854
rect 162250 75218 162486 75454
rect 162250 74898 162486 75134
rect 192970 75218 193206 75454
rect 192970 74898 193206 75134
rect 196706 54098 196942 54334
rect 197026 54098 197262 54334
rect 196706 53778 196942 54014
rect 197026 53778 197262 54014
rect 156986 50378 157222 50614
rect 157306 50378 157542 50614
rect 156986 50058 157222 50294
rect 157306 50058 157542 50294
rect 156986 14378 157222 14614
rect 157306 14378 157542 14614
rect 156986 14058 157222 14294
rect 157306 14058 157542 14294
rect 160706 18098 160942 18334
rect 161026 18098 161262 18334
rect 160706 17778 160942 18014
rect 161026 17778 161262 18014
rect 156986 -3462 157222 -3226
rect 157306 -3462 157542 -3226
rect 156986 -3782 157222 -3546
rect 157306 -3782 157542 -3546
rect 164426 21818 164662 22054
rect 164746 21818 164982 22054
rect 164426 21498 164662 21734
rect 164746 21498 164982 21734
rect 160706 -4422 160942 -4186
rect 161026 -4422 161262 -4186
rect 160706 -4742 160942 -4506
rect 161026 -4742 161262 -4506
rect 168146 25538 168382 25774
rect 168466 25538 168702 25774
rect 168146 25218 168382 25454
rect 168466 25218 168702 25454
rect 164426 -5382 164662 -5146
rect 164746 -5382 164982 -5146
rect 164426 -5702 164662 -5466
rect 164746 -5702 164982 -5466
rect 171866 29258 172102 29494
rect 172186 29258 172422 29494
rect 171866 28938 172102 29174
rect 172186 28938 172422 29174
rect 168146 -6342 168382 -6106
rect 168466 -6342 168702 -6106
rect 168146 -6662 168382 -6426
rect 168466 -6662 168702 -6426
rect 181826 39218 182062 39454
rect 182146 39218 182382 39454
rect 181826 38898 182062 39134
rect 182146 38898 182382 39134
rect 171866 -7302 172102 -7066
rect 172186 -7302 172422 -7066
rect 171866 -7622 172102 -7386
rect 172186 -7622 172422 -7386
rect 185546 42938 185782 43174
rect 185866 42938 186102 43174
rect 185546 42618 185782 42854
rect 185866 42618 186102 42854
rect 185546 6938 185782 7174
rect 185866 6938 186102 7174
rect 185546 6618 185782 6854
rect 185866 6618 186102 6854
rect 181826 3218 182062 3454
rect 182146 3218 182382 3454
rect 181826 2898 182062 3134
rect 182146 2898 182382 3134
rect 181826 -582 182062 -346
rect 182146 -582 182382 -346
rect 181826 -902 182062 -666
rect 182146 -902 182382 -666
rect 189266 46658 189502 46894
rect 189586 46658 189822 46894
rect 189266 46338 189502 46574
rect 189586 46338 189822 46574
rect 189266 10658 189502 10894
rect 189586 10658 189822 10894
rect 189266 10338 189502 10574
rect 189586 10338 189822 10574
rect 185546 -1542 185782 -1306
rect 185866 -1542 186102 -1306
rect 185546 -1862 185782 -1626
rect 185866 -1862 186102 -1626
rect 192986 50378 193222 50614
rect 193306 50378 193542 50614
rect 192986 50058 193222 50294
rect 193306 50058 193542 50294
rect 192986 14378 193222 14614
rect 193306 14378 193542 14614
rect 192986 14058 193222 14294
rect 193306 14058 193542 14294
rect 189266 -2502 189502 -2266
rect 189586 -2502 189822 -2266
rect 189266 -2822 189502 -2586
rect 189586 -2822 189822 -2586
rect 200426 237818 200662 238054
rect 200746 237818 200982 238054
rect 200426 237498 200662 237734
rect 200746 237498 200982 237734
rect 200426 201818 200662 202054
rect 200746 201818 200982 202054
rect 200426 201498 200662 201734
rect 200746 201498 200982 201734
rect 200426 165818 200662 166054
rect 200746 165818 200982 166054
rect 200426 165498 200662 165734
rect 200746 165498 200982 165734
rect 200426 129818 200662 130054
rect 200746 129818 200982 130054
rect 200426 129498 200662 129734
rect 200746 129498 200982 129734
rect 200426 93818 200662 94054
rect 200746 93818 200982 94054
rect 200426 93498 200662 93734
rect 200746 93498 200982 93734
rect 200426 57818 200662 58054
rect 200746 57818 200982 58054
rect 200426 57498 200662 57734
rect 200746 57498 200982 57734
rect 196706 18098 196942 18334
rect 197026 18098 197262 18334
rect 196706 17778 196942 18014
rect 197026 17778 197262 18014
rect 192986 -3462 193222 -3226
rect 193306 -3462 193542 -3226
rect 192986 -3782 193222 -3546
rect 193306 -3782 193542 -3546
rect 204146 241538 204382 241774
rect 204466 241538 204702 241774
rect 204146 241218 204382 241454
rect 204466 241218 204702 241454
rect 204146 205538 204382 205774
rect 204466 205538 204702 205774
rect 204146 205218 204382 205454
rect 204466 205218 204702 205454
rect 204146 169538 204382 169774
rect 204466 169538 204702 169774
rect 204146 169218 204382 169454
rect 204466 169218 204702 169454
rect 204146 133538 204382 133774
rect 204466 133538 204702 133774
rect 204146 133218 204382 133454
rect 204466 133218 204702 133454
rect 207866 245258 208102 245494
rect 208186 245258 208422 245494
rect 207866 244938 208102 245174
rect 208186 244938 208422 245174
rect 207866 209258 208102 209494
rect 208186 209258 208422 209494
rect 207866 208938 208102 209174
rect 208186 208938 208422 209174
rect 207866 173258 208102 173494
rect 208186 173258 208422 173494
rect 207866 172938 208102 173174
rect 208186 172938 208422 173174
rect 207866 137258 208102 137494
rect 208186 137258 208422 137494
rect 207866 136938 208102 137174
rect 208186 136938 208422 137174
rect 217826 255218 218062 255454
rect 218146 255218 218382 255454
rect 217826 254898 218062 255134
rect 218146 254898 218382 255134
rect 217826 219218 218062 219454
rect 218146 219218 218382 219454
rect 217826 218898 218062 219134
rect 218146 218898 218382 219134
rect 217826 183218 218062 183454
rect 218146 183218 218382 183454
rect 217826 182898 218062 183134
rect 218146 182898 218382 183134
rect 217826 147218 218062 147454
rect 218146 147218 218382 147454
rect 217826 146898 218062 147134
rect 218146 146898 218382 147134
rect 208330 114938 208566 115174
rect 208330 114618 208566 114854
rect 204146 97538 204382 97774
rect 204466 97538 204702 97774
rect 204146 97218 204382 97454
rect 204466 97218 204702 97454
rect 217826 111218 218062 111454
rect 218146 111218 218382 111454
rect 217826 110898 218062 111134
rect 218146 110898 218382 111134
rect 208330 78938 208566 79174
rect 208330 78618 208566 78854
rect 204146 61538 204382 61774
rect 204466 61538 204702 61774
rect 204146 61218 204382 61454
rect 204466 61218 204702 61454
rect 200426 21818 200662 22054
rect 200746 21818 200982 22054
rect 200426 21498 200662 21734
rect 200746 21498 200982 21734
rect 196706 -4422 196942 -4186
rect 197026 -4422 197262 -4186
rect 196706 -4742 196942 -4506
rect 197026 -4742 197262 -4506
rect 217826 75218 218062 75454
rect 218146 75218 218382 75454
rect 217826 74898 218062 75134
rect 218146 74898 218382 75134
rect 204146 25538 204382 25774
rect 204466 25538 204702 25774
rect 204146 25218 204382 25454
rect 204466 25218 204702 25454
rect 200426 -5382 200662 -5146
rect 200746 -5382 200982 -5146
rect 200426 -5702 200662 -5466
rect 200746 -5702 200982 -5466
rect 207866 29258 208102 29494
rect 208186 29258 208422 29494
rect 207866 28938 208102 29174
rect 208186 28938 208422 29174
rect 204146 -6342 204382 -6106
rect 204466 -6342 204702 -6106
rect 204146 -6662 204382 -6426
rect 204466 -6662 204702 -6426
rect 217826 39218 218062 39454
rect 218146 39218 218382 39454
rect 217826 38898 218062 39134
rect 218146 38898 218382 39134
rect 207866 -7302 208102 -7066
rect 208186 -7302 208422 -7066
rect 207866 -7622 208102 -7386
rect 208186 -7622 208422 -7386
rect 217826 3218 218062 3454
rect 218146 3218 218382 3454
rect 217826 2898 218062 3134
rect 218146 2898 218382 3134
rect 217826 -582 218062 -346
rect 218146 -582 218382 -346
rect 217826 -902 218062 -666
rect 218146 -902 218382 -666
rect 221546 705562 221782 705798
rect 221866 705562 222102 705798
rect 221546 705242 221782 705478
rect 221866 705242 222102 705478
rect 221546 690938 221782 691174
rect 221866 690938 222102 691174
rect 221546 690618 221782 690854
rect 221866 690618 222102 690854
rect 221546 654938 221782 655174
rect 221866 654938 222102 655174
rect 221546 654618 221782 654854
rect 221866 654618 222102 654854
rect 221546 618938 221782 619174
rect 221866 618938 222102 619174
rect 221546 618618 221782 618854
rect 221866 618618 222102 618854
rect 221546 582938 221782 583174
rect 221866 582938 222102 583174
rect 221546 582618 221782 582854
rect 221866 582618 222102 582854
rect 221546 546938 221782 547174
rect 221866 546938 222102 547174
rect 221546 546618 221782 546854
rect 221866 546618 222102 546854
rect 221546 510938 221782 511174
rect 221866 510938 222102 511174
rect 221546 510618 221782 510854
rect 221866 510618 222102 510854
rect 221546 474938 221782 475174
rect 221866 474938 222102 475174
rect 221546 474618 221782 474854
rect 221866 474618 222102 474854
rect 221546 438938 221782 439174
rect 221866 438938 222102 439174
rect 221546 438618 221782 438854
rect 221866 438618 222102 438854
rect 221546 402938 221782 403174
rect 221866 402938 222102 403174
rect 221546 402618 221782 402854
rect 221866 402618 222102 402854
rect 221546 366938 221782 367174
rect 221866 366938 222102 367174
rect 221546 366618 221782 366854
rect 221866 366618 222102 366854
rect 221546 330938 221782 331174
rect 221866 330938 222102 331174
rect 221546 330618 221782 330854
rect 221866 330618 222102 330854
rect 225266 706522 225502 706758
rect 225586 706522 225822 706758
rect 225266 706202 225502 706438
rect 225586 706202 225822 706438
rect 225266 694658 225502 694894
rect 225586 694658 225822 694894
rect 225266 694338 225502 694574
rect 225586 694338 225822 694574
rect 225266 658658 225502 658894
rect 225586 658658 225822 658894
rect 225266 658338 225502 658574
rect 225586 658338 225822 658574
rect 225266 622658 225502 622894
rect 225586 622658 225822 622894
rect 225266 622338 225502 622574
rect 225586 622338 225822 622574
rect 225266 586658 225502 586894
rect 225586 586658 225822 586894
rect 225266 586338 225502 586574
rect 225586 586338 225822 586574
rect 225266 550658 225502 550894
rect 225586 550658 225822 550894
rect 225266 550338 225502 550574
rect 225586 550338 225822 550574
rect 225266 514658 225502 514894
rect 225586 514658 225822 514894
rect 225266 514338 225502 514574
rect 225586 514338 225822 514574
rect 225266 478658 225502 478894
rect 225586 478658 225822 478894
rect 225266 478338 225502 478574
rect 225586 478338 225822 478574
rect 225266 442658 225502 442894
rect 225586 442658 225822 442894
rect 225266 442338 225502 442574
rect 225586 442338 225822 442574
rect 225266 406658 225502 406894
rect 225586 406658 225822 406894
rect 225266 406338 225502 406574
rect 225586 406338 225822 406574
rect 225266 370658 225502 370894
rect 225586 370658 225822 370894
rect 225266 370338 225502 370574
rect 225586 370338 225822 370574
rect 225266 334658 225502 334894
rect 225586 334658 225822 334894
rect 225266 334338 225502 334574
rect 225586 334338 225822 334574
rect 221546 294938 221782 295174
rect 221866 294938 222102 295174
rect 221546 294618 221782 294854
rect 221866 294618 222102 294854
rect 221546 258938 221782 259174
rect 221866 258938 222102 259174
rect 221546 258618 221782 258854
rect 221866 258618 222102 258854
rect 221546 222938 221782 223174
rect 221866 222938 222102 223174
rect 221546 222618 221782 222854
rect 221866 222618 222102 222854
rect 221546 186938 221782 187174
rect 221866 186938 222102 187174
rect 221546 186618 221782 186854
rect 221866 186618 222102 186854
rect 221546 150938 221782 151174
rect 221866 150938 222102 151174
rect 221546 150618 221782 150854
rect 221866 150618 222102 150854
rect 225266 298658 225502 298894
rect 225586 298658 225822 298894
rect 225266 298338 225502 298574
rect 225586 298338 225822 298574
rect 225266 262658 225502 262894
rect 225586 262658 225822 262894
rect 225266 262338 225502 262574
rect 225586 262338 225822 262574
rect 225266 226658 225502 226894
rect 225586 226658 225822 226894
rect 225266 226338 225502 226574
rect 225586 226338 225822 226574
rect 225266 190658 225502 190894
rect 225586 190658 225822 190894
rect 225266 190338 225502 190574
rect 225586 190338 225822 190574
rect 225266 154658 225502 154894
rect 225586 154658 225822 154894
rect 225266 154338 225502 154574
rect 225586 154338 225822 154574
rect 221546 114938 221782 115174
rect 221866 114938 222102 115174
rect 221546 114618 221782 114854
rect 221866 114618 222102 114854
rect 221546 78938 221782 79174
rect 221866 78938 222102 79174
rect 221546 78618 221782 78854
rect 221866 78618 222102 78854
rect 221546 42938 221782 43174
rect 221866 42938 222102 43174
rect 221546 42618 221782 42854
rect 221866 42618 222102 42854
rect 221546 6938 221782 7174
rect 221866 6938 222102 7174
rect 221546 6618 221782 6854
rect 221866 6618 222102 6854
rect 221546 -1542 221782 -1306
rect 221866 -1542 222102 -1306
rect 221546 -1862 221782 -1626
rect 221866 -1862 222102 -1626
rect 225266 118658 225502 118894
rect 225586 118658 225822 118894
rect 225266 118338 225502 118574
rect 225586 118338 225822 118574
rect 225266 82658 225502 82894
rect 225586 82658 225822 82894
rect 225266 82338 225502 82574
rect 225586 82338 225822 82574
rect 225266 46658 225502 46894
rect 225586 46658 225822 46894
rect 225266 46338 225502 46574
rect 225586 46338 225822 46574
rect 225266 10658 225502 10894
rect 225586 10658 225822 10894
rect 225266 10338 225502 10574
rect 225586 10338 225822 10574
rect 225266 -2502 225502 -2266
rect 225586 -2502 225822 -2266
rect 225266 -2822 225502 -2586
rect 225586 -2822 225822 -2586
rect 228986 707482 229222 707718
rect 229306 707482 229542 707718
rect 228986 707162 229222 707398
rect 229306 707162 229542 707398
rect 228986 698378 229222 698614
rect 229306 698378 229542 698614
rect 228986 698058 229222 698294
rect 229306 698058 229542 698294
rect 228986 662378 229222 662614
rect 229306 662378 229542 662614
rect 228986 662058 229222 662294
rect 229306 662058 229542 662294
rect 228986 626378 229222 626614
rect 229306 626378 229542 626614
rect 228986 626058 229222 626294
rect 229306 626058 229542 626294
rect 228986 590378 229222 590614
rect 229306 590378 229542 590614
rect 228986 590058 229222 590294
rect 229306 590058 229542 590294
rect 228986 554378 229222 554614
rect 229306 554378 229542 554614
rect 228986 554058 229222 554294
rect 229306 554058 229542 554294
rect 228986 518378 229222 518614
rect 229306 518378 229542 518614
rect 228986 518058 229222 518294
rect 229306 518058 229542 518294
rect 228986 482378 229222 482614
rect 229306 482378 229542 482614
rect 228986 482058 229222 482294
rect 229306 482058 229542 482294
rect 228986 446378 229222 446614
rect 229306 446378 229542 446614
rect 228986 446058 229222 446294
rect 229306 446058 229542 446294
rect 228986 410378 229222 410614
rect 229306 410378 229542 410614
rect 228986 410058 229222 410294
rect 229306 410058 229542 410294
rect 228986 374378 229222 374614
rect 229306 374378 229542 374614
rect 228986 374058 229222 374294
rect 229306 374058 229542 374294
rect 228986 338378 229222 338614
rect 229306 338378 229542 338614
rect 228986 338058 229222 338294
rect 229306 338058 229542 338294
rect 228986 302378 229222 302614
rect 229306 302378 229542 302614
rect 228986 302058 229222 302294
rect 229306 302058 229542 302294
rect 228986 266378 229222 266614
rect 229306 266378 229542 266614
rect 228986 266058 229222 266294
rect 229306 266058 229542 266294
rect 228986 230378 229222 230614
rect 229306 230378 229542 230614
rect 228986 230058 229222 230294
rect 229306 230058 229542 230294
rect 228986 194378 229222 194614
rect 229306 194378 229542 194614
rect 228986 194058 229222 194294
rect 229306 194058 229542 194294
rect 228986 158378 229222 158614
rect 229306 158378 229542 158614
rect 228986 158058 229222 158294
rect 229306 158058 229542 158294
rect 228986 122378 229222 122614
rect 229306 122378 229542 122614
rect 228986 122058 229222 122294
rect 229306 122058 229542 122294
rect 228986 86378 229222 86614
rect 229306 86378 229542 86614
rect 228986 86058 229222 86294
rect 229306 86058 229542 86294
rect 228986 50378 229222 50614
rect 229306 50378 229542 50614
rect 228986 50058 229222 50294
rect 229306 50058 229542 50294
rect 228986 14378 229222 14614
rect 229306 14378 229542 14614
rect 228986 14058 229222 14294
rect 229306 14058 229542 14294
rect 228986 -3462 229222 -3226
rect 229306 -3462 229542 -3226
rect 228986 -3782 229222 -3546
rect 229306 -3782 229542 -3546
rect 232706 708442 232942 708678
rect 233026 708442 233262 708678
rect 232706 708122 232942 708358
rect 233026 708122 233262 708358
rect 232706 666098 232942 666334
rect 233026 666098 233262 666334
rect 232706 665778 232942 666014
rect 233026 665778 233262 666014
rect 232706 630098 232942 630334
rect 233026 630098 233262 630334
rect 232706 629778 232942 630014
rect 233026 629778 233262 630014
rect 232706 594098 232942 594334
rect 233026 594098 233262 594334
rect 232706 593778 232942 594014
rect 233026 593778 233262 594014
rect 232706 558098 232942 558334
rect 233026 558098 233262 558334
rect 232706 557778 232942 558014
rect 233026 557778 233262 558014
rect 232706 522098 232942 522334
rect 233026 522098 233262 522334
rect 232706 521778 232942 522014
rect 233026 521778 233262 522014
rect 232706 486098 232942 486334
rect 233026 486098 233262 486334
rect 232706 485778 232942 486014
rect 233026 485778 233262 486014
rect 232706 450098 232942 450334
rect 233026 450098 233262 450334
rect 232706 449778 232942 450014
rect 233026 449778 233262 450014
rect 232706 414098 232942 414334
rect 233026 414098 233262 414334
rect 232706 413778 232942 414014
rect 233026 413778 233262 414014
rect 232706 378098 232942 378334
rect 233026 378098 233262 378334
rect 232706 377778 232942 378014
rect 233026 377778 233262 378014
rect 232706 342098 232942 342334
rect 233026 342098 233262 342334
rect 232706 341778 232942 342014
rect 233026 341778 233262 342014
rect 232706 306098 232942 306334
rect 233026 306098 233262 306334
rect 232706 305778 232942 306014
rect 233026 305778 233262 306014
rect 232706 270098 232942 270334
rect 233026 270098 233262 270334
rect 232706 269778 232942 270014
rect 233026 269778 233262 270014
rect 232706 234098 232942 234334
rect 233026 234098 233262 234334
rect 232706 233778 232942 234014
rect 233026 233778 233262 234014
rect 232706 198098 232942 198334
rect 233026 198098 233262 198334
rect 232706 197778 232942 198014
rect 233026 197778 233262 198014
rect 232706 162098 232942 162334
rect 233026 162098 233262 162334
rect 232706 161778 232942 162014
rect 233026 161778 233262 162014
rect 232706 126098 232942 126334
rect 233026 126098 233262 126334
rect 232706 125778 232942 126014
rect 233026 125778 233262 126014
rect 232706 90098 232942 90334
rect 233026 90098 233262 90334
rect 232706 89778 232942 90014
rect 233026 89778 233262 90014
rect 232706 54098 232942 54334
rect 233026 54098 233262 54334
rect 232706 53778 232942 54014
rect 233026 53778 233262 54014
rect 232706 18098 232942 18334
rect 233026 18098 233262 18334
rect 232706 17778 232942 18014
rect 233026 17778 233262 18014
rect 232706 -4422 232942 -4186
rect 233026 -4422 233262 -4186
rect 232706 -4742 232942 -4506
rect 233026 -4742 233262 -4506
rect 236426 709402 236662 709638
rect 236746 709402 236982 709638
rect 236426 709082 236662 709318
rect 236746 709082 236982 709318
rect 236426 669818 236662 670054
rect 236746 669818 236982 670054
rect 236426 669498 236662 669734
rect 236746 669498 236982 669734
rect 236426 633818 236662 634054
rect 236746 633818 236982 634054
rect 236426 633498 236662 633734
rect 236746 633498 236982 633734
rect 236426 597818 236662 598054
rect 236746 597818 236982 598054
rect 236426 597498 236662 597734
rect 236746 597498 236982 597734
rect 236426 561818 236662 562054
rect 236746 561818 236982 562054
rect 236426 561498 236662 561734
rect 236746 561498 236982 561734
rect 236426 525818 236662 526054
rect 236746 525818 236982 526054
rect 236426 525498 236662 525734
rect 236746 525498 236982 525734
rect 236426 489818 236662 490054
rect 236746 489818 236982 490054
rect 236426 489498 236662 489734
rect 236746 489498 236982 489734
rect 236426 453818 236662 454054
rect 236746 453818 236982 454054
rect 236426 453498 236662 453734
rect 236746 453498 236982 453734
rect 236426 417818 236662 418054
rect 236746 417818 236982 418054
rect 236426 417498 236662 417734
rect 236746 417498 236982 417734
rect 236426 381818 236662 382054
rect 236746 381818 236982 382054
rect 236426 381498 236662 381734
rect 236746 381498 236982 381734
rect 236426 345818 236662 346054
rect 236746 345818 236982 346054
rect 236426 345498 236662 345734
rect 236746 345498 236982 345734
rect 236426 309818 236662 310054
rect 236746 309818 236982 310054
rect 236426 309498 236662 309734
rect 236746 309498 236982 309734
rect 236426 273818 236662 274054
rect 236746 273818 236982 274054
rect 236426 273498 236662 273734
rect 236746 273498 236982 273734
rect 236426 237818 236662 238054
rect 236746 237818 236982 238054
rect 236426 237498 236662 237734
rect 236746 237498 236982 237734
rect 236426 201818 236662 202054
rect 236746 201818 236982 202054
rect 236426 201498 236662 201734
rect 236746 201498 236982 201734
rect 236426 165818 236662 166054
rect 236746 165818 236982 166054
rect 236426 165498 236662 165734
rect 236746 165498 236982 165734
rect 236426 129818 236662 130054
rect 236746 129818 236982 130054
rect 236426 129498 236662 129734
rect 236746 129498 236982 129734
rect 236426 93818 236662 94054
rect 236746 93818 236982 94054
rect 236426 93498 236662 93734
rect 236746 93498 236982 93734
rect 236426 57818 236662 58054
rect 236746 57818 236982 58054
rect 236426 57498 236662 57734
rect 236746 57498 236982 57734
rect 236426 21818 236662 22054
rect 236746 21818 236982 22054
rect 236426 21498 236662 21734
rect 236746 21498 236982 21734
rect 236426 -5382 236662 -5146
rect 236746 -5382 236982 -5146
rect 236426 -5702 236662 -5466
rect 236746 -5702 236982 -5466
rect 240146 710362 240382 710598
rect 240466 710362 240702 710598
rect 240146 710042 240382 710278
rect 240466 710042 240702 710278
rect 240146 673538 240382 673774
rect 240466 673538 240702 673774
rect 240146 673218 240382 673454
rect 240466 673218 240702 673454
rect 240146 637538 240382 637774
rect 240466 637538 240702 637774
rect 240146 637218 240382 637454
rect 240466 637218 240702 637454
rect 240146 601538 240382 601774
rect 240466 601538 240702 601774
rect 240146 601218 240382 601454
rect 240466 601218 240702 601454
rect 240146 565538 240382 565774
rect 240466 565538 240702 565774
rect 240146 565218 240382 565454
rect 240466 565218 240702 565454
rect 240146 529538 240382 529774
rect 240466 529538 240702 529774
rect 240146 529218 240382 529454
rect 240466 529218 240702 529454
rect 240146 493538 240382 493774
rect 240466 493538 240702 493774
rect 240146 493218 240382 493454
rect 240466 493218 240702 493454
rect 240146 457538 240382 457774
rect 240466 457538 240702 457774
rect 240146 457218 240382 457454
rect 240466 457218 240702 457454
rect 240146 421538 240382 421774
rect 240466 421538 240702 421774
rect 240146 421218 240382 421454
rect 240466 421218 240702 421454
rect 240146 385538 240382 385774
rect 240466 385538 240702 385774
rect 240146 385218 240382 385454
rect 240466 385218 240702 385454
rect 240146 349538 240382 349774
rect 240466 349538 240702 349774
rect 240146 349218 240382 349454
rect 240466 349218 240702 349454
rect 240146 313538 240382 313774
rect 240466 313538 240702 313774
rect 240146 313218 240382 313454
rect 240466 313218 240702 313454
rect 240146 277538 240382 277774
rect 240466 277538 240702 277774
rect 240146 277218 240382 277454
rect 240466 277218 240702 277454
rect 240146 241538 240382 241774
rect 240466 241538 240702 241774
rect 240146 241218 240382 241454
rect 240466 241218 240702 241454
rect 240146 205538 240382 205774
rect 240466 205538 240702 205774
rect 240146 205218 240382 205454
rect 240466 205218 240702 205454
rect 240146 169538 240382 169774
rect 240466 169538 240702 169774
rect 240146 169218 240382 169454
rect 240466 169218 240702 169454
rect 240146 133538 240382 133774
rect 240466 133538 240702 133774
rect 240146 133218 240382 133454
rect 240466 133218 240702 133454
rect 240146 97538 240382 97774
rect 240466 97538 240702 97774
rect 240146 97218 240382 97454
rect 240466 97218 240702 97454
rect 240146 61538 240382 61774
rect 240466 61538 240702 61774
rect 240146 61218 240382 61454
rect 240466 61218 240702 61454
rect 240146 25538 240382 25774
rect 240466 25538 240702 25774
rect 240146 25218 240382 25454
rect 240466 25218 240702 25454
rect 240146 -6342 240382 -6106
rect 240466 -6342 240702 -6106
rect 240146 -6662 240382 -6426
rect 240466 -6662 240702 -6426
rect 243866 711322 244102 711558
rect 244186 711322 244422 711558
rect 243866 711002 244102 711238
rect 244186 711002 244422 711238
rect 243866 677258 244102 677494
rect 244186 677258 244422 677494
rect 243866 676938 244102 677174
rect 244186 676938 244422 677174
rect 253826 704602 254062 704838
rect 254146 704602 254382 704838
rect 253826 704282 254062 704518
rect 254146 704282 254382 704518
rect 253826 687218 254062 687454
rect 254146 687218 254382 687454
rect 253826 686898 254062 687134
rect 254146 686898 254382 687134
rect 243866 641258 244102 641494
rect 244186 641258 244422 641494
rect 243866 640938 244102 641174
rect 244186 640938 244422 641174
rect 243866 605258 244102 605494
rect 244186 605258 244422 605494
rect 243866 604938 244102 605174
rect 244186 604938 244422 605174
rect 243866 569258 244102 569494
rect 244186 569258 244422 569494
rect 243866 568938 244102 569174
rect 244186 568938 244422 569174
rect 243866 533258 244102 533494
rect 244186 533258 244422 533494
rect 243866 532938 244102 533174
rect 244186 532938 244422 533174
rect 243866 497258 244102 497494
rect 244186 497258 244422 497494
rect 243866 496938 244102 497174
rect 244186 496938 244422 497174
rect 243866 461258 244102 461494
rect 244186 461258 244422 461494
rect 243866 460938 244102 461174
rect 244186 460938 244422 461174
rect 243866 425258 244102 425494
rect 244186 425258 244422 425494
rect 243866 424938 244102 425174
rect 244186 424938 244422 425174
rect 243866 389258 244102 389494
rect 244186 389258 244422 389494
rect 243866 388938 244102 389174
rect 244186 388938 244422 389174
rect 243866 353258 244102 353494
rect 244186 353258 244422 353494
rect 243866 352938 244102 353174
rect 244186 352938 244422 353174
rect 243866 317258 244102 317494
rect 244186 317258 244422 317494
rect 243866 316938 244102 317174
rect 244186 316938 244422 317174
rect 243866 281258 244102 281494
rect 244186 281258 244422 281494
rect 243866 280938 244102 281174
rect 244186 280938 244422 281174
rect 243866 245258 244102 245494
rect 244186 245258 244422 245494
rect 243866 244938 244102 245174
rect 244186 244938 244422 245174
rect 243866 209258 244102 209494
rect 244186 209258 244422 209494
rect 243866 208938 244102 209174
rect 244186 208938 244422 209174
rect 243866 173258 244102 173494
rect 244186 173258 244422 173494
rect 243866 172938 244102 173174
rect 244186 172938 244422 173174
rect 243866 137258 244102 137494
rect 244186 137258 244422 137494
rect 243866 136938 244102 137174
rect 244186 136938 244422 137174
rect 243866 101258 244102 101494
rect 244186 101258 244422 101494
rect 243866 100938 244102 101174
rect 244186 100938 244422 101174
rect 243866 65258 244102 65494
rect 244186 65258 244422 65494
rect 243866 64938 244102 65174
rect 244186 64938 244422 65174
rect 253826 651218 254062 651454
rect 254146 651218 254382 651454
rect 253826 650898 254062 651134
rect 254146 650898 254382 651134
rect 257546 705562 257782 705798
rect 257866 705562 258102 705798
rect 257546 705242 257782 705478
rect 257866 705242 258102 705478
rect 257546 690938 257782 691174
rect 257866 690938 258102 691174
rect 257546 690618 257782 690854
rect 257866 690618 258102 690854
rect 257546 654938 257782 655174
rect 257866 654938 258102 655174
rect 257546 654618 257782 654854
rect 257866 654618 258102 654854
rect 261266 706522 261502 706758
rect 261586 706522 261822 706758
rect 261266 706202 261502 706438
rect 261586 706202 261822 706438
rect 261266 694658 261502 694894
rect 261586 694658 261822 694894
rect 261266 694338 261502 694574
rect 261586 694338 261822 694574
rect 261266 658658 261502 658894
rect 261586 658658 261822 658894
rect 261266 658338 261502 658574
rect 261586 658338 261822 658574
rect 264986 707482 265222 707718
rect 265306 707482 265542 707718
rect 264986 707162 265222 707398
rect 265306 707162 265542 707398
rect 264986 698378 265222 698614
rect 265306 698378 265542 698614
rect 264986 698058 265222 698294
rect 265306 698058 265542 698294
rect 264986 662378 265222 662614
rect 265306 662378 265542 662614
rect 264986 662058 265222 662294
rect 265306 662058 265542 662294
rect 268706 708442 268942 708678
rect 269026 708442 269262 708678
rect 268706 708122 268942 708358
rect 269026 708122 269262 708358
rect 268706 666098 268942 666334
rect 269026 666098 269262 666334
rect 268706 665778 268942 666014
rect 269026 665778 269262 666014
rect 272426 709402 272662 709638
rect 272746 709402 272982 709638
rect 272426 709082 272662 709318
rect 272746 709082 272982 709318
rect 272426 669818 272662 670054
rect 272746 669818 272982 670054
rect 272426 669498 272662 669734
rect 272746 669498 272982 669734
rect 276146 710362 276382 710598
rect 276466 710362 276702 710598
rect 276146 710042 276382 710278
rect 276466 710042 276702 710278
rect 276146 673538 276382 673774
rect 276466 673538 276702 673774
rect 276146 673218 276382 673454
rect 276466 673218 276702 673454
rect 279866 711322 280102 711558
rect 280186 711322 280422 711558
rect 279866 711002 280102 711238
rect 280186 711002 280422 711238
rect 279866 677258 280102 677494
rect 280186 677258 280422 677494
rect 279866 676938 280102 677174
rect 280186 676938 280422 677174
rect 289826 704602 290062 704838
rect 290146 704602 290382 704838
rect 289826 704282 290062 704518
rect 290146 704282 290382 704518
rect 289826 687218 290062 687454
rect 290146 687218 290382 687454
rect 289826 686898 290062 687134
rect 290146 686898 290382 687134
rect 289826 651218 290062 651454
rect 290146 651218 290382 651454
rect 289826 650898 290062 651134
rect 290146 650898 290382 651134
rect 293546 705562 293782 705798
rect 293866 705562 294102 705798
rect 293546 705242 293782 705478
rect 293866 705242 294102 705478
rect 293546 690938 293782 691174
rect 293866 690938 294102 691174
rect 293546 690618 293782 690854
rect 293866 690618 294102 690854
rect 293546 654938 293782 655174
rect 293866 654938 294102 655174
rect 293546 654618 293782 654854
rect 293866 654618 294102 654854
rect 297266 706522 297502 706758
rect 297586 706522 297822 706758
rect 297266 706202 297502 706438
rect 297586 706202 297822 706438
rect 297266 694658 297502 694894
rect 297586 694658 297822 694894
rect 297266 694338 297502 694574
rect 297586 694338 297822 694574
rect 297266 658658 297502 658894
rect 297586 658658 297822 658894
rect 297266 658338 297502 658574
rect 297586 658338 297822 658574
rect 300986 707482 301222 707718
rect 301306 707482 301542 707718
rect 300986 707162 301222 707398
rect 301306 707162 301542 707398
rect 300986 698378 301222 698614
rect 301306 698378 301542 698614
rect 300986 698058 301222 698294
rect 301306 698058 301542 698294
rect 300986 662378 301222 662614
rect 301306 662378 301542 662614
rect 300986 662058 301222 662294
rect 301306 662058 301542 662294
rect 304706 708442 304942 708678
rect 305026 708442 305262 708678
rect 304706 708122 304942 708358
rect 305026 708122 305262 708358
rect 304706 666098 304942 666334
rect 305026 666098 305262 666334
rect 304706 665778 304942 666014
rect 305026 665778 305262 666014
rect 308426 709402 308662 709638
rect 308746 709402 308982 709638
rect 308426 709082 308662 709318
rect 308746 709082 308982 709318
rect 308426 669818 308662 670054
rect 308746 669818 308982 670054
rect 308426 669498 308662 669734
rect 308746 669498 308982 669734
rect 312146 710362 312382 710598
rect 312466 710362 312702 710598
rect 312146 710042 312382 710278
rect 312466 710042 312702 710278
rect 312146 673538 312382 673774
rect 312466 673538 312702 673774
rect 312146 673218 312382 673454
rect 312466 673218 312702 673454
rect 315866 711322 316102 711558
rect 316186 711322 316422 711558
rect 315866 711002 316102 711238
rect 316186 711002 316422 711238
rect 315866 677258 316102 677494
rect 316186 677258 316422 677494
rect 315866 676938 316102 677174
rect 316186 676938 316422 677174
rect 325826 704602 326062 704838
rect 326146 704602 326382 704838
rect 325826 704282 326062 704518
rect 326146 704282 326382 704518
rect 325826 687218 326062 687454
rect 326146 687218 326382 687454
rect 325826 686898 326062 687134
rect 326146 686898 326382 687134
rect 325826 651218 326062 651454
rect 326146 651218 326382 651454
rect 325826 650898 326062 651134
rect 326146 650898 326382 651134
rect 329546 705562 329782 705798
rect 329866 705562 330102 705798
rect 329546 705242 329782 705478
rect 329866 705242 330102 705478
rect 329546 690938 329782 691174
rect 329866 690938 330102 691174
rect 329546 690618 329782 690854
rect 329866 690618 330102 690854
rect 329546 654938 329782 655174
rect 329866 654938 330102 655174
rect 329546 654618 329782 654854
rect 329866 654618 330102 654854
rect 333266 706522 333502 706758
rect 333586 706522 333822 706758
rect 333266 706202 333502 706438
rect 333586 706202 333822 706438
rect 333266 694658 333502 694894
rect 333586 694658 333822 694894
rect 333266 694338 333502 694574
rect 333586 694338 333822 694574
rect 333266 658658 333502 658894
rect 333586 658658 333822 658894
rect 333266 658338 333502 658574
rect 333586 658338 333822 658574
rect 336986 707482 337222 707718
rect 337306 707482 337542 707718
rect 336986 707162 337222 707398
rect 337306 707162 337542 707398
rect 336986 698378 337222 698614
rect 337306 698378 337542 698614
rect 336986 698058 337222 698294
rect 337306 698058 337542 698294
rect 336986 662378 337222 662614
rect 337306 662378 337542 662614
rect 336986 662058 337222 662294
rect 337306 662058 337542 662294
rect 340706 708442 340942 708678
rect 341026 708442 341262 708678
rect 340706 708122 340942 708358
rect 341026 708122 341262 708358
rect 340706 666098 340942 666334
rect 341026 666098 341262 666334
rect 340706 665778 340942 666014
rect 341026 665778 341262 666014
rect 344426 709402 344662 709638
rect 344746 709402 344982 709638
rect 344426 709082 344662 709318
rect 344746 709082 344982 709318
rect 344426 669818 344662 670054
rect 344746 669818 344982 670054
rect 344426 669498 344662 669734
rect 344746 669498 344982 669734
rect 348146 710362 348382 710598
rect 348466 710362 348702 710598
rect 348146 710042 348382 710278
rect 348466 710042 348702 710278
rect 348146 673538 348382 673774
rect 348466 673538 348702 673774
rect 348146 673218 348382 673454
rect 348466 673218 348702 673454
rect 351866 711322 352102 711558
rect 352186 711322 352422 711558
rect 351866 711002 352102 711238
rect 352186 711002 352422 711238
rect 351866 677258 352102 677494
rect 352186 677258 352422 677494
rect 351866 676938 352102 677174
rect 352186 676938 352422 677174
rect 361826 704602 362062 704838
rect 362146 704602 362382 704838
rect 361826 704282 362062 704518
rect 362146 704282 362382 704518
rect 361826 687218 362062 687454
rect 362146 687218 362382 687454
rect 361826 686898 362062 687134
rect 362146 686898 362382 687134
rect 361826 651218 362062 651454
rect 362146 651218 362382 651454
rect 361826 650898 362062 651134
rect 362146 650898 362382 651134
rect 365546 705562 365782 705798
rect 365866 705562 366102 705798
rect 365546 705242 365782 705478
rect 365866 705242 366102 705478
rect 365546 690938 365782 691174
rect 365866 690938 366102 691174
rect 365546 690618 365782 690854
rect 365866 690618 366102 690854
rect 365546 654938 365782 655174
rect 365866 654938 366102 655174
rect 365546 654618 365782 654854
rect 365866 654618 366102 654854
rect 369266 706522 369502 706758
rect 369586 706522 369822 706758
rect 369266 706202 369502 706438
rect 369586 706202 369822 706438
rect 369266 694658 369502 694894
rect 369586 694658 369822 694894
rect 369266 694338 369502 694574
rect 369586 694338 369822 694574
rect 369266 658658 369502 658894
rect 369586 658658 369822 658894
rect 369266 658338 369502 658574
rect 369586 658338 369822 658574
rect 372986 707482 373222 707718
rect 373306 707482 373542 707718
rect 372986 707162 373222 707398
rect 373306 707162 373542 707398
rect 372986 698378 373222 698614
rect 373306 698378 373542 698614
rect 372986 698058 373222 698294
rect 373306 698058 373542 698294
rect 372986 662378 373222 662614
rect 373306 662378 373542 662614
rect 372986 662058 373222 662294
rect 373306 662058 373542 662294
rect 376706 708442 376942 708678
rect 377026 708442 377262 708678
rect 376706 708122 376942 708358
rect 377026 708122 377262 708358
rect 376706 666098 376942 666334
rect 377026 666098 377262 666334
rect 376706 665778 376942 666014
rect 377026 665778 377262 666014
rect 380426 709402 380662 709638
rect 380746 709402 380982 709638
rect 380426 709082 380662 709318
rect 380746 709082 380982 709318
rect 380426 669818 380662 670054
rect 380746 669818 380982 670054
rect 380426 669498 380662 669734
rect 380746 669498 380982 669734
rect 384146 710362 384382 710598
rect 384466 710362 384702 710598
rect 384146 710042 384382 710278
rect 384466 710042 384702 710278
rect 384146 673538 384382 673774
rect 384466 673538 384702 673774
rect 384146 673218 384382 673454
rect 384466 673218 384702 673454
rect 387866 711322 388102 711558
rect 388186 711322 388422 711558
rect 387866 711002 388102 711238
rect 388186 711002 388422 711238
rect 387866 677258 388102 677494
rect 388186 677258 388422 677494
rect 387866 676938 388102 677174
rect 388186 676938 388422 677174
rect 397826 704602 398062 704838
rect 398146 704602 398382 704838
rect 397826 704282 398062 704518
rect 398146 704282 398382 704518
rect 397826 687218 398062 687454
rect 398146 687218 398382 687454
rect 397826 686898 398062 687134
rect 398146 686898 398382 687134
rect 397826 651218 398062 651454
rect 398146 651218 398382 651454
rect 397826 650898 398062 651134
rect 398146 650898 398382 651134
rect 401546 705562 401782 705798
rect 401866 705562 402102 705798
rect 401546 705242 401782 705478
rect 401866 705242 402102 705478
rect 401546 690938 401782 691174
rect 401866 690938 402102 691174
rect 401546 690618 401782 690854
rect 401866 690618 402102 690854
rect 401546 654938 401782 655174
rect 401866 654938 402102 655174
rect 401546 654618 401782 654854
rect 401866 654618 402102 654854
rect 405266 706522 405502 706758
rect 405586 706522 405822 706758
rect 405266 706202 405502 706438
rect 405586 706202 405822 706438
rect 405266 694658 405502 694894
rect 405586 694658 405822 694894
rect 405266 694338 405502 694574
rect 405586 694338 405822 694574
rect 405266 658658 405502 658894
rect 405586 658658 405822 658894
rect 405266 658338 405502 658574
rect 405586 658338 405822 658574
rect 408986 707482 409222 707718
rect 409306 707482 409542 707718
rect 408986 707162 409222 707398
rect 409306 707162 409542 707398
rect 408986 698378 409222 698614
rect 409306 698378 409542 698614
rect 408986 698058 409222 698294
rect 409306 698058 409542 698294
rect 408986 662378 409222 662614
rect 409306 662378 409542 662614
rect 408986 662058 409222 662294
rect 409306 662058 409542 662294
rect 412706 708442 412942 708678
rect 413026 708442 413262 708678
rect 412706 708122 412942 708358
rect 413026 708122 413262 708358
rect 412706 666098 412942 666334
rect 413026 666098 413262 666334
rect 412706 665778 412942 666014
rect 413026 665778 413262 666014
rect 416426 709402 416662 709638
rect 416746 709402 416982 709638
rect 416426 709082 416662 709318
rect 416746 709082 416982 709318
rect 416426 669818 416662 670054
rect 416746 669818 416982 670054
rect 416426 669498 416662 669734
rect 416746 669498 416982 669734
rect 420146 710362 420382 710598
rect 420466 710362 420702 710598
rect 420146 710042 420382 710278
rect 420466 710042 420702 710278
rect 420146 673538 420382 673774
rect 420466 673538 420702 673774
rect 420146 673218 420382 673454
rect 420466 673218 420702 673454
rect 423866 711322 424102 711558
rect 424186 711322 424422 711558
rect 423866 711002 424102 711238
rect 424186 711002 424422 711238
rect 423866 677258 424102 677494
rect 424186 677258 424422 677494
rect 423866 676938 424102 677174
rect 424186 676938 424422 677174
rect 433826 704602 434062 704838
rect 434146 704602 434382 704838
rect 433826 704282 434062 704518
rect 434146 704282 434382 704518
rect 433826 687218 434062 687454
rect 434146 687218 434382 687454
rect 433826 686898 434062 687134
rect 434146 686898 434382 687134
rect 433826 651218 434062 651454
rect 434146 651218 434382 651454
rect 433826 650898 434062 651134
rect 434146 650898 434382 651134
rect 437546 705562 437782 705798
rect 437866 705562 438102 705798
rect 437546 705242 437782 705478
rect 437866 705242 438102 705478
rect 437546 690938 437782 691174
rect 437866 690938 438102 691174
rect 437546 690618 437782 690854
rect 437866 690618 438102 690854
rect 437546 654938 437782 655174
rect 437866 654938 438102 655174
rect 437546 654618 437782 654854
rect 437866 654618 438102 654854
rect 441266 706522 441502 706758
rect 441586 706522 441822 706758
rect 441266 706202 441502 706438
rect 441586 706202 441822 706438
rect 441266 694658 441502 694894
rect 441586 694658 441822 694894
rect 441266 694338 441502 694574
rect 441586 694338 441822 694574
rect 441266 658658 441502 658894
rect 441586 658658 441822 658894
rect 441266 658338 441502 658574
rect 441586 658338 441822 658574
rect 444986 707482 445222 707718
rect 445306 707482 445542 707718
rect 444986 707162 445222 707398
rect 445306 707162 445542 707398
rect 444986 698378 445222 698614
rect 445306 698378 445542 698614
rect 444986 698058 445222 698294
rect 445306 698058 445542 698294
rect 444986 662378 445222 662614
rect 445306 662378 445542 662614
rect 444986 662058 445222 662294
rect 445306 662058 445542 662294
rect 448706 708442 448942 708678
rect 449026 708442 449262 708678
rect 448706 708122 448942 708358
rect 449026 708122 449262 708358
rect 448706 666098 448942 666334
rect 449026 666098 449262 666334
rect 448706 665778 448942 666014
rect 449026 665778 449262 666014
rect 452426 709402 452662 709638
rect 452746 709402 452982 709638
rect 452426 709082 452662 709318
rect 452746 709082 452982 709318
rect 452426 669818 452662 670054
rect 452746 669818 452982 670054
rect 452426 669498 452662 669734
rect 452746 669498 452982 669734
rect 456146 710362 456382 710598
rect 456466 710362 456702 710598
rect 456146 710042 456382 710278
rect 456466 710042 456702 710278
rect 456146 673538 456382 673774
rect 456466 673538 456702 673774
rect 456146 673218 456382 673454
rect 456466 673218 456702 673454
rect 459866 711322 460102 711558
rect 460186 711322 460422 711558
rect 459866 711002 460102 711238
rect 460186 711002 460422 711238
rect 459866 677258 460102 677494
rect 460186 677258 460422 677494
rect 459866 676938 460102 677174
rect 460186 676938 460422 677174
rect 469826 704602 470062 704838
rect 470146 704602 470382 704838
rect 469826 704282 470062 704518
rect 470146 704282 470382 704518
rect 469826 687218 470062 687454
rect 470146 687218 470382 687454
rect 469826 686898 470062 687134
rect 470146 686898 470382 687134
rect 469826 651218 470062 651454
rect 470146 651218 470382 651454
rect 469826 650898 470062 651134
rect 470146 650898 470382 651134
rect 473546 705562 473782 705798
rect 473866 705562 474102 705798
rect 473546 705242 473782 705478
rect 473866 705242 474102 705478
rect 473546 690938 473782 691174
rect 473866 690938 474102 691174
rect 473546 690618 473782 690854
rect 473866 690618 474102 690854
rect 473546 654938 473782 655174
rect 473866 654938 474102 655174
rect 473546 654618 473782 654854
rect 473866 654618 474102 654854
rect 477266 706522 477502 706758
rect 477586 706522 477822 706758
rect 477266 706202 477502 706438
rect 477586 706202 477822 706438
rect 477266 694658 477502 694894
rect 477586 694658 477822 694894
rect 477266 694338 477502 694574
rect 477586 694338 477822 694574
rect 477266 658658 477502 658894
rect 477586 658658 477822 658894
rect 477266 658338 477502 658574
rect 477586 658338 477822 658574
rect 480986 707482 481222 707718
rect 481306 707482 481542 707718
rect 480986 707162 481222 707398
rect 481306 707162 481542 707398
rect 480986 698378 481222 698614
rect 481306 698378 481542 698614
rect 480986 698058 481222 698294
rect 481306 698058 481542 698294
rect 480986 662378 481222 662614
rect 481306 662378 481542 662614
rect 480986 662058 481222 662294
rect 481306 662058 481542 662294
rect 484706 708442 484942 708678
rect 485026 708442 485262 708678
rect 484706 708122 484942 708358
rect 485026 708122 485262 708358
rect 484706 666098 484942 666334
rect 485026 666098 485262 666334
rect 484706 665778 484942 666014
rect 485026 665778 485262 666014
rect 488426 709402 488662 709638
rect 488746 709402 488982 709638
rect 488426 709082 488662 709318
rect 488746 709082 488982 709318
rect 488426 669818 488662 670054
rect 488746 669818 488982 670054
rect 488426 669498 488662 669734
rect 488746 669498 488982 669734
rect 492146 710362 492382 710598
rect 492466 710362 492702 710598
rect 492146 710042 492382 710278
rect 492466 710042 492702 710278
rect 492146 673538 492382 673774
rect 492466 673538 492702 673774
rect 492146 673218 492382 673454
rect 492466 673218 492702 673454
rect 495866 711322 496102 711558
rect 496186 711322 496422 711558
rect 495866 711002 496102 711238
rect 496186 711002 496422 711238
rect 495866 677258 496102 677494
rect 496186 677258 496422 677494
rect 495866 676938 496102 677174
rect 496186 676938 496422 677174
rect 505826 704602 506062 704838
rect 506146 704602 506382 704838
rect 505826 704282 506062 704518
rect 506146 704282 506382 704518
rect 505826 687218 506062 687454
rect 506146 687218 506382 687454
rect 505826 686898 506062 687134
rect 506146 686898 506382 687134
rect 505826 651218 506062 651454
rect 506146 651218 506382 651454
rect 505826 650898 506062 651134
rect 506146 650898 506382 651134
rect 509546 705562 509782 705798
rect 509866 705562 510102 705798
rect 509546 705242 509782 705478
rect 509866 705242 510102 705478
rect 509546 690938 509782 691174
rect 509866 690938 510102 691174
rect 509546 690618 509782 690854
rect 509866 690618 510102 690854
rect 509546 654938 509782 655174
rect 509866 654938 510102 655174
rect 509546 654618 509782 654854
rect 509866 654618 510102 654854
rect 513266 706522 513502 706758
rect 513586 706522 513822 706758
rect 513266 706202 513502 706438
rect 513586 706202 513822 706438
rect 513266 694658 513502 694894
rect 513586 694658 513822 694894
rect 513266 694338 513502 694574
rect 513586 694338 513822 694574
rect 513266 658658 513502 658894
rect 513586 658658 513822 658894
rect 513266 658338 513502 658574
rect 513586 658338 513822 658574
rect 516986 707482 517222 707718
rect 517306 707482 517542 707718
rect 516986 707162 517222 707398
rect 517306 707162 517542 707398
rect 516986 698378 517222 698614
rect 517306 698378 517542 698614
rect 516986 698058 517222 698294
rect 517306 698058 517542 698294
rect 516986 662378 517222 662614
rect 517306 662378 517542 662614
rect 516986 662058 517222 662294
rect 517306 662058 517542 662294
rect 520706 708442 520942 708678
rect 521026 708442 521262 708678
rect 520706 708122 520942 708358
rect 521026 708122 521262 708358
rect 520706 666098 520942 666334
rect 521026 666098 521262 666334
rect 520706 665778 520942 666014
rect 521026 665778 521262 666014
rect 524426 709402 524662 709638
rect 524746 709402 524982 709638
rect 524426 709082 524662 709318
rect 524746 709082 524982 709318
rect 524426 669818 524662 670054
rect 524746 669818 524982 670054
rect 524426 669498 524662 669734
rect 524746 669498 524982 669734
rect 528146 710362 528382 710598
rect 528466 710362 528702 710598
rect 528146 710042 528382 710278
rect 528466 710042 528702 710278
rect 528146 673538 528382 673774
rect 528466 673538 528702 673774
rect 528146 673218 528382 673454
rect 528466 673218 528702 673454
rect 531866 711322 532102 711558
rect 532186 711322 532422 711558
rect 531866 711002 532102 711238
rect 532186 711002 532422 711238
rect 531866 677258 532102 677494
rect 532186 677258 532422 677494
rect 531866 676938 532102 677174
rect 532186 676938 532422 677174
rect 541826 704602 542062 704838
rect 542146 704602 542382 704838
rect 541826 704282 542062 704518
rect 542146 704282 542382 704518
rect 541826 687218 542062 687454
rect 542146 687218 542382 687454
rect 541826 686898 542062 687134
rect 542146 686898 542382 687134
rect 541826 651218 542062 651454
rect 542146 651218 542382 651454
rect 541826 650898 542062 651134
rect 542146 650898 542382 651134
rect 273210 618938 273446 619174
rect 273210 618618 273446 618854
rect 303930 618938 304166 619174
rect 303930 618618 304166 618854
rect 334650 618938 334886 619174
rect 334650 618618 334886 618854
rect 365370 618938 365606 619174
rect 365370 618618 365606 618854
rect 396090 618938 396326 619174
rect 396090 618618 396326 618854
rect 426810 618938 427046 619174
rect 426810 618618 427046 618854
rect 457530 618938 457766 619174
rect 457530 618618 457766 618854
rect 488250 618938 488486 619174
rect 488250 618618 488486 618854
rect 518970 618938 519206 619174
rect 518970 618618 519206 618854
rect 253826 615218 254062 615454
rect 254146 615218 254382 615454
rect 253826 614898 254062 615134
rect 254146 614898 254382 615134
rect 257850 615218 258086 615454
rect 257850 614898 258086 615134
rect 288570 615218 288806 615454
rect 288570 614898 288806 615134
rect 319290 615218 319526 615454
rect 319290 614898 319526 615134
rect 350010 615218 350246 615454
rect 350010 614898 350246 615134
rect 380730 615218 380966 615454
rect 380730 614898 380966 615134
rect 411450 615218 411686 615454
rect 411450 614898 411686 615134
rect 442170 615218 442406 615454
rect 442170 614898 442406 615134
rect 472890 615218 473126 615454
rect 472890 614898 473126 615134
rect 503610 615218 503846 615454
rect 503610 614898 503846 615134
rect 534330 615218 534566 615454
rect 534330 614898 534566 615134
rect 541826 615218 542062 615454
rect 542146 615218 542382 615454
rect 541826 614898 542062 615134
rect 542146 614898 542382 615134
rect 273210 582938 273446 583174
rect 273210 582618 273446 582854
rect 303930 582938 304166 583174
rect 303930 582618 304166 582854
rect 334650 582938 334886 583174
rect 334650 582618 334886 582854
rect 365370 582938 365606 583174
rect 365370 582618 365606 582854
rect 396090 582938 396326 583174
rect 396090 582618 396326 582854
rect 426810 582938 427046 583174
rect 426810 582618 427046 582854
rect 457530 582938 457766 583174
rect 457530 582618 457766 582854
rect 488250 582938 488486 583174
rect 488250 582618 488486 582854
rect 518970 582938 519206 583174
rect 518970 582618 519206 582854
rect 253826 579218 254062 579454
rect 254146 579218 254382 579454
rect 253826 578898 254062 579134
rect 254146 578898 254382 579134
rect 257850 579218 258086 579454
rect 257850 578898 258086 579134
rect 288570 579218 288806 579454
rect 288570 578898 288806 579134
rect 319290 579218 319526 579454
rect 319290 578898 319526 579134
rect 350010 579218 350246 579454
rect 350010 578898 350246 579134
rect 380730 579218 380966 579454
rect 380730 578898 380966 579134
rect 411450 579218 411686 579454
rect 411450 578898 411686 579134
rect 442170 579218 442406 579454
rect 442170 578898 442406 579134
rect 472890 579218 473126 579454
rect 472890 578898 473126 579134
rect 503610 579218 503846 579454
rect 503610 578898 503846 579134
rect 534330 579218 534566 579454
rect 534330 578898 534566 579134
rect 541826 579218 542062 579454
rect 542146 579218 542382 579454
rect 541826 578898 542062 579134
rect 542146 578898 542382 579134
rect 273210 546938 273446 547174
rect 273210 546618 273446 546854
rect 303930 546938 304166 547174
rect 303930 546618 304166 546854
rect 334650 546938 334886 547174
rect 334650 546618 334886 546854
rect 365370 546938 365606 547174
rect 365370 546618 365606 546854
rect 396090 546938 396326 547174
rect 396090 546618 396326 546854
rect 426810 546938 427046 547174
rect 426810 546618 427046 546854
rect 457530 546938 457766 547174
rect 457530 546618 457766 546854
rect 488250 546938 488486 547174
rect 488250 546618 488486 546854
rect 518970 546938 519206 547174
rect 518970 546618 519206 546854
rect 253826 543218 254062 543454
rect 254146 543218 254382 543454
rect 253826 542898 254062 543134
rect 254146 542898 254382 543134
rect 257850 543218 258086 543454
rect 257850 542898 258086 543134
rect 288570 543218 288806 543454
rect 288570 542898 288806 543134
rect 319290 543218 319526 543454
rect 319290 542898 319526 543134
rect 350010 543218 350246 543454
rect 350010 542898 350246 543134
rect 380730 543218 380966 543454
rect 380730 542898 380966 543134
rect 411450 543218 411686 543454
rect 411450 542898 411686 543134
rect 442170 543218 442406 543454
rect 442170 542898 442406 543134
rect 472890 543218 473126 543454
rect 472890 542898 473126 543134
rect 503610 543218 503846 543454
rect 503610 542898 503846 543134
rect 534330 543218 534566 543454
rect 534330 542898 534566 543134
rect 541826 543218 542062 543454
rect 542146 543218 542382 543454
rect 541826 542898 542062 543134
rect 542146 542898 542382 543134
rect 253826 507218 254062 507454
rect 254146 507218 254382 507454
rect 253826 506898 254062 507134
rect 254146 506898 254382 507134
rect 276146 529538 276382 529774
rect 276466 529538 276702 529774
rect 276146 529218 276382 529454
rect 276466 529218 276702 529454
rect 312146 529538 312382 529774
rect 312466 529538 312702 529774
rect 312146 529218 312382 529454
rect 312466 529218 312702 529454
rect 348146 529538 348382 529774
rect 348466 529538 348702 529774
rect 348146 529218 348382 529454
rect 348466 529218 348702 529454
rect 384146 529538 384382 529774
rect 384466 529538 384702 529774
rect 384146 529218 384382 529454
rect 384466 529218 384702 529454
rect 420146 529538 420382 529774
rect 420466 529538 420702 529774
rect 420146 529218 420382 529454
rect 420466 529218 420702 529454
rect 456146 529538 456382 529774
rect 456466 529538 456702 529774
rect 456146 529218 456382 529454
rect 456466 529218 456702 529454
rect 492146 529538 492382 529774
rect 492466 529538 492702 529774
rect 492146 529218 492382 529454
rect 492466 529218 492702 529454
rect 528146 529538 528382 529774
rect 528466 529538 528702 529774
rect 528146 529218 528382 529454
rect 528466 529218 528702 529454
rect 541826 507218 542062 507454
rect 542146 507218 542382 507454
rect 541826 506898 542062 507134
rect 542146 506898 542382 507134
rect 273210 474938 273446 475174
rect 273210 474618 273446 474854
rect 303930 474938 304166 475174
rect 303930 474618 304166 474854
rect 334650 474938 334886 475174
rect 334650 474618 334886 474854
rect 365370 474938 365606 475174
rect 365370 474618 365606 474854
rect 396090 474938 396326 475174
rect 396090 474618 396326 474854
rect 426810 474938 427046 475174
rect 426810 474618 427046 474854
rect 457530 474938 457766 475174
rect 457530 474618 457766 474854
rect 488250 474938 488486 475174
rect 488250 474618 488486 474854
rect 518970 474938 519206 475174
rect 518970 474618 519206 474854
rect 253826 471218 254062 471454
rect 254146 471218 254382 471454
rect 253826 470898 254062 471134
rect 254146 470898 254382 471134
rect 257850 471218 258086 471454
rect 257850 470898 258086 471134
rect 288570 471218 288806 471454
rect 288570 470898 288806 471134
rect 319290 471218 319526 471454
rect 319290 470898 319526 471134
rect 350010 471218 350246 471454
rect 350010 470898 350246 471134
rect 380730 471218 380966 471454
rect 380730 470898 380966 471134
rect 411450 471218 411686 471454
rect 411450 470898 411686 471134
rect 442170 471218 442406 471454
rect 442170 470898 442406 471134
rect 472890 471218 473126 471454
rect 472890 470898 473126 471134
rect 503610 471218 503846 471454
rect 503610 470898 503846 471134
rect 534330 471218 534566 471454
rect 534330 470898 534566 471134
rect 541826 471218 542062 471454
rect 542146 471218 542382 471454
rect 541826 470898 542062 471134
rect 542146 470898 542382 471134
rect 273210 438938 273446 439174
rect 273210 438618 273446 438854
rect 303930 438938 304166 439174
rect 303930 438618 304166 438854
rect 334650 438938 334886 439174
rect 334650 438618 334886 438854
rect 365370 438938 365606 439174
rect 365370 438618 365606 438854
rect 396090 438938 396326 439174
rect 396090 438618 396326 438854
rect 426810 438938 427046 439174
rect 426810 438618 427046 438854
rect 457530 438938 457766 439174
rect 457530 438618 457766 438854
rect 488250 438938 488486 439174
rect 488250 438618 488486 438854
rect 518970 438938 519206 439174
rect 518970 438618 519206 438854
rect 253826 435218 254062 435454
rect 254146 435218 254382 435454
rect 253826 434898 254062 435134
rect 254146 434898 254382 435134
rect 257850 435218 258086 435454
rect 257850 434898 258086 435134
rect 288570 435218 288806 435454
rect 288570 434898 288806 435134
rect 319290 435218 319526 435454
rect 319290 434898 319526 435134
rect 350010 435218 350246 435454
rect 350010 434898 350246 435134
rect 380730 435218 380966 435454
rect 380730 434898 380966 435134
rect 411450 435218 411686 435454
rect 411450 434898 411686 435134
rect 442170 435218 442406 435454
rect 442170 434898 442406 435134
rect 472890 435218 473126 435454
rect 472890 434898 473126 435134
rect 503610 435218 503846 435454
rect 503610 434898 503846 435134
rect 534330 435218 534566 435454
rect 534330 434898 534566 435134
rect 541826 435218 542062 435454
rect 542146 435218 542382 435454
rect 541826 434898 542062 435134
rect 542146 434898 542382 435134
rect 273210 402938 273446 403174
rect 273210 402618 273446 402854
rect 303930 402938 304166 403174
rect 303930 402618 304166 402854
rect 334650 402938 334886 403174
rect 334650 402618 334886 402854
rect 365370 402938 365606 403174
rect 365370 402618 365606 402854
rect 396090 402938 396326 403174
rect 396090 402618 396326 402854
rect 426810 402938 427046 403174
rect 426810 402618 427046 402854
rect 457530 402938 457766 403174
rect 457530 402618 457766 402854
rect 488250 402938 488486 403174
rect 488250 402618 488486 402854
rect 518970 402938 519206 403174
rect 518970 402618 519206 402854
rect 253826 399218 254062 399454
rect 254146 399218 254382 399454
rect 253826 398898 254062 399134
rect 254146 398898 254382 399134
rect 257850 399218 258086 399454
rect 257850 398898 258086 399134
rect 288570 399218 288806 399454
rect 288570 398898 288806 399134
rect 319290 399218 319526 399454
rect 319290 398898 319526 399134
rect 350010 399218 350246 399454
rect 350010 398898 350246 399134
rect 380730 399218 380966 399454
rect 380730 398898 380966 399134
rect 411450 399218 411686 399454
rect 411450 398898 411686 399134
rect 442170 399218 442406 399454
rect 442170 398898 442406 399134
rect 472890 399218 473126 399454
rect 472890 398898 473126 399134
rect 503610 399218 503846 399454
rect 503610 398898 503846 399134
rect 534330 399218 534566 399454
rect 534330 398898 534566 399134
rect 541826 399218 542062 399454
rect 542146 399218 542382 399454
rect 541826 398898 542062 399134
rect 542146 398898 542382 399134
rect 253826 363218 254062 363454
rect 254146 363218 254382 363454
rect 253826 362898 254062 363134
rect 254146 362898 254382 363134
rect 253826 327218 254062 327454
rect 254146 327218 254382 327454
rect 253826 326898 254062 327134
rect 254146 326898 254382 327134
rect 253826 291218 254062 291454
rect 254146 291218 254382 291454
rect 253826 290898 254062 291134
rect 254146 290898 254382 291134
rect 253826 255218 254062 255454
rect 254146 255218 254382 255454
rect 253826 254898 254062 255134
rect 254146 254898 254382 255134
rect 253826 219218 254062 219454
rect 254146 219218 254382 219454
rect 253826 218898 254062 219134
rect 254146 218898 254382 219134
rect 253826 183218 254062 183454
rect 254146 183218 254382 183454
rect 253826 182898 254062 183134
rect 254146 182898 254382 183134
rect 253826 147218 254062 147454
rect 254146 147218 254382 147454
rect 253826 146898 254062 147134
rect 254146 146898 254382 147134
rect 253826 111218 254062 111454
rect 254146 111218 254382 111454
rect 253826 110898 254062 111134
rect 254146 110898 254382 111134
rect 253826 75218 254062 75454
rect 254146 75218 254382 75454
rect 253826 74898 254062 75134
rect 254146 74898 254382 75134
rect 243866 29258 244102 29494
rect 244186 29258 244422 29494
rect 243866 28938 244102 29174
rect 244186 28938 244422 29174
rect 243866 -7302 244102 -7066
rect 244186 -7302 244422 -7066
rect 243866 -7622 244102 -7386
rect 244186 -7622 244422 -7386
rect 253826 39218 254062 39454
rect 254146 39218 254382 39454
rect 253826 38898 254062 39134
rect 254146 38898 254382 39134
rect 253826 3218 254062 3454
rect 254146 3218 254382 3454
rect 253826 2898 254062 3134
rect 254146 2898 254382 3134
rect 253826 -582 254062 -346
rect 254146 -582 254382 -346
rect 253826 -902 254062 -666
rect 254146 -902 254382 -666
rect 257546 366938 257782 367174
rect 257866 366938 258102 367174
rect 257546 366618 257782 366854
rect 257866 366618 258102 366854
rect 257546 330938 257782 331174
rect 257866 330938 258102 331174
rect 257546 330618 257782 330854
rect 257866 330618 258102 330854
rect 261266 370658 261502 370894
rect 261586 370658 261822 370894
rect 261266 370338 261502 370574
rect 261586 370338 261822 370574
rect 261266 334658 261502 334894
rect 261586 334658 261822 334894
rect 261266 334338 261502 334574
rect 261586 334338 261822 334574
rect 264986 374378 265222 374614
rect 265306 374378 265542 374614
rect 264986 374058 265222 374294
rect 265306 374058 265542 374294
rect 264986 338378 265222 338614
rect 265306 338378 265542 338614
rect 264986 338058 265222 338294
rect 265306 338058 265542 338294
rect 268706 378098 268942 378334
rect 269026 378098 269262 378334
rect 268706 377778 268942 378014
rect 269026 377778 269262 378014
rect 268706 342098 268942 342334
rect 269026 342098 269262 342334
rect 268706 341778 268942 342014
rect 269026 341778 269262 342014
rect 289826 363218 290062 363454
rect 290146 363218 290382 363454
rect 289826 362898 290062 363134
rect 290146 362898 290382 363134
rect 289826 327218 290062 327454
rect 290146 327218 290382 327454
rect 289826 326898 290062 327134
rect 290146 326898 290382 327134
rect 293546 366938 293782 367174
rect 293866 366938 294102 367174
rect 293546 366618 293782 366854
rect 293866 366618 294102 366854
rect 293546 330938 293782 331174
rect 293866 330938 294102 331174
rect 293546 330618 293782 330854
rect 293866 330618 294102 330854
rect 297266 370658 297502 370894
rect 297586 370658 297822 370894
rect 297266 370338 297502 370574
rect 297586 370338 297822 370574
rect 297266 334658 297502 334894
rect 297586 334658 297822 334894
rect 297266 334338 297502 334574
rect 297586 334338 297822 334574
rect 300986 374378 301222 374614
rect 301306 374378 301542 374614
rect 300986 374058 301222 374294
rect 301306 374058 301542 374294
rect 300986 338378 301222 338614
rect 301306 338378 301542 338614
rect 300986 338058 301222 338294
rect 301306 338058 301542 338294
rect 304706 378098 304942 378334
rect 305026 378098 305262 378334
rect 304706 377778 304942 378014
rect 305026 377778 305262 378014
rect 304706 342098 304942 342334
rect 305026 342098 305262 342334
rect 304706 341778 304942 342014
rect 305026 341778 305262 342014
rect 325826 363218 326062 363454
rect 326146 363218 326382 363454
rect 325826 362898 326062 363134
rect 326146 362898 326382 363134
rect 325826 327218 326062 327454
rect 326146 327218 326382 327454
rect 325826 326898 326062 327134
rect 326146 326898 326382 327134
rect 329546 366938 329782 367174
rect 329866 366938 330102 367174
rect 329546 366618 329782 366854
rect 329866 366618 330102 366854
rect 329546 330938 329782 331174
rect 329866 330938 330102 331174
rect 329546 330618 329782 330854
rect 329866 330618 330102 330854
rect 333266 370658 333502 370894
rect 333586 370658 333822 370894
rect 333266 370338 333502 370574
rect 333586 370338 333822 370574
rect 333266 334658 333502 334894
rect 333586 334658 333822 334894
rect 333266 334338 333502 334574
rect 333586 334338 333822 334574
rect 336986 374378 337222 374614
rect 337306 374378 337542 374614
rect 336986 374058 337222 374294
rect 337306 374058 337542 374294
rect 336986 338378 337222 338614
rect 337306 338378 337542 338614
rect 336986 338058 337222 338294
rect 337306 338058 337542 338294
rect 340706 378098 340942 378334
rect 341026 378098 341262 378334
rect 340706 377778 340942 378014
rect 341026 377778 341262 378014
rect 340706 342098 340942 342334
rect 341026 342098 341262 342334
rect 340706 341778 340942 342014
rect 341026 341778 341262 342014
rect 361826 363218 362062 363454
rect 362146 363218 362382 363454
rect 361826 362898 362062 363134
rect 362146 362898 362382 363134
rect 361826 327218 362062 327454
rect 362146 327218 362382 327454
rect 361826 326898 362062 327134
rect 362146 326898 362382 327134
rect 365546 366938 365782 367174
rect 365866 366938 366102 367174
rect 365546 366618 365782 366854
rect 365866 366618 366102 366854
rect 365546 330938 365782 331174
rect 365866 330938 366102 331174
rect 365546 330618 365782 330854
rect 365866 330618 366102 330854
rect 369266 370658 369502 370894
rect 369586 370658 369822 370894
rect 369266 370338 369502 370574
rect 369586 370338 369822 370574
rect 369266 334658 369502 334894
rect 369586 334658 369822 334894
rect 369266 334338 369502 334574
rect 369586 334338 369822 334574
rect 372986 374378 373222 374614
rect 373306 374378 373542 374614
rect 372986 374058 373222 374294
rect 373306 374058 373542 374294
rect 372986 338378 373222 338614
rect 373306 338378 373542 338614
rect 372986 338058 373222 338294
rect 373306 338058 373542 338294
rect 376706 378098 376942 378334
rect 377026 378098 377262 378334
rect 376706 377778 376942 378014
rect 377026 377778 377262 378014
rect 376706 342098 376942 342334
rect 377026 342098 377262 342334
rect 376706 341778 376942 342014
rect 377026 341778 377262 342014
rect 397826 363218 398062 363454
rect 398146 363218 398382 363454
rect 397826 362898 398062 363134
rect 398146 362898 398382 363134
rect 397826 327218 398062 327454
rect 398146 327218 398382 327454
rect 397826 326898 398062 327134
rect 398146 326898 398382 327134
rect 401546 366938 401782 367174
rect 401866 366938 402102 367174
rect 401546 366618 401782 366854
rect 401866 366618 402102 366854
rect 401546 330938 401782 331174
rect 401866 330938 402102 331174
rect 401546 330618 401782 330854
rect 401866 330618 402102 330854
rect 405266 370658 405502 370894
rect 405586 370658 405822 370894
rect 405266 370338 405502 370574
rect 405586 370338 405822 370574
rect 405266 334658 405502 334894
rect 405586 334658 405822 334894
rect 405266 334338 405502 334574
rect 405586 334338 405822 334574
rect 408986 374378 409222 374614
rect 409306 374378 409542 374614
rect 408986 374058 409222 374294
rect 409306 374058 409542 374294
rect 408986 338378 409222 338614
rect 409306 338378 409542 338614
rect 408986 338058 409222 338294
rect 409306 338058 409542 338294
rect 412706 378098 412942 378334
rect 413026 378098 413262 378334
rect 412706 377778 412942 378014
rect 413026 377778 413262 378014
rect 412706 342098 412942 342334
rect 413026 342098 413262 342334
rect 412706 341778 412942 342014
rect 413026 341778 413262 342014
rect 433826 363218 434062 363454
rect 434146 363218 434382 363454
rect 433826 362898 434062 363134
rect 434146 362898 434382 363134
rect 433826 327218 434062 327454
rect 434146 327218 434382 327454
rect 433826 326898 434062 327134
rect 434146 326898 434382 327134
rect 437546 366938 437782 367174
rect 437866 366938 438102 367174
rect 437546 366618 437782 366854
rect 437866 366618 438102 366854
rect 437546 330938 437782 331174
rect 437866 330938 438102 331174
rect 437546 330618 437782 330854
rect 437866 330618 438102 330854
rect 441266 370658 441502 370894
rect 441586 370658 441822 370894
rect 441266 370338 441502 370574
rect 441586 370338 441822 370574
rect 441266 334658 441502 334894
rect 441586 334658 441822 334894
rect 441266 334338 441502 334574
rect 441586 334338 441822 334574
rect 444986 374378 445222 374614
rect 445306 374378 445542 374614
rect 444986 374058 445222 374294
rect 445306 374058 445542 374294
rect 444986 338378 445222 338614
rect 445306 338378 445542 338614
rect 444986 338058 445222 338294
rect 445306 338058 445542 338294
rect 448706 378098 448942 378334
rect 449026 378098 449262 378334
rect 448706 377778 448942 378014
rect 449026 377778 449262 378014
rect 448706 342098 448942 342334
rect 449026 342098 449262 342334
rect 448706 341778 448942 342014
rect 449026 341778 449262 342014
rect 469826 363218 470062 363454
rect 470146 363218 470382 363454
rect 469826 362898 470062 363134
rect 470146 362898 470382 363134
rect 469826 327218 470062 327454
rect 470146 327218 470382 327454
rect 469826 326898 470062 327134
rect 470146 326898 470382 327134
rect 473546 366938 473782 367174
rect 473866 366938 474102 367174
rect 473546 366618 473782 366854
rect 473866 366618 474102 366854
rect 473546 330938 473782 331174
rect 473866 330938 474102 331174
rect 473546 330618 473782 330854
rect 473866 330618 474102 330854
rect 477266 370658 477502 370894
rect 477586 370658 477822 370894
rect 477266 370338 477502 370574
rect 477586 370338 477822 370574
rect 477266 334658 477502 334894
rect 477586 334658 477822 334894
rect 477266 334338 477502 334574
rect 477586 334338 477822 334574
rect 480986 374378 481222 374614
rect 481306 374378 481542 374614
rect 480986 374058 481222 374294
rect 481306 374058 481542 374294
rect 480986 338378 481222 338614
rect 481306 338378 481542 338614
rect 480986 338058 481222 338294
rect 481306 338058 481542 338294
rect 484706 378098 484942 378334
rect 485026 378098 485262 378334
rect 484706 377778 484942 378014
rect 485026 377778 485262 378014
rect 484706 342098 484942 342334
rect 485026 342098 485262 342334
rect 484706 341778 484942 342014
rect 485026 341778 485262 342014
rect 505826 363218 506062 363454
rect 506146 363218 506382 363454
rect 505826 362898 506062 363134
rect 506146 362898 506382 363134
rect 505826 327218 506062 327454
rect 506146 327218 506382 327454
rect 505826 326898 506062 327134
rect 506146 326898 506382 327134
rect 509546 366938 509782 367174
rect 509866 366938 510102 367174
rect 509546 366618 509782 366854
rect 509866 366618 510102 366854
rect 509546 330938 509782 331174
rect 509866 330938 510102 331174
rect 509546 330618 509782 330854
rect 509866 330618 510102 330854
rect 513266 370658 513502 370894
rect 513586 370658 513822 370894
rect 513266 370338 513502 370574
rect 513586 370338 513822 370574
rect 513266 334658 513502 334894
rect 513586 334658 513822 334894
rect 513266 334338 513502 334574
rect 513586 334338 513822 334574
rect 516986 374378 517222 374614
rect 517306 374378 517542 374614
rect 516986 374058 517222 374294
rect 517306 374058 517542 374294
rect 516986 338378 517222 338614
rect 517306 338378 517542 338614
rect 516986 338058 517222 338294
rect 517306 338058 517542 338294
rect 520706 378098 520942 378334
rect 521026 378098 521262 378334
rect 520706 377778 520942 378014
rect 521026 377778 521262 378014
rect 520706 342098 520942 342334
rect 521026 342098 521262 342334
rect 520706 341778 520942 342014
rect 521026 341778 521262 342014
rect 541826 363218 542062 363454
rect 542146 363218 542382 363454
rect 541826 362898 542062 363134
rect 542146 362898 542382 363134
rect 541826 327218 542062 327454
rect 542146 327218 542382 327454
rect 541826 326898 542062 327134
rect 542146 326898 542382 327134
rect 545546 705562 545782 705798
rect 545866 705562 546102 705798
rect 545546 705242 545782 705478
rect 545866 705242 546102 705478
rect 545546 690938 545782 691174
rect 545866 690938 546102 691174
rect 545546 690618 545782 690854
rect 545866 690618 546102 690854
rect 545546 654938 545782 655174
rect 545866 654938 546102 655174
rect 545546 654618 545782 654854
rect 545866 654618 546102 654854
rect 549266 706522 549502 706758
rect 549586 706522 549822 706758
rect 549266 706202 549502 706438
rect 549586 706202 549822 706438
rect 549266 694658 549502 694894
rect 549586 694658 549822 694894
rect 549266 694338 549502 694574
rect 549586 694338 549822 694574
rect 549266 658658 549502 658894
rect 549586 658658 549822 658894
rect 549266 658338 549502 658574
rect 549586 658338 549822 658574
rect 552986 707482 553222 707718
rect 553306 707482 553542 707718
rect 552986 707162 553222 707398
rect 553306 707162 553542 707398
rect 552986 698378 553222 698614
rect 553306 698378 553542 698614
rect 552986 698058 553222 698294
rect 553306 698058 553542 698294
rect 552986 662378 553222 662614
rect 553306 662378 553542 662614
rect 552986 662058 553222 662294
rect 553306 662058 553542 662294
rect 552986 626378 553222 626614
rect 553306 626378 553542 626614
rect 552986 626058 553222 626294
rect 553306 626058 553542 626294
rect 545546 618938 545782 619174
rect 545866 618938 546102 619174
rect 545546 618618 545782 618854
rect 545866 618618 546102 618854
rect 549690 618938 549926 619174
rect 549690 618618 549926 618854
rect 552986 590378 553222 590614
rect 553306 590378 553542 590614
rect 552986 590058 553222 590294
rect 553306 590058 553542 590294
rect 545546 582938 545782 583174
rect 545866 582938 546102 583174
rect 545546 582618 545782 582854
rect 545866 582618 546102 582854
rect 549690 582938 549926 583174
rect 549690 582618 549926 582854
rect 552986 554378 553222 554614
rect 553306 554378 553542 554614
rect 552986 554058 553222 554294
rect 553306 554058 553542 554294
rect 545546 546938 545782 547174
rect 545866 546938 546102 547174
rect 545546 546618 545782 546854
rect 545866 546618 546102 546854
rect 549690 546938 549926 547174
rect 549690 546618 549926 546854
rect 545546 510938 545782 511174
rect 545866 510938 546102 511174
rect 545546 510618 545782 510854
rect 545866 510618 546102 510854
rect 552986 518378 553222 518614
rect 553306 518378 553542 518614
rect 552986 518058 553222 518294
rect 553306 518058 553542 518294
rect 552986 482378 553222 482614
rect 553306 482378 553542 482614
rect 552986 482058 553222 482294
rect 553306 482058 553542 482294
rect 545546 474938 545782 475174
rect 545866 474938 546102 475174
rect 545546 474618 545782 474854
rect 545866 474618 546102 474854
rect 549690 474938 549926 475174
rect 549690 474618 549926 474854
rect 552986 446378 553222 446614
rect 553306 446378 553542 446614
rect 552986 446058 553222 446294
rect 553306 446058 553542 446294
rect 545546 438938 545782 439174
rect 545866 438938 546102 439174
rect 545546 438618 545782 438854
rect 545866 438618 546102 438854
rect 549690 438938 549926 439174
rect 549690 438618 549926 438854
rect 552986 410378 553222 410614
rect 553306 410378 553542 410614
rect 552986 410058 553222 410294
rect 553306 410058 553542 410294
rect 545546 402938 545782 403174
rect 545866 402938 546102 403174
rect 545546 402618 545782 402854
rect 545866 402618 546102 402854
rect 549690 402938 549926 403174
rect 549690 402618 549926 402854
rect 545546 366938 545782 367174
rect 545866 366938 546102 367174
rect 545546 366618 545782 366854
rect 545866 366618 546102 366854
rect 545546 330938 545782 331174
rect 545866 330938 546102 331174
rect 545546 330618 545782 330854
rect 545866 330618 546102 330854
rect 549266 370658 549502 370894
rect 549586 370658 549822 370894
rect 549266 370338 549502 370574
rect 549586 370338 549822 370574
rect 549266 334658 549502 334894
rect 549586 334658 549822 334894
rect 549266 334338 549502 334574
rect 549586 334338 549822 334574
rect 552986 374378 553222 374614
rect 553306 374378 553542 374614
rect 552986 374058 553222 374294
rect 553306 374058 553542 374294
rect 552986 338378 553222 338614
rect 553306 338378 553542 338614
rect 552986 338058 553222 338294
rect 553306 338058 553542 338294
rect 552986 302378 553222 302614
rect 553306 302378 553542 302614
rect 552986 302058 553222 302294
rect 553306 302058 553542 302294
rect 257546 294938 257782 295174
rect 257866 294938 258102 295174
rect 257546 294618 257782 294854
rect 257866 294618 258102 294854
rect 279610 294938 279846 295174
rect 279610 294618 279846 294854
rect 310330 294938 310566 295174
rect 310330 294618 310566 294854
rect 341050 294938 341286 295174
rect 341050 294618 341286 294854
rect 371770 294938 372006 295174
rect 371770 294618 372006 294854
rect 402490 294938 402726 295174
rect 402490 294618 402726 294854
rect 433210 294938 433446 295174
rect 433210 294618 433446 294854
rect 463930 294938 464166 295174
rect 463930 294618 464166 294854
rect 494650 294938 494886 295174
rect 494650 294618 494886 294854
rect 525370 294938 525606 295174
rect 525370 294618 525606 294854
rect 264250 291218 264486 291454
rect 264250 290898 264486 291134
rect 294970 291218 295206 291454
rect 294970 290898 295206 291134
rect 325690 291218 325926 291454
rect 325690 290898 325926 291134
rect 356410 291218 356646 291454
rect 356410 290898 356646 291134
rect 387130 291218 387366 291454
rect 387130 290898 387366 291134
rect 417850 291218 418086 291454
rect 417850 290898 418086 291134
rect 448570 291218 448806 291454
rect 448570 290898 448806 291134
rect 479290 291218 479526 291454
rect 479290 290898 479526 291134
rect 510010 291218 510246 291454
rect 510010 290898 510246 291134
rect 540730 291218 540966 291454
rect 540730 290898 540966 291134
rect 552986 266378 553222 266614
rect 553306 266378 553542 266614
rect 552986 266058 553222 266294
rect 553306 266058 553542 266294
rect 257546 258938 257782 259174
rect 257866 258938 258102 259174
rect 257546 258618 257782 258854
rect 257866 258618 258102 258854
rect 279610 258938 279846 259174
rect 279610 258618 279846 258854
rect 310330 258938 310566 259174
rect 310330 258618 310566 258854
rect 341050 258938 341286 259174
rect 341050 258618 341286 258854
rect 371770 258938 372006 259174
rect 371770 258618 372006 258854
rect 402490 258938 402726 259174
rect 402490 258618 402726 258854
rect 433210 258938 433446 259174
rect 433210 258618 433446 258854
rect 463930 258938 464166 259174
rect 463930 258618 464166 258854
rect 494650 258938 494886 259174
rect 494650 258618 494886 258854
rect 525370 258938 525606 259174
rect 525370 258618 525606 258854
rect 264250 255218 264486 255454
rect 264250 254898 264486 255134
rect 294970 255218 295206 255454
rect 294970 254898 295206 255134
rect 325690 255218 325926 255454
rect 325690 254898 325926 255134
rect 356410 255218 356646 255454
rect 356410 254898 356646 255134
rect 387130 255218 387366 255454
rect 387130 254898 387366 255134
rect 417850 255218 418086 255454
rect 417850 254898 418086 255134
rect 448570 255218 448806 255454
rect 448570 254898 448806 255134
rect 479290 255218 479526 255454
rect 479290 254898 479526 255134
rect 510010 255218 510246 255454
rect 510010 254898 510246 255134
rect 540730 255218 540966 255454
rect 540730 254898 540966 255134
rect 552986 230378 553222 230614
rect 553306 230378 553542 230614
rect 552986 230058 553222 230294
rect 553306 230058 553542 230294
rect 257546 222938 257782 223174
rect 257866 222938 258102 223174
rect 257546 222618 257782 222854
rect 257866 222618 258102 222854
rect 279610 222938 279846 223174
rect 279610 222618 279846 222854
rect 310330 222938 310566 223174
rect 310330 222618 310566 222854
rect 341050 222938 341286 223174
rect 341050 222618 341286 222854
rect 371770 222938 372006 223174
rect 371770 222618 372006 222854
rect 402490 222938 402726 223174
rect 402490 222618 402726 222854
rect 433210 222938 433446 223174
rect 433210 222618 433446 222854
rect 463930 222938 464166 223174
rect 463930 222618 464166 222854
rect 494650 222938 494886 223174
rect 494650 222618 494886 222854
rect 525370 222938 525606 223174
rect 525370 222618 525606 222854
rect 264250 219218 264486 219454
rect 264250 218898 264486 219134
rect 294970 219218 295206 219454
rect 294970 218898 295206 219134
rect 325690 219218 325926 219454
rect 325690 218898 325926 219134
rect 356410 219218 356646 219454
rect 356410 218898 356646 219134
rect 387130 219218 387366 219454
rect 387130 218898 387366 219134
rect 417850 219218 418086 219454
rect 417850 218898 418086 219134
rect 448570 219218 448806 219454
rect 448570 218898 448806 219134
rect 479290 219218 479526 219454
rect 479290 218898 479526 219134
rect 510010 219218 510246 219454
rect 510010 218898 510246 219134
rect 540730 219218 540966 219454
rect 540730 218898 540966 219134
rect 552986 194378 553222 194614
rect 553306 194378 553542 194614
rect 552986 194058 553222 194294
rect 553306 194058 553542 194294
rect 257546 186938 257782 187174
rect 257866 186938 258102 187174
rect 257546 186618 257782 186854
rect 257866 186618 258102 186854
rect 279610 186938 279846 187174
rect 279610 186618 279846 186854
rect 310330 186938 310566 187174
rect 310330 186618 310566 186854
rect 341050 186938 341286 187174
rect 341050 186618 341286 186854
rect 371770 186938 372006 187174
rect 371770 186618 372006 186854
rect 402490 186938 402726 187174
rect 402490 186618 402726 186854
rect 433210 186938 433446 187174
rect 433210 186618 433446 186854
rect 463930 186938 464166 187174
rect 463930 186618 464166 186854
rect 494650 186938 494886 187174
rect 494650 186618 494886 186854
rect 525370 186938 525606 187174
rect 525370 186618 525606 186854
rect 264250 183218 264486 183454
rect 264250 182898 264486 183134
rect 294970 183218 295206 183454
rect 294970 182898 295206 183134
rect 325690 183218 325926 183454
rect 325690 182898 325926 183134
rect 356410 183218 356646 183454
rect 356410 182898 356646 183134
rect 387130 183218 387366 183454
rect 387130 182898 387366 183134
rect 417850 183218 418086 183454
rect 417850 182898 418086 183134
rect 448570 183218 448806 183454
rect 448570 182898 448806 183134
rect 479290 183218 479526 183454
rect 479290 182898 479526 183134
rect 510010 183218 510246 183454
rect 510010 182898 510246 183134
rect 540730 183218 540966 183454
rect 540730 182898 540966 183134
rect 552986 158378 553222 158614
rect 553306 158378 553542 158614
rect 552986 158058 553222 158294
rect 553306 158058 553542 158294
rect 257546 150938 257782 151174
rect 257866 150938 258102 151174
rect 257546 150618 257782 150854
rect 257866 150618 258102 150854
rect 279610 150938 279846 151174
rect 279610 150618 279846 150854
rect 310330 150938 310566 151174
rect 310330 150618 310566 150854
rect 341050 150938 341286 151174
rect 341050 150618 341286 150854
rect 371770 150938 372006 151174
rect 371770 150618 372006 150854
rect 402490 150938 402726 151174
rect 402490 150618 402726 150854
rect 433210 150938 433446 151174
rect 433210 150618 433446 150854
rect 463930 150938 464166 151174
rect 463930 150618 464166 150854
rect 494650 150938 494886 151174
rect 494650 150618 494886 150854
rect 525370 150938 525606 151174
rect 525370 150618 525606 150854
rect 264250 147218 264486 147454
rect 264250 146898 264486 147134
rect 294970 147218 295206 147454
rect 294970 146898 295206 147134
rect 325690 147218 325926 147454
rect 325690 146898 325926 147134
rect 356410 147218 356646 147454
rect 356410 146898 356646 147134
rect 387130 147218 387366 147454
rect 387130 146898 387366 147134
rect 417850 147218 418086 147454
rect 417850 146898 418086 147134
rect 448570 147218 448806 147454
rect 448570 146898 448806 147134
rect 479290 147218 479526 147454
rect 479290 146898 479526 147134
rect 510010 147218 510246 147454
rect 510010 146898 510246 147134
rect 540730 147218 540966 147454
rect 540730 146898 540966 147134
rect 552986 122378 553222 122614
rect 553306 122378 553542 122614
rect 552986 122058 553222 122294
rect 553306 122058 553542 122294
rect 257546 114938 257782 115174
rect 257866 114938 258102 115174
rect 257546 114618 257782 114854
rect 257866 114618 258102 114854
rect 279610 114938 279846 115174
rect 279610 114618 279846 114854
rect 310330 114938 310566 115174
rect 310330 114618 310566 114854
rect 341050 114938 341286 115174
rect 341050 114618 341286 114854
rect 371770 114938 372006 115174
rect 371770 114618 372006 114854
rect 402490 114938 402726 115174
rect 402490 114618 402726 114854
rect 433210 114938 433446 115174
rect 433210 114618 433446 114854
rect 463930 114938 464166 115174
rect 463930 114618 464166 114854
rect 494650 114938 494886 115174
rect 494650 114618 494886 114854
rect 525370 114938 525606 115174
rect 525370 114618 525606 114854
rect 264250 111218 264486 111454
rect 264250 110898 264486 111134
rect 294970 111218 295206 111454
rect 294970 110898 295206 111134
rect 325690 111218 325926 111454
rect 325690 110898 325926 111134
rect 356410 111218 356646 111454
rect 356410 110898 356646 111134
rect 387130 111218 387366 111454
rect 387130 110898 387366 111134
rect 417850 111218 418086 111454
rect 417850 110898 418086 111134
rect 448570 111218 448806 111454
rect 448570 110898 448806 111134
rect 479290 111218 479526 111454
rect 479290 110898 479526 111134
rect 510010 111218 510246 111454
rect 510010 110898 510246 111134
rect 540730 111218 540966 111454
rect 540730 110898 540966 111134
rect 552986 86378 553222 86614
rect 553306 86378 553542 86614
rect 552986 86058 553222 86294
rect 553306 86058 553542 86294
rect 257546 78938 257782 79174
rect 257866 78938 258102 79174
rect 257546 78618 257782 78854
rect 257866 78618 258102 78854
rect 279610 78938 279846 79174
rect 279610 78618 279846 78854
rect 310330 78938 310566 79174
rect 310330 78618 310566 78854
rect 341050 78938 341286 79174
rect 341050 78618 341286 78854
rect 371770 78938 372006 79174
rect 371770 78618 372006 78854
rect 402490 78938 402726 79174
rect 402490 78618 402726 78854
rect 433210 78938 433446 79174
rect 433210 78618 433446 78854
rect 463930 78938 464166 79174
rect 463930 78618 464166 78854
rect 494650 78938 494886 79174
rect 494650 78618 494886 78854
rect 525370 78938 525606 79174
rect 525370 78618 525606 78854
rect 264250 75218 264486 75454
rect 264250 74898 264486 75134
rect 294970 75218 295206 75454
rect 294970 74898 295206 75134
rect 325690 75218 325926 75454
rect 325690 74898 325926 75134
rect 356410 75218 356646 75454
rect 356410 74898 356646 75134
rect 387130 75218 387366 75454
rect 387130 74898 387366 75134
rect 417850 75218 418086 75454
rect 417850 74898 418086 75134
rect 448570 75218 448806 75454
rect 448570 74898 448806 75134
rect 479290 75218 479526 75454
rect 479290 74898 479526 75134
rect 510010 75218 510246 75454
rect 510010 74898 510246 75134
rect 540730 75218 540966 75454
rect 540730 74898 540966 75134
rect 552986 50378 553222 50614
rect 553306 50378 553542 50614
rect 257546 42938 257782 43174
rect 257866 42938 258102 43174
rect 257546 42618 257782 42854
rect 257866 42618 258102 42854
rect 257546 6938 257782 7174
rect 257866 6938 258102 7174
rect 257546 6618 257782 6854
rect 257866 6618 258102 6854
rect 552986 50058 553222 50294
rect 553306 50058 553542 50294
rect 261266 10658 261502 10894
rect 261586 10658 261822 10894
rect 261266 10338 261502 10574
rect 261586 10338 261822 10574
rect 257546 -1542 257782 -1306
rect 257866 -1542 258102 -1306
rect 257546 -1862 257782 -1626
rect 257866 -1862 258102 -1626
rect 261266 -2502 261502 -2266
rect 261586 -2502 261822 -2266
rect 261266 -2822 261502 -2586
rect 261586 -2822 261822 -2586
rect 264986 14378 265222 14614
rect 265306 14378 265542 14614
rect 264986 14058 265222 14294
rect 265306 14058 265542 14294
rect 264986 -3462 265222 -3226
rect 265306 -3462 265542 -3226
rect 264986 -3782 265222 -3546
rect 265306 -3782 265542 -3546
rect 268706 18098 268942 18334
rect 269026 18098 269262 18334
rect 268706 17778 268942 18014
rect 269026 17778 269262 18014
rect 268706 -4422 268942 -4186
rect 269026 -4422 269262 -4186
rect 268706 -4742 268942 -4506
rect 269026 -4742 269262 -4506
rect 272426 21818 272662 22054
rect 272746 21818 272982 22054
rect 272426 21498 272662 21734
rect 272746 21498 272982 21734
rect 272426 -5382 272662 -5146
rect 272746 -5382 272982 -5146
rect 272426 -5702 272662 -5466
rect 272746 -5702 272982 -5466
rect 279610 42938 279846 43174
rect 279610 42618 279846 42854
rect 276146 25538 276382 25774
rect 276466 25538 276702 25774
rect 276146 25218 276382 25454
rect 276466 25218 276702 25454
rect 276146 -6342 276382 -6106
rect 276466 -6342 276702 -6106
rect 276146 -6662 276382 -6426
rect 276466 -6662 276702 -6426
rect 279866 29258 280102 29494
rect 280186 29258 280422 29494
rect 279866 28938 280102 29174
rect 280186 28938 280422 29174
rect 279866 -7302 280102 -7066
rect 280186 -7302 280422 -7066
rect 279866 -7622 280102 -7386
rect 280186 -7622 280422 -7386
rect 289826 39218 290062 39454
rect 290146 39218 290382 39454
rect 289826 38898 290062 39134
rect 290146 38898 290382 39134
rect 289826 3218 290062 3454
rect 290146 3218 290382 3454
rect 289826 2898 290062 3134
rect 290146 2898 290382 3134
rect 289826 -582 290062 -346
rect 290146 -582 290382 -346
rect 289826 -902 290062 -666
rect 290146 -902 290382 -666
rect 293546 6938 293782 7174
rect 293866 6938 294102 7174
rect 293546 6618 293782 6854
rect 293866 6618 294102 6854
rect 293546 -1542 293782 -1306
rect 293866 -1542 294102 -1306
rect 293546 -1862 293782 -1626
rect 293866 -1862 294102 -1626
rect 297266 10658 297502 10894
rect 297586 10658 297822 10894
rect 297266 10338 297502 10574
rect 297586 10338 297822 10574
rect 297266 -2502 297502 -2266
rect 297586 -2502 297822 -2266
rect 297266 -2822 297502 -2586
rect 297586 -2822 297822 -2586
rect 300986 14378 301222 14614
rect 301306 14378 301542 14614
rect 300986 14058 301222 14294
rect 301306 14058 301542 14294
rect 300986 -3462 301222 -3226
rect 301306 -3462 301542 -3226
rect 300986 -3782 301222 -3546
rect 301306 -3782 301542 -3546
rect 304706 18098 304942 18334
rect 305026 18098 305262 18334
rect 304706 17778 304942 18014
rect 305026 17778 305262 18014
rect 304706 -4422 304942 -4186
rect 305026 -4422 305262 -4186
rect 304706 -4742 304942 -4506
rect 305026 -4742 305262 -4506
rect 310330 42938 310566 43174
rect 310330 42618 310566 42854
rect 308426 21818 308662 22054
rect 308746 21818 308982 22054
rect 308426 21498 308662 21734
rect 308746 21498 308982 21734
rect 308426 -5382 308662 -5146
rect 308746 -5382 308982 -5146
rect 308426 -5702 308662 -5466
rect 308746 -5702 308982 -5466
rect 312146 25538 312382 25774
rect 312466 25538 312702 25774
rect 312146 25218 312382 25454
rect 312466 25218 312702 25454
rect 312146 -6342 312382 -6106
rect 312466 -6342 312702 -6106
rect 312146 -6662 312382 -6426
rect 312466 -6662 312702 -6426
rect 315866 29258 316102 29494
rect 316186 29258 316422 29494
rect 315866 28938 316102 29174
rect 316186 28938 316422 29174
rect 315866 -7302 316102 -7066
rect 316186 -7302 316422 -7066
rect 315866 -7622 316102 -7386
rect 316186 -7622 316422 -7386
rect 325826 39218 326062 39454
rect 326146 39218 326382 39454
rect 325826 38898 326062 39134
rect 326146 38898 326382 39134
rect 325826 3218 326062 3454
rect 326146 3218 326382 3454
rect 325826 2898 326062 3134
rect 326146 2898 326382 3134
rect 325826 -582 326062 -346
rect 326146 -582 326382 -346
rect 325826 -902 326062 -666
rect 326146 -902 326382 -666
rect 329546 6938 329782 7174
rect 329866 6938 330102 7174
rect 329546 6618 329782 6854
rect 329866 6618 330102 6854
rect 329546 -1542 329782 -1306
rect 329866 -1542 330102 -1306
rect 329546 -1862 329782 -1626
rect 329866 -1862 330102 -1626
rect 333266 10658 333502 10894
rect 333586 10658 333822 10894
rect 333266 10338 333502 10574
rect 333586 10338 333822 10574
rect 333266 -2502 333502 -2266
rect 333586 -2502 333822 -2266
rect 333266 -2822 333502 -2586
rect 333586 -2822 333822 -2586
rect 341050 42938 341286 43174
rect 341050 42618 341286 42854
rect 336986 14378 337222 14614
rect 337306 14378 337542 14614
rect 336986 14058 337222 14294
rect 337306 14058 337542 14294
rect 336986 -3462 337222 -3226
rect 337306 -3462 337542 -3226
rect 336986 -3782 337222 -3546
rect 337306 -3782 337542 -3546
rect 340706 18098 340942 18334
rect 341026 18098 341262 18334
rect 340706 17778 340942 18014
rect 341026 17778 341262 18014
rect 340706 -4422 340942 -4186
rect 341026 -4422 341262 -4186
rect 340706 -4742 340942 -4506
rect 341026 -4742 341262 -4506
rect 344426 21818 344662 22054
rect 344746 21818 344982 22054
rect 344426 21498 344662 21734
rect 344746 21498 344982 21734
rect 344426 -5382 344662 -5146
rect 344746 -5382 344982 -5146
rect 344426 -5702 344662 -5466
rect 344746 -5702 344982 -5466
rect 348146 25538 348382 25774
rect 348466 25538 348702 25774
rect 348146 25218 348382 25454
rect 348466 25218 348702 25454
rect 348146 -6342 348382 -6106
rect 348466 -6342 348702 -6106
rect 348146 -6662 348382 -6426
rect 348466 -6662 348702 -6426
rect 351866 29258 352102 29494
rect 352186 29258 352422 29494
rect 351866 28938 352102 29174
rect 352186 28938 352422 29174
rect 351866 -7302 352102 -7066
rect 352186 -7302 352422 -7066
rect 351866 -7622 352102 -7386
rect 352186 -7622 352422 -7386
rect 361826 39218 362062 39454
rect 362146 39218 362382 39454
rect 361826 38898 362062 39134
rect 362146 38898 362382 39134
rect 361826 3218 362062 3454
rect 362146 3218 362382 3454
rect 361826 2898 362062 3134
rect 362146 2898 362382 3134
rect 361826 -582 362062 -346
rect 362146 -582 362382 -346
rect 361826 -902 362062 -666
rect 362146 -902 362382 -666
rect 365546 6938 365782 7174
rect 365866 6938 366102 7174
rect 365546 6618 365782 6854
rect 365866 6618 366102 6854
rect 365546 -1542 365782 -1306
rect 365866 -1542 366102 -1306
rect 365546 -1862 365782 -1626
rect 365866 -1862 366102 -1626
rect 371770 42938 372006 43174
rect 371770 42618 372006 42854
rect 369266 10658 369502 10894
rect 369586 10658 369822 10894
rect 369266 10338 369502 10574
rect 369586 10338 369822 10574
rect 369266 -2502 369502 -2266
rect 369586 -2502 369822 -2266
rect 369266 -2822 369502 -2586
rect 369586 -2822 369822 -2586
rect 372986 14378 373222 14614
rect 373306 14378 373542 14614
rect 372986 14058 373222 14294
rect 373306 14058 373542 14294
rect 372986 -3462 373222 -3226
rect 373306 -3462 373542 -3226
rect 372986 -3782 373222 -3546
rect 373306 -3782 373542 -3546
rect 376706 18098 376942 18334
rect 377026 18098 377262 18334
rect 376706 17778 376942 18014
rect 377026 17778 377262 18014
rect 376706 -4422 376942 -4186
rect 377026 -4422 377262 -4186
rect 376706 -4742 376942 -4506
rect 377026 -4742 377262 -4506
rect 380426 21818 380662 22054
rect 380746 21818 380982 22054
rect 380426 21498 380662 21734
rect 380746 21498 380982 21734
rect 380426 -5382 380662 -5146
rect 380746 -5382 380982 -5146
rect 380426 -5702 380662 -5466
rect 380746 -5702 380982 -5466
rect 384146 25538 384382 25774
rect 384466 25538 384702 25774
rect 384146 25218 384382 25454
rect 384466 25218 384702 25454
rect 384146 -6342 384382 -6106
rect 384466 -6342 384702 -6106
rect 384146 -6662 384382 -6426
rect 384466 -6662 384702 -6426
rect 387866 29258 388102 29494
rect 388186 29258 388422 29494
rect 387866 28938 388102 29174
rect 388186 28938 388422 29174
rect 387866 -7302 388102 -7066
rect 388186 -7302 388422 -7066
rect 387866 -7622 388102 -7386
rect 388186 -7622 388422 -7386
rect 397826 39218 398062 39454
rect 398146 39218 398382 39454
rect 397826 38898 398062 39134
rect 398146 38898 398382 39134
rect 397826 3218 398062 3454
rect 398146 3218 398382 3454
rect 397826 2898 398062 3134
rect 398146 2898 398382 3134
rect 397826 -582 398062 -346
rect 398146 -582 398382 -346
rect 397826 -902 398062 -666
rect 398146 -902 398382 -666
rect 402490 42938 402726 43174
rect 402490 42618 402726 42854
rect 401546 6938 401782 7174
rect 401866 6938 402102 7174
rect 401546 6618 401782 6854
rect 401866 6618 402102 6854
rect 401546 -1542 401782 -1306
rect 401866 -1542 402102 -1306
rect 401546 -1862 401782 -1626
rect 401866 -1862 402102 -1626
rect 405266 10658 405502 10894
rect 405586 10658 405822 10894
rect 405266 10338 405502 10574
rect 405586 10338 405822 10574
rect 405266 -2502 405502 -2266
rect 405586 -2502 405822 -2266
rect 405266 -2822 405502 -2586
rect 405586 -2822 405822 -2586
rect 408986 14378 409222 14614
rect 409306 14378 409542 14614
rect 408986 14058 409222 14294
rect 409306 14058 409542 14294
rect 408986 -3462 409222 -3226
rect 409306 -3462 409542 -3226
rect 408986 -3782 409222 -3546
rect 409306 -3782 409542 -3546
rect 412706 18098 412942 18334
rect 413026 18098 413262 18334
rect 412706 17778 412942 18014
rect 413026 17778 413262 18014
rect 412706 -4422 412942 -4186
rect 413026 -4422 413262 -4186
rect 412706 -4742 412942 -4506
rect 413026 -4742 413262 -4506
rect 416426 21818 416662 22054
rect 416746 21818 416982 22054
rect 416426 21498 416662 21734
rect 416746 21498 416982 21734
rect 416426 -5382 416662 -5146
rect 416746 -5382 416982 -5146
rect 416426 -5702 416662 -5466
rect 416746 -5702 416982 -5466
rect 420146 25538 420382 25774
rect 420466 25538 420702 25774
rect 420146 25218 420382 25454
rect 420466 25218 420702 25454
rect 420146 -6342 420382 -6106
rect 420466 -6342 420702 -6106
rect 420146 -6662 420382 -6426
rect 420466 -6662 420702 -6426
rect 433210 42938 433446 43174
rect 433210 42618 433446 42854
rect 423866 29258 424102 29494
rect 424186 29258 424422 29494
rect 423866 28938 424102 29174
rect 424186 28938 424422 29174
rect 423866 -7302 424102 -7066
rect 424186 -7302 424422 -7066
rect 423866 -7622 424102 -7386
rect 424186 -7622 424422 -7386
rect 433826 39218 434062 39454
rect 434146 39218 434382 39454
rect 433826 38898 434062 39134
rect 434146 38898 434382 39134
rect 433826 3218 434062 3454
rect 434146 3218 434382 3454
rect 433826 2898 434062 3134
rect 434146 2898 434382 3134
rect 433826 -582 434062 -346
rect 434146 -582 434382 -346
rect 433826 -902 434062 -666
rect 434146 -902 434382 -666
rect 437546 6938 437782 7174
rect 437866 6938 438102 7174
rect 437546 6618 437782 6854
rect 437866 6618 438102 6854
rect 437546 -1542 437782 -1306
rect 437866 -1542 438102 -1306
rect 437546 -1862 437782 -1626
rect 437866 -1862 438102 -1626
rect 441266 10658 441502 10894
rect 441586 10658 441822 10894
rect 441266 10338 441502 10574
rect 441586 10338 441822 10574
rect 441266 -2502 441502 -2266
rect 441586 -2502 441822 -2266
rect 441266 -2822 441502 -2586
rect 441586 -2822 441822 -2586
rect 444986 14378 445222 14614
rect 445306 14378 445542 14614
rect 444986 14058 445222 14294
rect 445306 14058 445542 14294
rect 444986 -3462 445222 -3226
rect 445306 -3462 445542 -3226
rect 444986 -3782 445222 -3546
rect 445306 -3782 445542 -3546
rect 448706 18098 448942 18334
rect 449026 18098 449262 18334
rect 448706 17778 448942 18014
rect 449026 17778 449262 18014
rect 448706 -4422 448942 -4186
rect 449026 -4422 449262 -4186
rect 448706 -4742 448942 -4506
rect 449026 -4742 449262 -4506
rect 452426 21818 452662 22054
rect 452746 21818 452982 22054
rect 452426 21498 452662 21734
rect 452746 21498 452982 21734
rect 452426 -5382 452662 -5146
rect 452746 -5382 452982 -5146
rect 452426 -5702 452662 -5466
rect 452746 -5702 452982 -5466
rect 456146 25538 456382 25774
rect 456466 25538 456702 25774
rect 456146 25218 456382 25454
rect 456466 25218 456702 25454
rect 456146 -6342 456382 -6106
rect 456466 -6342 456702 -6106
rect 456146 -6662 456382 -6426
rect 456466 -6662 456702 -6426
rect 463930 42938 464166 43174
rect 463930 42618 464166 42854
rect 459866 29258 460102 29494
rect 460186 29258 460422 29494
rect 459866 28938 460102 29174
rect 460186 28938 460422 29174
rect 459866 -7302 460102 -7066
rect 460186 -7302 460422 -7066
rect 459866 -7622 460102 -7386
rect 460186 -7622 460422 -7386
rect 469826 39218 470062 39454
rect 470146 39218 470382 39454
rect 469826 38898 470062 39134
rect 470146 38898 470382 39134
rect 469826 3218 470062 3454
rect 470146 3218 470382 3454
rect 469826 2898 470062 3134
rect 470146 2898 470382 3134
rect 469826 -582 470062 -346
rect 470146 -582 470382 -346
rect 469826 -902 470062 -666
rect 470146 -902 470382 -666
rect 473546 6938 473782 7174
rect 473866 6938 474102 7174
rect 473546 6618 473782 6854
rect 473866 6618 474102 6854
rect 473546 -1542 473782 -1306
rect 473866 -1542 474102 -1306
rect 473546 -1862 473782 -1626
rect 473866 -1862 474102 -1626
rect 477266 10658 477502 10894
rect 477586 10658 477822 10894
rect 477266 10338 477502 10574
rect 477586 10338 477822 10574
rect 477266 -2502 477502 -2266
rect 477586 -2502 477822 -2266
rect 477266 -2822 477502 -2586
rect 477586 -2822 477822 -2586
rect 480986 14378 481222 14614
rect 481306 14378 481542 14614
rect 480986 14058 481222 14294
rect 481306 14058 481542 14294
rect 480986 -3462 481222 -3226
rect 481306 -3462 481542 -3226
rect 480986 -3782 481222 -3546
rect 481306 -3782 481542 -3546
rect 484706 18098 484942 18334
rect 485026 18098 485262 18334
rect 484706 17778 484942 18014
rect 485026 17778 485262 18014
rect 484706 -4422 484942 -4186
rect 485026 -4422 485262 -4186
rect 484706 -4742 484942 -4506
rect 485026 -4742 485262 -4506
rect 488426 21818 488662 22054
rect 488746 21818 488982 22054
rect 488426 21498 488662 21734
rect 488746 21498 488982 21734
rect 488426 -5382 488662 -5146
rect 488746 -5382 488982 -5146
rect 488426 -5702 488662 -5466
rect 488746 -5702 488982 -5466
rect 494650 42938 494886 43174
rect 494650 42618 494886 42854
rect 492146 25538 492382 25774
rect 492466 25538 492702 25774
rect 492146 25218 492382 25454
rect 492466 25218 492702 25454
rect 492146 -6342 492382 -6106
rect 492466 -6342 492702 -6106
rect 492146 -6662 492382 -6426
rect 492466 -6662 492702 -6426
rect 495866 29258 496102 29494
rect 496186 29258 496422 29494
rect 495866 28938 496102 29174
rect 496186 28938 496422 29174
rect 495866 -7302 496102 -7066
rect 496186 -7302 496422 -7066
rect 495866 -7622 496102 -7386
rect 496186 -7622 496422 -7386
rect 505826 39218 506062 39454
rect 506146 39218 506382 39454
rect 505826 38898 506062 39134
rect 506146 38898 506382 39134
rect 505826 3218 506062 3454
rect 506146 3218 506382 3454
rect 505826 2898 506062 3134
rect 506146 2898 506382 3134
rect 505826 -582 506062 -346
rect 506146 -582 506382 -346
rect 505826 -902 506062 -666
rect 506146 -902 506382 -666
rect 509546 6938 509782 7174
rect 509866 6938 510102 7174
rect 509546 6618 509782 6854
rect 509866 6618 510102 6854
rect 509546 -1542 509782 -1306
rect 509866 -1542 510102 -1306
rect 509546 -1862 509782 -1626
rect 509866 -1862 510102 -1626
rect 513266 10658 513502 10894
rect 513586 10658 513822 10894
rect 513266 10338 513502 10574
rect 513586 10338 513822 10574
rect 513266 -2502 513502 -2266
rect 513586 -2502 513822 -2266
rect 513266 -2822 513502 -2586
rect 513586 -2822 513822 -2586
rect 516986 14378 517222 14614
rect 517306 14378 517542 14614
rect 516986 14058 517222 14294
rect 517306 14058 517542 14294
rect 516986 -3462 517222 -3226
rect 517306 -3462 517542 -3226
rect 516986 -3782 517222 -3546
rect 517306 -3782 517542 -3546
rect 520706 18098 520942 18334
rect 521026 18098 521262 18334
rect 520706 17778 520942 18014
rect 521026 17778 521262 18014
rect 520706 -4422 520942 -4186
rect 521026 -4422 521262 -4186
rect 520706 -4742 520942 -4506
rect 521026 -4742 521262 -4506
rect 525370 42938 525606 43174
rect 525370 42618 525606 42854
rect 524426 21818 524662 22054
rect 524746 21818 524982 22054
rect 524426 21498 524662 21734
rect 524746 21498 524982 21734
rect 524426 -5382 524662 -5146
rect 524746 -5382 524982 -5146
rect 524426 -5702 524662 -5466
rect 524746 -5702 524982 -5466
rect 528146 25538 528382 25774
rect 528466 25538 528702 25774
rect 528146 25218 528382 25454
rect 528466 25218 528702 25454
rect 528146 -6342 528382 -6106
rect 528466 -6342 528702 -6106
rect 528146 -6662 528382 -6426
rect 528466 -6662 528702 -6426
rect 531866 29258 532102 29494
rect 532186 29258 532422 29494
rect 531866 28938 532102 29174
rect 532186 28938 532422 29174
rect 531866 -7302 532102 -7066
rect 532186 -7302 532422 -7066
rect 531866 -7622 532102 -7386
rect 532186 -7622 532422 -7386
rect 541826 39218 542062 39454
rect 542146 39218 542382 39454
rect 541826 38898 542062 39134
rect 542146 38898 542382 39134
rect 541826 3218 542062 3454
rect 542146 3218 542382 3454
rect 541826 2898 542062 3134
rect 542146 2898 542382 3134
rect 541826 -582 542062 -346
rect 542146 -582 542382 -346
rect 541826 -902 542062 -666
rect 542146 -902 542382 -666
rect 545546 6938 545782 7174
rect 545866 6938 546102 7174
rect 545546 6618 545782 6854
rect 545866 6618 546102 6854
rect 545546 -1542 545782 -1306
rect 545866 -1542 546102 -1306
rect 545546 -1862 545782 -1626
rect 545866 -1862 546102 -1626
rect 549266 10658 549502 10894
rect 549586 10658 549822 10894
rect 549266 10338 549502 10574
rect 549586 10338 549822 10574
rect 549266 -2502 549502 -2266
rect 549586 -2502 549822 -2266
rect 549266 -2822 549502 -2586
rect 549586 -2822 549822 -2586
rect 552986 14378 553222 14614
rect 553306 14378 553542 14614
rect 552986 14058 553222 14294
rect 553306 14058 553542 14294
rect 552986 -3462 553222 -3226
rect 553306 -3462 553542 -3226
rect 552986 -3782 553222 -3546
rect 553306 -3782 553542 -3546
rect 556706 708442 556942 708678
rect 557026 708442 557262 708678
rect 556706 708122 556942 708358
rect 557026 708122 557262 708358
rect 556706 666098 556942 666334
rect 557026 666098 557262 666334
rect 556706 665778 556942 666014
rect 557026 665778 557262 666014
rect 556706 630098 556942 630334
rect 557026 630098 557262 630334
rect 556706 629778 556942 630014
rect 557026 629778 557262 630014
rect 556706 594098 556942 594334
rect 557026 594098 557262 594334
rect 556706 593778 556942 594014
rect 557026 593778 557262 594014
rect 556706 558098 556942 558334
rect 557026 558098 557262 558334
rect 556706 557778 556942 558014
rect 557026 557778 557262 558014
rect 556706 522098 556942 522334
rect 557026 522098 557262 522334
rect 556706 521778 556942 522014
rect 557026 521778 557262 522014
rect 556706 486098 556942 486334
rect 557026 486098 557262 486334
rect 556706 485778 556942 486014
rect 557026 485778 557262 486014
rect 556706 450098 556942 450334
rect 557026 450098 557262 450334
rect 556706 449778 556942 450014
rect 557026 449778 557262 450014
rect 556706 414098 556942 414334
rect 557026 414098 557262 414334
rect 556706 413778 556942 414014
rect 557026 413778 557262 414014
rect 556706 378098 556942 378334
rect 557026 378098 557262 378334
rect 556706 377778 556942 378014
rect 557026 377778 557262 378014
rect 556706 342098 556942 342334
rect 557026 342098 557262 342334
rect 556706 341778 556942 342014
rect 557026 341778 557262 342014
rect 556706 306098 556942 306334
rect 557026 306098 557262 306334
rect 556706 305778 556942 306014
rect 557026 305778 557262 306014
rect 556706 270098 556942 270334
rect 557026 270098 557262 270334
rect 556706 269778 556942 270014
rect 557026 269778 557262 270014
rect 556706 234098 556942 234334
rect 557026 234098 557262 234334
rect 556706 233778 556942 234014
rect 557026 233778 557262 234014
rect 556706 198098 556942 198334
rect 557026 198098 557262 198334
rect 556706 197778 556942 198014
rect 557026 197778 557262 198014
rect 556706 162098 556942 162334
rect 557026 162098 557262 162334
rect 556706 161778 556942 162014
rect 557026 161778 557262 162014
rect 556706 126098 556942 126334
rect 557026 126098 557262 126334
rect 556706 125778 556942 126014
rect 557026 125778 557262 126014
rect 556706 90098 556942 90334
rect 557026 90098 557262 90334
rect 556706 89778 556942 90014
rect 557026 89778 557262 90014
rect 556706 54098 556942 54334
rect 557026 54098 557262 54334
rect 556706 53778 556942 54014
rect 557026 53778 557262 54014
rect 556706 18098 556942 18334
rect 557026 18098 557262 18334
rect 556706 17778 556942 18014
rect 557026 17778 557262 18014
rect 556706 -4422 556942 -4186
rect 557026 -4422 557262 -4186
rect 556706 -4742 556942 -4506
rect 557026 -4742 557262 -4506
rect 560426 709402 560662 709638
rect 560746 709402 560982 709638
rect 560426 709082 560662 709318
rect 560746 709082 560982 709318
rect 560426 669818 560662 670054
rect 560746 669818 560982 670054
rect 560426 669498 560662 669734
rect 560746 669498 560982 669734
rect 560426 633818 560662 634054
rect 560746 633818 560982 634054
rect 560426 633498 560662 633734
rect 560746 633498 560982 633734
rect 560426 597818 560662 598054
rect 560746 597818 560982 598054
rect 560426 597498 560662 597734
rect 560746 597498 560982 597734
rect 560426 561818 560662 562054
rect 560746 561818 560982 562054
rect 560426 561498 560662 561734
rect 560746 561498 560982 561734
rect 560426 525818 560662 526054
rect 560746 525818 560982 526054
rect 560426 525498 560662 525734
rect 560746 525498 560982 525734
rect 560426 489818 560662 490054
rect 560746 489818 560982 490054
rect 560426 489498 560662 489734
rect 560746 489498 560982 489734
rect 560426 453818 560662 454054
rect 560746 453818 560982 454054
rect 560426 453498 560662 453734
rect 560746 453498 560982 453734
rect 560426 417818 560662 418054
rect 560746 417818 560982 418054
rect 560426 417498 560662 417734
rect 560746 417498 560982 417734
rect 560426 381818 560662 382054
rect 560746 381818 560982 382054
rect 560426 381498 560662 381734
rect 560746 381498 560982 381734
rect 560426 345818 560662 346054
rect 560746 345818 560982 346054
rect 560426 345498 560662 345734
rect 560746 345498 560982 345734
rect 560426 309818 560662 310054
rect 560746 309818 560982 310054
rect 560426 309498 560662 309734
rect 560746 309498 560982 309734
rect 560426 273818 560662 274054
rect 560746 273818 560982 274054
rect 560426 273498 560662 273734
rect 560746 273498 560982 273734
rect 560426 237818 560662 238054
rect 560746 237818 560982 238054
rect 560426 237498 560662 237734
rect 560746 237498 560982 237734
rect 560426 201818 560662 202054
rect 560746 201818 560982 202054
rect 560426 201498 560662 201734
rect 560746 201498 560982 201734
rect 560426 165818 560662 166054
rect 560746 165818 560982 166054
rect 560426 165498 560662 165734
rect 560746 165498 560982 165734
rect 560426 129818 560662 130054
rect 560746 129818 560982 130054
rect 560426 129498 560662 129734
rect 560746 129498 560982 129734
rect 560426 93818 560662 94054
rect 560746 93818 560982 94054
rect 560426 93498 560662 93734
rect 560746 93498 560982 93734
rect 560426 57818 560662 58054
rect 560746 57818 560982 58054
rect 560426 57498 560662 57734
rect 560746 57498 560982 57734
rect 560426 21818 560662 22054
rect 560746 21818 560982 22054
rect 560426 21498 560662 21734
rect 560746 21498 560982 21734
rect 560426 -5382 560662 -5146
rect 560746 -5382 560982 -5146
rect 560426 -5702 560662 -5466
rect 560746 -5702 560982 -5466
rect 564146 710362 564382 710598
rect 564466 710362 564702 710598
rect 564146 710042 564382 710278
rect 564466 710042 564702 710278
rect 564146 673538 564382 673774
rect 564466 673538 564702 673774
rect 564146 673218 564382 673454
rect 564466 673218 564702 673454
rect 564146 637538 564382 637774
rect 564466 637538 564702 637774
rect 564146 637218 564382 637454
rect 564466 637218 564702 637454
rect 567866 711322 568102 711558
rect 568186 711322 568422 711558
rect 567866 711002 568102 711238
rect 568186 711002 568422 711238
rect 567866 677258 568102 677494
rect 568186 677258 568422 677494
rect 567866 676938 568102 677174
rect 568186 676938 568422 677174
rect 567866 641258 568102 641494
rect 568186 641258 568422 641494
rect 567866 640938 568102 641174
rect 568186 640938 568422 641174
rect 565050 615218 565286 615454
rect 565050 614898 565286 615134
rect 564146 601538 564382 601774
rect 564466 601538 564702 601774
rect 564146 601218 564382 601454
rect 564466 601218 564702 601454
rect 567866 605258 568102 605494
rect 568186 605258 568422 605494
rect 567866 604938 568102 605174
rect 568186 604938 568422 605174
rect 565050 579218 565286 579454
rect 565050 578898 565286 579134
rect 564146 565538 564382 565774
rect 564466 565538 564702 565774
rect 564146 565218 564382 565454
rect 564466 565218 564702 565454
rect 567866 569258 568102 569494
rect 568186 569258 568422 569494
rect 567866 568938 568102 569174
rect 568186 568938 568422 569174
rect 565050 543218 565286 543454
rect 565050 542898 565286 543134
rect 564146 529538 564382 529774
rect 564466 529538 564702 529774
rect 564146 529218 564382 529454
rect 564466 529218 564702 529454
rect 564146 493538 564382 493774
rect 564466 493538 564702 493774
rect 564146 493218 564382 493454
rect 564466 493218 564702 493454
rect 567866 533258 568102 533494
rect 568186 533258 568422 533494
rect 567866 532938 568102 533174
rect 568186 532938 568422 533174
rect 567866 497258 568102 497494
rect 568186 497258 568422 497494
rect 567866 496938 568102 497174
rect 568186 496938 568422 497174
rect 565050 471218 565286 471454
rect 565050 470898 565286 471134
rect 564146 457538 564382 457774
rect 564466 457538 564702 457774
rect 564146 457218 564382 457454
rect 564466 457218 564702 457454
rect 567866 461258 568102 461494
rect 568186 461258 568422 461494
rect 567866 460938 568102 461174
rect 568186 460938 568422 461174
rect 565050 435218 565286 435454
rect 565050 434898 565286 435134
rect 564146 421538 564382 421774
rect 564466 421538 564702 421774
rect 564146 421218 564382 421454
rect 564466 421218 564702 421454
rect 567866 425258 568102 425494
rect 568186 425258 568422 425494
rect 567866 424938 568102 425174
rect 568186 424938 568422 425174
rect 565050 399218 565286 399454
rect 565050 398898 565286 399134
rect 564146 385538 564382 385774
rect 564466 385538 564702 385774
rect 564146 385218 564382 385454
rect 564466 385218 564702 385454
rect 564146 349538 564382 349774
rect 564466 349538 564702 349774
rect 564146 349218 564382 349454
rect 564466 349218 564702 349454
rect 564146 313538 564382 313774
rect 564466 313538 564702 313774
rect 564146 313218 564382 313454
rect 564466 313218 564702 313454
rect 564146 277538 564382 277774
rect 564466 277538 564702 277774
rect 564146 277218 564382 277454
rect 564466 277218 564702 277454
rect 564146 241538 564382 241774
rect 564466 241538 564702 241774
rect 564146 241218 564382 241454
rect 564466 241218 564702 241454
rect 564146 205538 564382 205774
rect 564466 205538 564702 205774
rect 564146 205218 564382 205454
rect 564466 205218 564702 205454
rect 564146 169538 564382 169774
rect 564466 169538 564702 169774
rect 564146 169218 564382 169454
rect 564466 169218 564702 169454
rect 564146 133538 564382 133774
rect 564466 133538 564702 133774
rect 564146 133218 564382 133454
rect 564466 133218 564702 133454
rect 564146 97538 564382 97774
rect 564466 97538 564702 97774
rect 564146 97218 564382 97454
rect 564466 97218 564702 97454
rect 564146 61538 564382 61774
rect 564466 61538 564702 61774
rect 564146 61218 564382 61454
rect 564466 61218 564702 61454
rect 564146 25538 564382 25774
rect 564466 25538 564702 25774
rect 564146 25218 564382 25454
rect 564466 25218 564702 25454
rect 564146 -6342 564382 -6106
rect 564466 -6342 564702 -6106
rect 564146 -6662 564382 -6426
rect 564466 -6662 564702 -6426
rect 567866 389258 568102 389494
rect 568186 389258 568422 389494
rect 567866 388938 568102 389174
rect 568186 388938 568422 389174
rect 567866 353258 568102 353494
rect 568186 353258 568422 353494
rect 567866 352938 568102 353174
rect 568186 352938 568422 353174
rect 567866 317258 568102 317494
rect 568186 317258 568422 317494
rect 567866 316938 568102 317174
rect 568186 316938 568422 317174
rect 567866 281258 568102 281494
rect 568186 281258 568422 281494
rect 567866 280938 568102 281174
rect 568186 280938 568422 281174
rect 567866 245258 568102 245494
rect 568186 245258 568422 245494
rect 567866 244938 568102 245174
rect 568186 244938 568422 245174
rect 567866 209258 568102 209494
rect 568186 209258 568422 209494
rect 567866 208938 568102 209174
rect 568186 208938 568422 209174
rect 567866 173258 568102 173494
rect 568186 173258 568422 173494
rect 567866 172938 568102 173174
rect 568186 172938 568422 173174
rect 567866 137258 568102 137494
rect 568186 137258 568422 137494
rect 567866 136938 568102 137174
rect 568186 136938 568422 137174
rect 567866 101258 568102 101494
rect 568186 101258 568422 101494
rect 567866 100938 568102 101174
rect 568186 100938 568422 101174
rect 567866 65258 568102 65494
rect 568186 65258 568422 65494
rect 567866 64938 568102 65174
rect 568186 64938 568422 65174
rect 567866 29258 568102 29494
rect 568186 29258 568422 29494
rect 567866 28938 568102 29174
rect 568186 28938 568422 29174
rect 567866 -7302 568102 -7066
rect 568186 -7302 568422 -7066
rect 567866 -7622 568102 -7386
rect 568186 -7622 568422 -7386
rect 577826 704602 578062 704838
rect 578146 704602 578382 704838
rect 577826 704282 578062 704518
rect 578146 704282 578382 704518
rect 577826 687218 578062 687454
rect 578146 687218 578382 687454
rect 577826 686898 578062 687134
rect 578146 686898 578382 687134
rect 577826 651218 578062 651454
rect 578146 651218 578382 651454
rect 577826 650898 578062 651134
rect 578146 650898 578382 651134
rect 577826 615218 578062 615454
rect 578146 615218 578382 615454
rect 577826 614898 578062 615134
rect 578146 614898 578382 615134
rect 577826 579218 578062 579454
rect 578146 579218 578382 579454
rect 577826 578898 578062 579134
rect 578146 578898 578382 579134
rect 577826 543218 578062 543454
rect 578146 543218 578382 543454
rect 577826 542898 578062 543134
rect 578146 542898 578382 543134
rect 577826 507218 578062 507454
rect 578146 507218 578382 507454
rect 577826 506898 578062 507134
rect 578146 506898 578382 507134
rect 577826 471218 578062 471454
rect 578146 471218 578382 471454
rect 577826 470898 578062 471134
rect 578146 470898 578382 471134
rect 577826 435218 578062 435454
rect 578146 435218 578382 435454
rect 577826 434898 578062 435134
rect 578146 434898 578382 435134
rect 577826 399218 578062 399454
rect 578146 399218 578382 399454
rect 577826 398898 578062 399134
rect 578146 398898 578382 399134
rect 577826 363218 578062 363454
rect 578146 363218 578382 363454
rect 577826 362898 578062 363134
rect 578146 362898 578382 363134
rect 577826 327218 578062 327454
rect 578146 327218 578382 327454
rect 577826 326898 578062 327134
rect 578146 326898 578382 327134
rect 577826 291218 578062 291454
rect 578146 291218 578382 291454
rect 577826 290898 578062 291134
rect 578146 290898 578382 291134
rect 577826 255218 578062 255454
rect 578146 255218 578382 255454
rect 577826 254898 578062 255134
rect 578146 254898 578382 255134
rect 577826 219218 578062 219454
rect 578146 219218 578382 219454
rect 577826 218898 578062 219134
rect 578146 218898 578382 219134
rect 577826 183218 578062 183454
rect 578146 183218 578382 183454
rect 577826 182898 578062 183134
rect 578146 182898 578382 183134
rect 577826 147218 578062 147454
rect 578146 147218 578382 147454
rect 577826 146898 578062 147134
rect 578146 146898 578382 147134
rect 577826 111218 578062 111454
rect 578146 111218 578382 111454
rect 577826 110898 578062 111134
rect 578146 110898 578382 111134
rect 577826 75218 578062 75454
rect 578146 75218 578382 75454
rect 577826 74898 578062 75134
rect 578146 74898 578382 75134
rect 577826 39218 578062 39454
rect 578146 39218 578382 39454
rect 577826 38898 578062 39134
rect 578146 38898 578382 39134
rect 577826 3218 578062 3454
rect 578146 3218 578382 3454
rect 577826 2898 578062 3134
rect 578146 2898 578382 3134
rect 577826 -582 578062 -346
rect 578146 -582 578382 -346
rect 577826 -902 578062 -666
rect 578146 -902 578382 -666
rect 592062 711322 592298 711558
rect 592382 711322 592618 711558
rect 592062 711002 592298 711238
rect 592382 711002 592618 711238
rect 591102 710362 591338 710598
rect 591422 710362 591658 710598
rect 591102 710042 591338 710278
rect 591422 710042 591658 710278
rect 590142 709402 590378 709638
rect 590462 709402 590698 709638
rect 590142 709082 590378 709318
rect 590462 709082 590698 709318
rect 589182 708442 589418 708678
rect 589502 708442 589738 708678
rect 589182 708122 589418 708358
rect 589502 708122 589738 708358
rect 588222 707482 588458 707718
rect 588542 707482 588778 707718
rect 588222 707162 588458 707398
rect 588542 707162 588778 707398
rect 587262 706522 587498 706758
rect 587582 706522 587818 706758
rect 587262 706202 587498 706438
rect 587582 706202 587818 706438
rect 581546 705562 581782 705798
rect 581866 705562 582102 705798
rect 581546 705242 581782 705478
rect 581866 705242 582102 705478
rect 586302 705562 586538 705798
rect 586622 705562 586858 705798
rect 586302 705242 586538 705478
rect 586622 705242 586858 705478
rect 581546 690938 581782 691174
rect 581866 690938 582102 691174
rect 581546 690618 581782 690854
rect 581866 690618 582102 690854
rect 581546 654938 581782 655174
rect 581866 654938 582102 655174
rect 581546 654618 581782 654854
rect 581866 654618 582102 654854
rect 581546 618938 581782 619174
rect 581866 618938 582102 619174
rect 581546 618618 581782 618854
rect 581866 618618 582102 618854
rect 581546 582938 581782 583174
rect 581866 582938 582102 583174
rect 581546 582618 581782 582854
rect 581866 582618 582102 582854
rect 581546 546938 581782 547174
rect 581866 546938 582102 547174
rect 581546 546618 581782 546854
rect 581866 546618 582102 546854
rect 581546 510938 581782 511174
rect 581866 510938 582102 511174
rect 581546 510618 581782 510854
rect 581866 510618 582102 510854
rect 581546 474938 581782 475174
rect 581866 474938 582102 475174
rect 581546 474618 581782 474854
rect 581866 474618 582102 474854
rect 581546 438938 581782 439174
rect 581866 438938 582102 439174
rect 581546 438618 581782 438854
rect 581866 438618 582102 438854
rect 581546 402938 581782 403174
rect 581866 402938 582102 403174
rect 581546 402618 581782 402854
rect 581866 402618 582102 402854
rect 581546 366938 581782 367174
rect 581866 366938 582102 367174
rect 581546 366618 581782 366854
rect 581866 366618 582102 366854
rect 581546 330938 581782 331174
rect 581866 330938 582102 331174
rect 581546 330618 581782 330854
rect 581866 330618 582102 330854
rect 581546 294938 581782 295174
rect 581866 294938 582102 295174
rect 581546 294618 581782 294854
rect 581866 294618 582102 294854
rect 581546 258938 581782 259174
rect 581866 258938 582102 259174
rect 581546 258618 581782 258854
rect 581866 258618 582102 258854
rect 581546 222938 581782 223174
rect 581866 222938 582102 223174
rect 581546 222618 581782 222854
rect 581866 222618 582102 222854
rect 581546 186938 581782 187174
rect 581866 186938 582102 187174
rect 581546 186618 581782 186854
rect 581866 186618 582102 186854
rect 581546 150938 581782 151174
rect 581866 150938 582102 151174
rect 581546 150618 581782 150854
rect 581866 150618 582102 150854
rect 581546 114938 581782 115174
rect 581866 114938 582102 115174
rect 581546 114618 581782 114854
rect 581866 114618 582102 114854
rect 581546 78938 581782 79174
rect 581866 78938 582102 79174
rect 581546 78618 581782 78854
rect 581866 78618 582102 78854
rect 581546 42938 581782 43174
rect 581866 42938 582102 43174
rect 581546 42618 581782 42854
rect 581866 42618 582102 42854
rect 581546 6938 581782 7174
rect 581866 6938 582102 7174
rect 581546 6618 581782 6854
rect 581866 6618 582102 6854
rect 585342 704602 585578 704838
rect 585662 704602 585898 704838
rect 585342 704282 585578 704518
rect 585662 704282 585898 704518
rect 585342 687218 585578 687454
rect 585662 687218 585898 687454
rect 585342 686898 585578 687134
rect 585662 686898 585898 687134
rect 585342 651218 585578 651454
rect 585662 651218 585898 651454
rect 585342 650898 585578 651134
rect 585662 650898 585898 651134
rect 585342 615218 585578 615454
rect 585662 615218 585898 615454
rect 585342 614898 585578 615134
rect 585662 614898 585898 615134
rect 585342 579218 585578 579454
rect 585662 579218 585898 579454
rect 585342 578898 585578 579134
rect 585662 578898 585898 579134
rect 585342 543218 585578 543454
rect 585662 543218 585898 543454
rect 585342 542898 585578 543134
rect 585662 542898 585898 543134
rect 585342 507218 585578 507454
rect 585662 507218 585898 507454
rect 585342 506898 585578 507134
rect 585662 506898 585898 507134
rect 585342 471218 585578 471454
rect 585662 471218 585898 471454
rect 585342 470898 585578 471134
rect 585662 470898 585898 471134
rect 585342 435218 585578 435454
rect 585662 435218 585898 435454
rect 585342 434898 585578 435134
rect 585662 434898 585898 435134
rect 585342 399218 585578 399454
rect 585662 399218 585898 399454
rect 585342 398898 585578 399134
rect 585662 398898 585898 399134
rect 585342 363218 585578 363454
rect 585662 363218 585898 363454
rect 585342 362898 585578 363134
rect 585662 362898 585898 363134
rect 585342 327218 585578 327454
rect 585662 327218 585898 327454
rect 585342 326898 585578 327134
rect 585662 326898 585898 327134
rect 585342 291218 585578 291454
rect 585662 291218 585898 291454
rect 585342 290898 585578 291134
rect 585662 290898 585898 291134
rect 585342 255218 585578 255454
rect 585662 255218 585898 255454
rect 585342 254898 585578 255134
rect 585662 254898 585898 255134
rect 585342 219218 585578 219454
rect 585662 219218 585898 219454
rect 585342 218898 585578 219134
rect 585662 218898 585898 219134
rect 585342 183218 585578 183454
rect 585662 183218 585898 183454
rect 585342 182898 585578 183134
rect 585662 182898 585898 183134
rect 585342 147218 585578 147454
rect 585662 147218 585898 147454
rect 585342 146898 585578 147134
rect 585662 146898 585898 147134
rect 585342 111218 585578 111454
rect 585662 111218 585898 111454
rect 585342 110898 585578 111134
rect 585662 110898 585898 111134
rect 585342 75218 585578 75454
rect 585662 75218 585898 75454
rect 585342 74898 585578 75134
rect 585662 74898 585898 75134
rect 585342 39218 585578 39454
rect 585662 39218 585898 39454
rect 585342 38898 585578 39134
rect 585662 38898 585898 39134
rect 585342 3218 585578 3454
rect 585662 3218 585898 3454
rect 585342 2898 585578 3134
rect 585662 2898 585898 3134
rect 585342 -582 585578 -346
rect 585662 -582 585898 -346
rect 585342 -902 585578 -666
rect 585662 -902 585898 -666
rect 586302 690938 586538 691174
rect 586622 690938 586858 691174
rect 586302 690618 586538 690854
rect 586622 690618 586858 690854
rect 586302 654938 586538 655174
rect 586622 654938 586858 655174
rect 586302 654618 586538 654854
rect 586622 654618 586858 654854
rect 586302 618938 586538 619174
rect 586622 618938 586858 619174
rect 586302 618618 586538 618854
rect 586622 618618 586858 618854
rect 586302 582938 586538 583174
rect 586622 582938 586858 583174
rect 586302 582618 586538 582854
rect 586622 582618 586858 582854
rect 586302 546938 586538 547174
rect 586622 546938 586858 547174
rect 586302 546618 586538 546854
rect 586622 546618 586858 546854
rect 586302 510938 586538 511174
rect 586622 510938 586858 511174
rect 586302 510618 586538 510854
rect 586622 510618 586858 510854
rect 586302 474938 586538 475174
rect 586622 474938 586858 475174
rect 586302 474618 586538 474854
rect 586622 474618 586858 474854
rect 586302 438938 586538 439174
rect 586622 438938 586858 439174
rect 586302 438618 586538 438854
rect 586622 438618 586858 438854
rect 586302 402938 586538 403174
rect 586622 402938 586858 403174
rect 586302 402618 586538 402854
rect 586622 402618 586858 402854
rect 586302 366938 586538 367174
rect 586622 366938 586858 367174
rect 586302 366618 586538 366854
rect 586622 366618 586858 366854
rect 586302 330938 586538 331174
rect 586622 330938 586858 331174
rect 586302 330618 586538 330854
rect 586622 330618 586858 330854
rect 586302 294938 586538 295174
rect 586622 294938 586858 295174
rect 586302 294618 586538 294854
rect 586622 294618 586858 294854
rect 586302 258938 586538 259174
rect 586622 258938 586858 259174
rect 586302 258618 586538 258854
rect 586622 258618 586858 258854
rect 586302 222938 586538 223174
rect 586622 222938 586858 223174
rect 586302 222618 586538 222854
rect 586622 222618 586858 222854
rect 586302 186938 586538 187174
rect 586622 186938 586858 187174
rect 586302 186618 586538 186854
rect 586622 186618 586858 186854
rect 586302 150938 586538 151174
rect 586622 150938 586858 151174
rect 586302 150618 586538 150854
rect 586622 150618 586858 150854
rect 586302 114938 586538 115174
rect 586622 114938 586858 115174
rect 586302 114618 586538 114854
rect 586622 114618 586858 114854
rect 586302 78938 586538 79174
rect 586622 78938 586858 79174
rect 586302 78618 586538 78854
rect 586622 78618 586858 78854
rect 586302 42938 586538 43174
rect 586622 42938 586858 43174
rect 586302 42618 586538 42854
rect 586622 42618 586858 42854
rect 586302 6938 586538 7174
rect 586622 6938 586858 7174
rect 586302 6618 586538 6854
rect 586622 6618 586858 6854
rect 581546 -1542 581782 -1306
rect 581866 -1542 582102 -1306
rect 581546 -1862 581782 -1626
rect 581866 -1862 582102 -1626
rect 586302 -1542 586538 -1306
rect 586622 -1542 586858 -1306
rect 586302 -1862 586538 -1626
rect 586622 -1862 586858 -1626
rect 587262 694658 587498 694894
rect 587582 694658 587818 694894
rect 587262 694338 587498 694574
rect 587582 694338 587818 694574
rect 587262 658658 587498 658894
rect 587582 658658 587818 658894
rect 587262 658338 587498 658574
rect 587582 658338 587818 658574
rect 587262 622658 587498 622894
rect 587582 622658 587818 622894
rect 587262 622338 587498 622574
rect 587582 622338 587818 622574
rect 587262 586658 587498 586894
rect 587582 586658 587818 586894
rect 587262 586338 587498 586574
rect 587582 586338 587818 586574
rect 587262 550658 587498 550894
rect 587582 550658 587818 550894
rect 587262 550338 587498 550574
rect 587582 550338 587818 550574
rect 587262 514658 587498 514894
rect 587582 514658 587818 514894
rect 587262 514338 587498 514574
rect 587582 514338 587818 514574
rect 587262 478658 587498 478894
rect 587582 478658 587818 478894
rect 587262 478338 587498 478574
rect 587582 478338 587818 478574
rect 587262 442658 587498 442894
rect 587582 442658 587818 442894
rect 587262 442338 587498 442574
rect 587582 442338 587818 442574
rect 587262 406658 587498 406894
rect 587582 406658 587818 406894
rect 587262 406338 587498 406574
rect 587582 406338 587818 406574
rect 587262 370658 587498 370894
rect 587582 370658 587818 370894
rect 587262 370338 587498 370574
rect 587582 370338 587818 370574
rect 587262 334658 587498 334894
rect 587582 334658 587818 334894
rect 587262 334338 587498 334574
rect 587582 334338 587818 334574
rect 587262 298658 587498 298894
rect 587582 298658 587818 298894
rect 587262 298338 587498 298574
rect 587582 298338 587818 298574
rect 587262 262658 587498 262894
rect 587582 262658 587818 262894
rect 587262 262338 587498 262574
rect 587582 262338 587818 262574
rect 587262 226658 587498 226894
rect 587582 226658 587818 226894
rect 587262 226338 587498 226574
rect 587582 226338 587818 226574
rect 587262 190658 587498 190894
rect 587582 190658 587818 190894
rect 587262 190338 587498 190574
rect 587582 190338 587818 190574
rect 587262 154658 587498 154894
rect 587582 154658 587818 154894
rect 587262 154338 587498 154574
rect 587582 154338 587818 154574
rect 587262 118658 587498 118894
rect 587582 118658 587818 118894
rect 587262 118338 587498 118574
rect 587582 118338 587818 118574
rect 587262 82658 587498 82894
rect 587582 82658 587818 82894
rect 587262 82338 587498 82574
rect 587582 82338 587818 82574
rect 587262 46658 587498 46894
rect 587582 46658 587818 46894
rect 587262 46338 587498 46574
rect 587582 46338 587818 46574
rect 587262 10658 587498 10894
rect 587582 10658 587818 10894
rect 587262 10338 587498 10574
rect 587582 10338 587818 10574
rect 587262 -2502 587498 -2266
rect 587582 -2502 587818 -2266
rect 587262 -2822 587498 -2586
rect 587582 -2822 587818 -2586
rect 588222 698378 588458 698614
rect 588542 698378 588778 698614
rect 588222 698058 588458 698294
rect 588542 698058 588778 698294
rect 588222 662378 588458 662614
rect 588542 662378 588778 662614
rect 588222 662058 588458 662294
rect 588542 662058 588778 662294
rect 588222 626378 588458 626614
rect 588542 626378 588778 626614
rect 588222 626058 588458 626294
rect 588542 626058 588778 626294
rect 588222 590378 588458 590614
rect 588542 590378 588778 590614
rect 588222 590058 588458 590294
rect 588542 590058 588778 590294
rect 588222 554378 588458 554614
rect 588542 554378 588778 554614
rect 588222 554058 588458 554294
rect 588542 554058 588778 554294
rect 588222 518378 588458 518614
rect 588542 518378 588778 518614
rect 588222 518058 588458 518294
rect 588542 518058 588778 518294
rect 588222 482378 588458 482614
rect 588542 482378 588778 482614
rect 588222 482058 588458 482294
rect 588542 482058 588778 482294
rect 588222 446378 588458 446614
rect 588542 446378 588778 446614
rect 588222 446058 588458 446294
rect 588542 446058 588778 446294
rect 588222 410378 588458 410614
rect 588542 410378 588778 410614
rect 588222 410058 588458 410294
rect 588542 410058 588778 410294
rect 588222 374378 588458 374614
rect 588542 374378 588778 374614
rect 588222 374058 588458 374294
rect 588542 374058 588778 374294
rect 588222 338378 588458 338614
rect 588542 338378 588778 338614
rect 588222 338058 588458 338294
rect 588542 338058 588778 338294
rect 588222 302378 588458 302614
rect 588542 302378 588778 302614
rect 588222 302058 588458 302294
rect 588542 302058 588778 302294
rect 588222 266378 588458 266614
rect 588542 266378 588778 266614
rect 588222 266058 588458 266294
rect 588542 266058 588778 266294
rect 588222 230378 588458 230614
rect 588542 230378 588778 230614
rect 588222 230058 588458 230294
rect 588542 230058 588778 230294
rect 588222 194378 588458 194614
rect 588542 194378 588778 194614
rect 588222 194058 588458 194294
rect 588542 194058 588778 194294
rect 588222 158378 588458 158614
rect 588542 158378 588778 158614
rect 588222 158058 588458 158294
rect 588542 158058 588778 158294
rect 588222 122378 588458 122614
rect 588542 122378 588778 122614
rect 588222 122058 588458 122294
rect 588542 122058 588778 122294
rect 588222 86378 588458 86614
rect 588542 86378 588778 86614
rect 588222 86058 588458 86294
rect 588542 86058 588778 86294
rect 588222 50378 588458 50614
rect 588542 50378 588778 50614
rect 588222 50058 588458 50294
rect 588542 50058 588778 50294
rect 588222 14378 588458 14614
rect 588542 14378 588778 14614
rect 588222 14058 588458 14294
rect 588542 14058 588778 14294
rect 588222 -3462 588458 -3226
rect 588542 -3462 588778 -3226
rect 588222 -3782 588458 -3546
rect 588542 -3782 588778 -3546
rect 589182 666098 589418 666334
rect 589502 666098 589738 666334
rect 589182 665778 589418 666014
rect 589502 665778 589738 666014
rect 589182 630098 589418 630334
rect 589502 630098 589738 630334
rect 589182 629778 589418 630014
rect 589502 629778 589738 630014
rect 589182 594098 589418 594334
rect 589502 594098 589738 594334
rect 589182 593778 589418 594014
rect 589502 593778 589738 594014
rect 589182 558098 589418 558334
rect 589502 558098 589738 558334
rect 589182 557778 589418 558014
rect 589502 557778 589738 558014
rect 589182 522098 589418 522334
rect 589502 522098 589738 522334
rect 589182 521778 589418 522014
rect 589502 521778 589738 522014
rect 589182 486098 589418 486334
rect 589502 486098 589738 486334
rect 589182 485778 589418 486014
rect 589502 485778 589738 486014
rect 589182 450098 589418 450334
rect 589502 450098 589738 450334
rect 589182 449778 589418 450014
rect 589502 449778 589738 450014
rect 589182 414098 589418 414334
rect 589502 414098 589738 414334
rect 589182 413778 589418 414014
rect 589502 413778 589738 414014
rect 589182 378098 589418 378334
rect 589502 378098 589738 378334
rect 589182 377778 589418 378014
rect 589502 377778 589738 378014
rect 589182 342098 589418 342334
rect 589502 342098 589738 342334
rect 589182 341778 589418 342014
rect 589502 341778 589738 342014
rect 589182 306098 589418 306334
rect 589502 306098 589738 306334
rect 589182 305778 589418 306014
rect 589502 305778 589738 306014
rect 589182 270098 589418 270334
rect 589502 270098 589738 270334
rect 589182 269778 589418 270014
rect 589502 269778 589738 270014
rect 589182 234098 589418 234334
rect 589502 234098 589738 234334
rect 589182 233778 589418 234014
rect 589502 233778 589738 234014
rect 589182 198098 589418 198334
rect 589502 198098 589738 198334
rect 589182 197778 589418 198014
rect 589502 197778 589738 198014
rect 589182 162098 589418 162334
rect 589502 162098 589738 162334
rect 589182 161778 589418 162014
rect 589502 161778 589738 162014
rect 589182 126098 589418 126334
rect 589502 126098 589738 126334
rect 589182 125778 589418 126014
rect 589502 125778 589738 126014
rect 589182 90098 589418 90334
rect 589502 90098 589738 90334
rect 589182 89778 589418 90014
rect 589502 89778 589738 90014
rect 589182 54098 589418 54334
rect 589502 54098 589738 54334
rect 589182 53778 589418 54014
rect 589502 53778 589738 54014
rect 589182 18098 589418 18334
rect 589502 18098 589738 18334
rect 589182 17778 589418 18014
rect 589502 17778 589738 18014
rect 589182 -4422 589418 -4186
rect 589502 -4422 589738 -4186
rect 589182 -4742 589418 -4506
rect 589502 -4742 589738 -4506
rect 590142 669818 590378 670054
rect 590462 669818 590698 670054
rect 590142 669498 590378 669734
rect 590462 669498 590698 669734
rect 590142 633818 590378 634054
rect 590462 633818 590698 634054
rect 590142 633498 590378 633734
rect 590462 633498 590698 633734
rect 590142 597818 590378 598054
rect 590462 597818 590698 598054
rect 590142 597498 590378 597734
rect 590462 597498 590698 597734
rect 590142 561818 590378 562054
rect 590462 561818 590698 562054
rect 590142 561498 590378 561734
rect 590462 561498 590698 561734
rect 590142 525818 590378 526054
rect 590462 525818 590698 526054
rect 590142 525498 590378 525734
rect 590462 525498 590698 525734
rect 590142 489818 590378 490054
rect 590462 489818 590698 490054
rect 590142 489498 590378 489734
rect 590462 489498 590698 489734
rect 590142 453818 590378 454054
rect 590462 453818 590698 454054
rect 590142 453498 590378 453734
rect 590462 453498 590698 453734
rect 590142 417818 590378 418054
rect 590462 417818 590698 418054
rect 590142 417498 590378 417734
rect 590462 417498 590698 417734
rect 590142 381818 590378 382054
rect 590462 381818 590698 382054
rect 590142 381498 590378 381734
rect 590462 381498 590698 381734
rect 590142 345818 590378 346054
rect 590462 345818 590698 346054
rect 590142 345498 590378 345734
rect 590462 345498 590698 345734
rect 590142 309818 590378 310054
rect 590462 309818 590698 310054
rect 590142 309498 590378 309734
rect 590462 309498 590698 309734
rect 590142 273818 590378 274054
rect 590462 273818 590698 274054
rect 590142 273498 590378 273734
rect 590462 273498 590698 273734
rect 590142 237818 590378 238054
rect 590462 237818 590698 238054
rect 590142 237498 590378 237734
rect 590462 237498 590698 237734
rect 590142 201818 590378 202054
rect 590462 201818 590698 202054
rect 590142 201498 590378 201734
rect 590462 201498 590698 201734
rect 590142 165818 590378 166054
rect 590462 165818 590698 166054
rect 590142 165498 590378 165734
rect 590462 165498 590698 165734
rect 590142 129818 590378 130054
rect 590462 129818 590698 130054
rect 590142 129498 590378 129734
rect 590462 129498 590698 129734
rect 590142 93818 590378 94054
rect 590462 93818 590698 94054
rect 590142 93498 590378 93734
rect 590462 93498 590698 93734
rect 590142 57818 590378 58054
rect 590462 57818 590698 58054
rect 590142 57498 590378 57734
rect 590462 57498 590698 57734
rect 590142 21818 590378 22054
rect 590462 21818 590698 22054
rect 590142 21498 590378 21734
rect 590462 21498 590698 21734
rect 590142 -5382 590378 -5146
rect 590462 -5382 590698 -5146
rect 590142 -5702 590378 -5466
rect 590462 -5702 590698 -5466
rect 591102 673538 591338 673774
rect 591422 673538 591658 673774
rect 591102 673218 591338 673454
rect 591422 673218 591658 673454
rect 591102 637538 591338 637774
rect 591422 637538 591658 637774
rect 591102 637218 591338 637454
rect 591422 637218 591658 637454
rect 591102 601538 591338 601774
rect 591422 601538 591658 601774
rect 591102 601218 591338 601454
rect 591422 601218 591658 601454
rect 591102 565538 591338 565774
rect 591422 565538 591658 565774
rect 591102 565218 591338 565454
rect 591422 565218 591658 565454
rect 591102 529538 591338 529774
rect 591422 529538 591658 529774
rect 591102 529218 591338 529454
rect 591422 529218 591658 529454
rect 591102 493538 591338 493774
rect 591422 493538 591658 493774
rect 591102 493218 591338 493454
rect 591422 493218 591658 493454
rect 591102 457538 591338 457774
rect 591422 457538 591658 457774
rect 591102 457218 591338 457454
rect 591422 457218 591658 457454
rect 591102 421538 591338 421774
rect 591422 421538 591658 421774
rect 591102 421218 591338 421454
rect 591422 421218 591658 421454
rect 591102 385538 591338 385774
rect 591422 385538 591658 385774
rect 591102 385218 591338 385454
rect 591422 385218 591658 385454
rect 591102 349538 591338 349774
rect 591422 349538 591658 349774
rect 591102 349218 591338 349454
rect 591422 349218 591658 349454
rect 591102 313538 591338 313774
rect 591422 313538 591658 313774
rect 591102 313218 591338 313454
rect 591422 313218 591658 313454
rect 591102 277538 591338 277774
rect 591422 277538 591658 277774
rect 591102 277218 591338 277454
rect 591422 277218 591658 277454
rect 591102 241538 591338 241774
rect 591422 241538 591658 241774
rect 591102 241218 591338 241454
rect 591422 241218 591658 241454
rect 591102 205538 591338 205774
rect 591422 205538 591658 205774
rect 591102 205218 591338 205454
rect 591422 205218 591658 205454
rect 591102 169538 591338 169774
rect 591422 169538 591658 169774
rect 591102 169218 591338 169454
rect 591422 169218 591658 169454
rect 591102 133538 591338 133774
rect 591422 133538 591658 133774
rect 591102 133218 591338 133454
rect 591422 133218 591658 133454
rect 591102 97538 591338 97774
rect 591422 97538 591658 97774
rect 591102 97218 591338 97454
rect 591422 97218 591658 97454
rect 591102 61538 591338 61774
rect 591422 61538 591658 61774
rect 591102 61218 591338 61454
rect 591422 61218 591658 61454
rect 591102 25538 591338 25774
rect 591422 25538 591658 25774
rect 591102 25218 591338 25454
rect 591422 25218 591658 25454
rect 591102 -6342 591338 -6106
rect 591422 -6342 591658 -6106
rect 591102 -6662 591338 -6426
rect 591422 -6662 591658 -6426
rect 592062 677258 592298 677494
rect 592382 677258 592618 677494
rect 592062 676938 592298 677174
rect 592382 676938 592618 677174
rect 592062 641258 592298 641494
rect 592382 641258 592618 641494
rect 592062 640938 592298 641174
rect 592382 640938 592618 641174
rect 592062 605258 592298 605494
rect 592382 605258 592618 605494
rect 592062 604938 592298 605174
rect 592382 604938 592618 605174
rect 592062 569258 592298 569494
rect 592382 569258 592618 569494
rect 592062 568938 592298 569174
rect 592382 568938 592618 569174
rect 592062 533258 592298 533494
rect 592382 533258 592618 533494
rect 592062 532938 592298 533174
rect 592382 532938 592618 533174
rect 592062 497258 592298 497494
rect 592382 497258 592618 497494
rect 592062 496938 592298 497174
rect 592382 496938 592618 497174
rect 592062 461258 592298 461494
rect 592382 461258 592618 461494
rect 592062 460938 592298 461174
rect 592382 460938 592618 461174
rect 592062 425258 592298 425494
rect 592382 425258 592618 425494
rect 592062 424938 592298 425174
rect 592382 424938 592618 425174
rect 592062 389258 592298 389494
rect 592382 389258 592618 389494
rect 592062 388938 592298 389174
rect 592382 388938 592618 389174
rect 592062 353258 592298 353494
rect 592382 353258 592618 353494
rect 592062 352938 592298 353174
rect 592382 352938 592618 353174
rect 592062 317258 592298 317494
rect 592382 317258 592618 317494
rect 592062 316938 592298 317174
rect 592382 316938 592618 317174
rect 592062 281258 592298 281494
rect 592382 281258 592618 281494
rect 592062 280938 592298 281174
rect 592382 280938 592618 281174
rect 592062 245258 592298 245494
rect 592382 245258 592618 245494
rect 592062 244938 592298 245174
rect 592382 244938 592618 245174
rect 592062 209258 592298 209494
rect 592382 209258 592618 209494
rect 592062 208938 592298 209174
rect 592382 208938 592618 209174
rect 592062 173258 592298 173494
rect 592382 173258 592618 173494
rect 592062 172938 592298 173174
rect 592382 172938 592618 173174
rect 592062 137258 592298 137494
rect 592382 137258 592618 137494
rect 592062 136938 592298 137174
rect 592382 136938 592618 137174
rect 592062 101258 592298 101494
rect 592382 101258 592618 101494
rect 592062 100938 592298 101174
rect 592382 100938 592618 101174
rect 592062 65258 592298 65494
rect 592382 65258 592618 65494
rect 592062 64938 592298 65174
rect 592382 64938 592618 65174
rect 592062 29258 592298 29494
rect 592382 29258 592618 29494
rect 592062 28938 592298 29174
rect 592382 28938 592618 29174
rect 592062 -7302 592298 -7066
rect 592382 -7302 592618 -7066
rect 592062 -7622 592298 -7386
rect 592382 -7622 592618 -7386
<< metal5 >>
rect -8726 711558 592650 711590
rect -8726 711322 -8694 711558
rect -8458 711322 -8374 711558
rect -8138 711322 27866 711558
rect 28102 711322 28186 711558
rect 28422 711322 63866 711558
rect 64102 711322 64186 711558
rect 64422 711322 99866 711558
rect 100102 711322 100186 711558
rect 100422 711322 135866 711558
rect 136102 711322 136186 711558
rect 136422 711322 171866 711558
rect 172102 711322 172186 711558
rect 172422 711322 207866 711558
rect 208102 711322 208186 711558
rect 208422 711322 243866 711558
rect 244102 711322 244186 711558
rect 244422 711322 279866 711558
rect 280102 711322 280186 711558
rect 280422 711322 315866 711558
rect 316102 711322 316186 711558
rect 316422 711322 351866 711558
rect 352102 711322 352186 711558
rect 352422 711322 387866 711558
rect 388102 711322 388186 711558
rect 388422 711322 423866 711558
rect 424102 711322 424186 711558
rect 424422 711322 459866 711558
rect 460102 711322 460186 711558
rect 460422 711322 495866 711558
rect 496102 711322 496186 711558
rect 496422 711322 531866 711558
rect 532102 711322 532186 711558
rect 532422 711322 567866 711558
rect 568102 711322 568186 711558
rect 568422 711322 592062 711558
rect 592298 711322 592382 711558
rect 592618 711322 592650 711558
rect -8726 711238 592650 711322
rect -8726 711002 -8694 711238
rect -8458 711002 -8374 711238
rect -8138 711002 27866 711238
rect 28102 711002 28186 711238
rect 28422 711002 63866 711238
rect 64102 711002 64186 711238
rect 64422 711002 99866 711238
rect 100102 711002 100186 711238
rect 100422 711002 135866 711238
rect 136102 711002 136186 711238
rect 136422 711002 171866 711238
rect 172102 711002 172186 711238
rect 172422 711002 207866 711238
rect 208102 711002 208186 711238
rect 208422 711002 243866 711238
rect 244102 711002 244186 711238
rect 244422 711002 279866 711238
rect 280102 711002 280186 711238
rect 280422 711002 315866 711238
rect 316102 711002 316186 711238
rect 316422 711002 351866 711238
rect 352102 711002 352186 711238
rect 352422 711002 387866 711238
rect 388102 711002 388186 711238
rect 388422 711002 423866 711238
rect 424102 711002 424186 711238
rect 424422 711002 459866 711238
rect 460102 711002 460186 711238
rect 460422 711002 495866 711238
rect 496102 711002 496186 711238
rect 496422 711002 531866 711238
rect 532102 711002 532186 711238
rect 532422 711002 567866 711238
rect 568102 711002 568186 711238
rect 568422 711002 592062 711238
rect 592298 711002 592382 711238
rect 592618 711002 592650 711238
rect -8726 710970 592650 711002
rect -7766 710598 591690 710630
rect -7766 710362 -7734 710598
rect -7498 710362 -7414 710598
rect -7178 710362 24146 710598
rect 24382 710362 24466 710598
rect 24702 710362 60146 710598
rect 60382 710362 60466 710598
rect 60702 710362 96146 710598
rect 96382 710362 96466 710598
rect 96702 710362 132146 710598
rect 132382 710362 132466 710598
rect 132702 710362 168146 710598
rect 168382 710362 168466 710598
rect 168702 710362 204146 710598
rect 204382 710362 204466 710598
rect 204702 710362 240146 710598
rect 240382 710362 240466 710598
rect 240702 710362 276146 710598
rect 276382 710362 276466 710598
rect 276702 710362 312146 710598
rect 312382 710362 312466 710598
rect 312702 710362 348146 710598
rect 348382 710362 348466 710598
rect 348702 710362 384146 710598
rect 384382 710362 384466 710598
rect 384702 710362 420146 710598
rect 420382 710362 420466 710598
rect 420702 710362 456146 710598
rect 456382 710362 456466 710598
rect 456702 710362 492146 710598
rect 492382 710362 492466 710598
rect 492702 710362 528146 710598
rect 528382 710362 528466 710598
rect 528702 710362 564146 710598
rect 564382 710362 564466 710598
rect 564702 710362 591102 710598
rect 591338 710362 591422 710598
rect 591658 710362 591690 710598
rect -7766 710278 591690 710362
rect -7766 710042 -7734 710278
rect -7498 710042 -7414 710278
rect -7178 710042 24146 710278
rect 24382 710042 24466 710278
rect 24702 710042 60146 710278
rect 60382 710042 60466 710278
rect 60702 710042 96146 710278
rect 96382 710042 96466 710278
rect 96702 710042 132146 710278
rect 132382 710042 132466 710278
rect 132702 710042 168146 710278
rect 168382 710042 168466 710278
rect 168702 710042 204146 710278
rect 204382 710042 204466 710278
rect 204702 710042 240146 710278
rect 240382 710042 240466 710278
rect 240702 710042 276146 710278
rect 276382 710042 276466 710278
rect 276702 710042 312146 710278
rect 312382 710042 312466 710278
rect 312702 710042 348146 710278
rect 348382 710042 348466 710278
rect 348702 710042 384146 710278
rect 384382 710042 384466 710278
rect 384702 710042 420146 710278
rect 420382 710042 420466 710278
rect 420702 710042 456146 710278
rect 456382 710042 456466 710278
rect 456702 710042 492146 710278
rect 492382 710042 492466 710278
rect 492702 710042 528146 710278
rect 528382 710042 528466 710278
rect 528702 710042 564146 710278
rect 564382 710042 564466 710278
rect 564702 710042 591102 710278
rect 591338 710042 591422 710278
rect 591658 710042 591690 710278
rect -7766 710010 591690 710042
rect -6806 709638 590730 709670
rect -6806 709402 -6774 709638
rect -6538 709402 -6454 709638
rect -6218 709402 20426 709638
rect 20662 709402 20746 709638
rect 20982 709402 56426 709638
rect 56662 709402 56746 709638
rect 56982 709402 92426 709638
rect 92662 709402 92746 709638
rect 92982 709402 128426 709638
rect 128662 709402 128746 709638
rect 128982 709402 164426 709638
rect 164662 709402 164746 709638
rect 164982 709402 200426 709638
rect 200662 709402 200746 709638
rect 200982 709402 236426 709638
rect 236662 709402 236746 709638
rect 236982 709402 272426 709638
rect 272662 709402 272746 709638
rect 272982 709402 308426 709638
rect 308662 709402 308746 709638
rect 308982 709402 344426 709638
rect 344662 709402 344746 709638
rect 344982 709402 380426 709638
rect 380662 709402 380746 709638
rect 380982 709402 416426 709638
rect 416662 709402 416746 709638
rect 416982 709402 452426 709638
rect 452662 709402 452746 709638
rect 452982 709402 488426 709638
rect 488662 709402 488746 709638
rect 488982 709402 524426 709638
rect 524662 709402 524746 709638
rect 524982 709402 560426 709638
rect 560662 709402 560746 709638
rect 560982 709402 590142 709638
rect 590378 709402 590462 709638
rect 590698 709402 590730 709638
rect -6806 709318 590730 709402
rect -6806 709082 -6774 709318
rect -6538 709082 -6454 709318
rect -6218 709082 20426 709318
rect 20662 709082 20746 709318
rect 20982 709082 56426 709318
rect 56662 709082 56746 709318
rect 56982 709082 92426 709318
rect 92662 709082 92746 709318
rect 92982 709082 128426 709318
rect 128662 709082 128746 709318
rect 128982 709082 164426 709318
rect 164662 709082 164746 709318
rect 164982 709082 200426 709318
rect 200662 709082 200746 709318
rect 200982 709082 236426 709318
rect 236662 709082 236746 709318
rect 236982 709082 272426 709318
rect 272662 709082 272746 709318
rect 272982 709082 308426 709318
rect 308662 709082 308746 709318
rect 308982 709082 344426 709318
rect 344662 709082 344746 709318
rect 344982 709082 380426 709318
rect 380662 709082 380746 709318
rect 380982 709082 416426 709318
rect 416662 709082 416746 709318
rect 416982 709082 452426 709318
rect 452662 709082 452746 709318
rect 452982 709082 488426 709318
rect 488662 709082 488746 709318
rect 488982 709082 524426 709318
rect 524662 709082 524746 709318
rect 524982 709082 560426 709318
rect 560662 709082 560746 709318
rect 560982 709082 590142 709318
rect 590378 709082 590462 709318
rect 590698 709082 590730 709318
rect -6806 709050 590730 709082
rect -5846 708678 589770 708710
rect -5846 708442 -5814 708678
rect -5578 708442 -5494 708678
rect -5258 708442 16706 708678
rect 16942 708442 17026 708678
rect 17262 708442 52706 708678
rect 52942 708442 53026 708678
rect 53262 708442 88706 708678
rect 88942 708442 89026 708678
rect 89262 708442 124706 708678
rect 124942 708442 125026 708678
rect 125262 708442 160706 708678
rect 160942 708442 161026 708678
rect 161262 708442 196706 708678
rect 196942 708442 197026 708678
rect 197262 708442 232706 708678
rect 232942 708442 233026 708678
rect 233262 708442 268706 708678
rect 268942 708442 269026 708678
rect 269262 708442 304706 708678
rect 304942 708442 305026 708678
rect 305262 708442 340706 708678
rect 340942 708442 341026 708678
rect 341262 708442 376706 708678
rect 376942 708442 377026 708678
rect 377262 708442 412706 708678
rect 412942 708442 413026 708678
rect 413262 708442 448706 708678
rect 448942 708442 449026 708678
rect 449262 708442 484706 708678
rect 484942 708442 485026 708678
rect 485262 708442 520706 708678
rect 520942 708442 521026 708678
rect 521262 708442 556706 708678
rect 556942 708442 557026 708678
rect 557262 708442 589182 708678
rect 589418 708442 589502 708678
rect 589738 708442 589770 708678
rect -5846 708358 589770 708442
rect -5846 708122 -5814 708358
rect -5578 708122 -5494 708358
rect -5258 708122 16706 708358
rect 16942 708122 17026 708358
rect 17262 708122 52706 708358
rect 52942 708122 53026 708358
rect 53262 708122 88706 708358
rect 88942 708122 89026 708358
rect 89262 708122 124706 708358
rect 124942 708122 125026 708358
rect 125262 708122 160706 708358
rect 160942 708122 161026 708358
rect 161262 708122 196706 708358
rect 196942 708122 197026 708358
rect 197262 708122 232706 708358
rect 232942 708122 233026 708358
rect 233262 708122 268706 708358
rect 268942 708122 269026 708358
rect 269262 708122 304706 708358
rect 304942 708122 305026 708358
rect 305262 708122 340706 708358
rect 340942 708122 341026 708358
rect 341262 708122 376706 708358
rect 376942 708122 377026 708358
rect 377262 708122 412706 708358
rect 412942 708122 413026 708358
rect 413262 708122 448706 708358
rect 448942 708122 449026 708358
rect 449262 708122 484706 708358
rect 484942 708122 485026 708358
rect 485262 708122 520706 708358
rect 520942 708122 521026 708358
rect 521262 708122 556706 708358
rect 556942 708122 557026 708358
rect 557262 708122 589182 708358
rect 589418 708122 589502 708358
rect 589738 708122 589770 708358
rect -5846 708090 589770 708122
rect -4886 707718 588810 707750
rect -4886 707482 -4854 707718
rect -4618 707482 -4534 707718
rect -4298 707482 12986 707718
rect 13222 707482 13306 707718
rect 13542 707482 48986 707718
rect 49222 707482 49306 707718
rect 49542 707482 84986 707718
rect 85222 707482 85306 707718
rect 85542 707482 120986 707718
rect 121222 707482 121306 707718
rect 121542 707482 156986 707718
rect 157222 707482 157306 707718
rect 157542 707482 192986 707718
rect 193222 707482 193306 707718
rect 193542 707482 228986 707718
rect 229222 707482 229306 707718
rect 229542 707482 264986 707718
rect 265222 707482 265306 707718
rect 265542 707482 300986 707718
rect 301222 707482 301306 707718
rect 301542 707482 336986 707718
rect 337222 707482 337306 707718
rect 337542 707482 372986 707718
rect 373222 707482 373306 707718
rect 373542 707482 408986 707718
rect 409222 707482 409306 707718
rect 409542 707482 444986 707718
rect 445222 707482 445306 707718
rect 445542 707482 480986 707718
rect 481222 707482 481306 707718
rect 481542 707482 516986 707718
rect 517222 707482 517306 707718
rect 517542 707482 552986 707718
rect 553222 707482 553306 707718
rect 553542 707482 588222 707718
rect 588458 707482 588542 707718
rect 588778 707482 588810 707718
rect -4886 707398 588810 707482
rect -4886 707162 -4854 707398
rect -4618 707162 -4534 707398
rect -4298 707162 12986 707398
rect 13222 707162 13306 707398
rect 13542 707162 48986 707398
rect 49222 707162 49306 707398
rect 49542 707162 84986 707398
rect 85222 707162 85306 707398
rect 85542 707162 120986 707398
rect 121222 707162 121306 707398
rect 121542 707162 156986 707398
rect 157222 707162 157306 707398
rect 157542 707162 192986 707398
rect 193222 707162 193306 707398
rect 193542 707162 228986 707398
rect 229222 707162 229306 707398
rect 229542 707162 264986 707398
rect 265222 707162 265306 707398
rect 265542 707162 300986 707398
rect 301222 707162 301306 707398
rect 301542 707162 336986 707398
rect 337222 707162 337306 707398
rect 337542 707162 372986 707398
rect 373222 707162 373306 707398
rect 373542 707162 408986 707398
rect 409222 707162 409306 707398
rect 409542 707162 444986 707398
rect 445222 707162 445306 707398
rect 445542 707162 480986 707398
rect 481222 707162 481306 707398
rect 481542 707162 516986 707398
rect 517222 707162 517306 707398
rect 517542 707162 552986 707398
rect 553222 707162 553306 707398
rect 553542 707162 588222 707398
rect 588458 707162 588542 707398
rect 588778 707162 588810 707398
rect -4886 707130 588810 707162
rect -3926 706758 587850 706790
rect -3926 706522 -3894 706758
rect -3658 706522 -3574 706758
rect -3338 706522 9266 706758
rect 9502 706522 9586 706758
rect 9822 706522 45266 706758
rect 45502 706522 45586 706758
rect 45822 706522 81266 706758
rect 81502 706522 81586 706758
rect 81822 706522 117266 706758
rect 117502 706522 117586 706758
rect 117822 706522 153266 706758
rect 153502 706522 153586 706758
rect 153822 706522 189266 706758
rect 189502 706522 189586 706758
rect 189822 706522 225266 706758
rect 225502 706522 225586 706758
rect 225822 706522 261266 706758
rect 261502 706522 261586 706758
rect 261822 706522 297266 706758
rect 297502 706522 297586 706758
rect 297822 706522 333266 706758
rect 333502 706522 333586 706758
rect 333822 706522 369266 706758
rect 369502 706522 369586 706758
rect 369822 706522 405266 706758
rect 405502 706522 405586 706758
rect 405822 706522 441266 706758
rect 441502 706522 441586 706758
rect 441822 706522 477266 706758
rect 477502 706522 477586 706758
rect 477822 706522 513266 706758
rect 513502 706522 513586 706758
rect 513822 706522 549266 706758
rect 549502 706522 549586 706758
rect 549822 706522 587262 706758
rect 587498 706522 587582 706758
rect 587818 706522 587850 706758
rect -3926 706438 587850 706522
rect -3926 706202 -3894 706438
rect -3658 706202 -3574 706438
rect -3338 706202 9266 706438
rect 9502 706202 9586 706438
rect 9822 706202 45266 706438
rect 45502 706202 45586 706438
rect 45822 706202 81266 706438
rect 81502 706202 81586 706438
rect 81822 706202 117266 706438
rect 117502 706202 117586 706438
rect 117822 706202 153266 706438
rect 153502 706202 153586 706438
rect 153822 706202 189266 706438
rect 189502 706202 189586 706438
rect 189822 706202 225266 706438
rect 225502 706202 225586 706438
rect 225822 706202 261266 706438
rect 261502 706202 261586 706438
rect 261822 706202 297266 706438
rect 297502 706202 297586 706438
rect 297822 706202 333266 706438
rect 333502 706202 333586 706438
rect 333822 706202 369266 706438
rect 369502 706202 369586 706438
rect 369822 706202 405266 706438
rect 405502 706202 405586 706438
rect 405822 706202 441266 706438
rect 441502 706202 441586 706438
rect 441822 706202 477266 706438
rect 477502 706202 477586 706438
rect 477822 706202 513266 706438
rect 513502 706202 513586 706438
rect 513822 706202 549266 706438
rect 549502 706202 549586 706438
rect 549822 706202 587262 706438
rect 587498 706202 587582 706438
rect 587818 706202 587850 706438
rect -3926 706170 587850 706202
rect -2966 705798 586890 705830
rect -2966 705562 -2934 705798
rect -2698 705562 -2614 705798
rect -2378 705562 5546 705798
rect 5782 705562 5866 705798
rect 6102 705562 41546 705798
rect 41782 705562 41866 705798
rect 42102 705562 77546 705798
rect 77782 705562 77866 705798
rect 78102 705562 113546 705798
rect 113782 705562 113866 705798
rect 114102 705562 149546 705798
rect 149782 705562 149866 705798
rect 150102 705562 185546 705798
rect 185782 705562 185866 705798
rect 186102 705562 221546 705798
rect 221782 705562 221866 705798
rect 222102 705562 257546 705798
rect 257782 705562 257866 705798
rect 258102 705562 293546 705798
rect 293782 705562 293866 705798
rect 294102 705562 329546 705798
rect 329782 705562 329866 705798
rect 330102 705562 365546 705798
rect 365782 705562 365866 705798
rect 366102 705562 401546 705798
rect 401782 705562 401866 705798
rect 402102 705562 437546 705798
rect 437782 705562 437866 705798
rect 438102 705562 473546 705798
rect 473782 705562 473866 705798
rect 474102 705562 509546 705798
rect 509782 705562 509866 705798
rect 510102 705562 545546 705798
rect 545782 705562 545866 705798
rect 546102 705562 581546 705798
rect 581782 705562 581866 705798
rect 582102 705562 586302 705798
rect 586538 705562 586622 705798
rect 586858 705562 586890 705798
rect -2966 705478 586890 705562
rect -2966 705242 -2934 705478
rect -2698 705242 -2614 705478
rect -2378 705242 5546 705478
rect 5782 705242 5866 705478
rect 6102 705242 41546 705478
rect 41782 705242 41866 705478
rect 42102 705242 77546 705478
rect 77782 705242 77866 705478
rect 78102 705242 113546 705478
rect 113782 705242 113866 705478
rect 114102 705242 149546 705478
rect 149782 705242 149866 705478
rect 150102 705242 185546 705478
rect 185782 705242 185866 705478
rect 186102 705242 221546 705478
rect 221782 705242 221866 705478
rect 222102 705242 257546 705478
rect 257782 705242 257866 705478
rect 258102 705242 293546 705478
rect 293782 705242 293866 705478
rect 294102 705242 329546 705478
rect 329782 705242 329866 705478
rect 330102 705242 365546 705478
rect 365782 705242 365866 705478
rect 366102 705242 401546 705478
rect 401782 705242 401866 705478
rect 402102 705242 437546 705478
rect 437782 705242 437866 705478
rect 438102 705242 473546 705478
rect 473782 705242 473866 705478
rect 474102 705242 509546 705478
rect 509782 705242 509866 705478
rect 510102 705242 545546 705478
rect 545782 705242 545866 705478
rect 546102 705242 581546 705478
rect 581782 705242 581866 705478
rect 582102 705242 586302 705478
rect 586538 705242 586622 705478
rect 586858 705242 586890 705478
rect -2966 705210 586890 705242
rect -2006 704838 585930 704870
rect -2006 704602 -1974 704838
rect -1738 704602 -1654 704838
rect -1418 704602 1826 704838
rect 2062 704602 2146 704838
rect 2382 704602 37826 704838
rect 38062 704602 38146 704838
rect 38382 704602 73826 704838
rect 74062 704602 74146 704838
rect 74382 704602 109826 704838
rect 110062 704602 110146 704838
rect 110382 704602 145826 704838
rect 146062 704602 146146 704838
rect 146382 704602 181826 704838
rect 182062 704602 182146 704838
rect 182382 704602 217826 704838
rect 218062 704602 218146 704838
rect 218382 704602 253826 704838
rect 254062 704602 254146 704838
rect 254382 704602 289826 704838
rect 290062 704602 290146 704838
rect 290382 704602 325826 704838
rect 326062 704602 326146 704838
rect 326382 704602 361826 704838
rect 362062 704602 362146 704838
rect 362382 704602 397826 704838
rect 398062 704602 398146 704838
rect 398382 704602 433826 704838
rect 434062 704602 434146 704838
rect 434382 704602 469826 704838
rect 470062 704602 470146 704838
rect 470382 704602 505826 704838
rect 506062 704602 506146 704838
rect 506382 704602 541826 704838
rect 542062 704602 542146 704838
rect 542382 704602 577826 704838
rect 578062 704602 578146 704838
rect 578382 704602 585342 704838
rect 585578 704602 585662 704838
rect 585898 704602 585930 704838
rect -2006 704518 585930 704602
rect -2006 704282 -1974 704518
rect -1738 704282 -1654 704518
rect -1418 704282 1826 704518
rect 2062 704282 2146 704518
rect 2382 704282 37826 704518
rect 38062 704282 38146 704518
rect 38382 704282 73826 704518
rect 74062 704282 74146 704518
rect 74382 704282 109826 704518
rect 110062 704282 110146 704518
rect 110382 704282 145826 704518
rect 146062 704282 146146 704518
rect 146382 704282 181826 704518
rect 182062 704282 182146 704518
rect 182382 704282 217826 704518
rect 218062 704282 218146 704518
rect 218382 704282 253826 704518
rect 254062 704282 254146 704518
rect 254382 704282 289826 704518
rect 290062 704282 290146 704518
rect 290382 704282 325826 704518
rect 326062 704282 326146 704518
rect 326382 704282 361826 704518
rect 362062 704282 362146 704518
rect 362382 704282 397826 704518
rect 398062 704282 398146 704518
rect 398382 704282 433826 704518
rect 434062 704282 434146 704518
rect 434382 704282 469826 704518
rect 470062 704282 470146 704518
rect 470382 704282 505826 704518
rect 506062 704282 506146 704518
rect 506382 704282 541826 704518
rect 542062 704282 542146 704518
rect 542382 704282 577826 704518
rect 578062 704282 578146 704518
rect 578382 704282 585342 704518
rect 585578 704282 585662 704518
rect 585898 704282 585930 704518
rect -2006 704250 585930 704282
rect -8726 698614 592650 698646
rect -8726 698378 -4854 698614
rect -4618 698378 -4534 698614
rect -4298 698378 12986 698614
rect 13222 698378 13306 698614
rect 13542 698378 48986 698614
rect 49222 698378 49306 698614
rect 49542 698378 84986 698614
rect 85222 698378 85306 698614
rect 85542 698378 120986 698614
rect 121222 698378 121306 698614
rect 121542 698378 156986 698614
rect 157222 698378 157306 698614
rect 157542 698378 192986 698614
rect 193222 698378 193306 698614
rect 193542 698378 228986 698614
rect 229222 698378 229306 698614
rect 229542 698378 264986 698614
rect 265222 698378 265306 698614
rect 265542 698378 300986 698614
rect 301222 698378 301306 698614
rect 301542 698378 336986 698614
rect 337222 698378 337306 698614
rect 337542 698378 372986 698614
rect 373222 698378 373306 698614
rect 373542 698378 408986 698614
rect 409222 698378 409306 698614
rect 409542 698378 444986 698614
rect 445222 698378 445306 698614
rect 445542 698378 480986 698614
rect 481222 698378 481306 698614
rect 481542 698378 516986 698614
rect 517222 698378 517306 698614
rect 517542 698378 552986 698614
rect 553222 698378 553306 698614
rect 553542 698378 588222 698614
rect 588458 698378 588542 698614
rect 588778 698378 592650 698614
rect -8726 698294 592650 698378
rect -8726 698058 -4854 698294
rect -4618 698058 -4534 698294
rect -4298 698058 12986 698294
rect 13222 698058 13306 698294
rect 13542 698058 48986 698294
rect 49222 698058 49306 698294
rect 49542 698058 84986 698294
rect 85222 698058 85306 698294
rect 85542 698058 120986 698294
rect 121222 698058 121306 698294
rect 121542 698058 156986 698294
rect 157222 698058 157306 698294
rect 157542 698058 192986 698294
rect 193222 698058 193306 698294
rect 193542 698058 228986 698294
rect 229222 698058 229306 698294
rect 229542 698058 264986 698294
rect 265222 698058 265306 698294
rect 265542 698058 300986 698294
rect 301222 698058 301306 698294
rect 301542 698058 336986 698294
rect 337222 698058 337306 698294
rect 337542 698058 372986 698294
rect 373222 698058 373306 698294
rect 373542 698058 408986 698294
rect 409222 698058 409306 698294
rect 409542 698058 444986 698294
rect 445222 698058 445306 698294
rect 445542 698058 480986 698294
rect 481222 698058 481306 698294
rect 481542 698058 516986 698294
rect 517222 698058 517306 698294
rect 517542 698058 552986 698294
rect 553222 698058 553306 698294
rect 553542 698058 588222 698294
rect 588458 698058 588542 698294
rect 588778 698058 592650 698294
rect -8726 698026 592650 698058
rect -8726 694894 592650 694926
rect -8726 694658 -3894 694894
rect -3658 694658 -3574 694894
rect -3338 694658 9266 694894
rect 9502 694658 9586 694894
rect 9822 694658 45266 694894
rect 45502 694658 45586 694894
rect 45822 694658 81266 694894
rect 81502 694658 81586 694894
rect 81822 694658 117266 694894
rect 117502 694658 117586 694894
rect 117822 694658 153266 694894
rect 153502 694658 153586 694894
rect 153822 694658 189266 694894
rect 189502 694658 189586 694894
rect 189822 694658 225266 694894
rect 225502 694658 225586 694894
rect 225822 694658 261266 694894
rect 261502 694658 261586 694894
rect 261822 694658 297266 694894
rect 297502 694658 297586 694894
rect 297822 694658 333266 694894
rect 333502 694658 333586 694894
rect 333822 694658 369266 694894
rect 369502 694658 369586 694894
rect 369822 694658 405266 694894
rect 405502 694658 405586 694894
rect 405822 694658 441266 694894
rect 441502 694658 441586 694894
rect 441822 694658 477266 694894
rect 477502 694658 477586 694894
rect 477822 694658 513266 694894
rect 513502 694658 513586 694894
rect 513822 694658 549266 694894
rect 549502 694658 549586 694894
rect 549822 694658 587262 694894
rect 587498 694658 587582 694894
rect 587818 694658 592650 694894
rect -8726 694574 592650 694658
rect -8726 694338 -3894 694574
rect -3658 694338 -3574 694574
rect -3338 694338 9266 694574
rect 9502 694338 9586 694574
rect 9822 694338 45266 694574
rect 45502 694338 45586 694574
rect 45822 694338 81266 694574
rect 81502 694338 81586 694574
rect 81822 694338 117266 694574
rect 117502 694338 117586 694574
rect 117822 694338 153266 694574
rect 153502 694338 153586 694574
rect 153822 694338 189266 694574
rect 189502 694338 189586 694574
rect 189822 694338 225266 694574
rect 225502 694338 225586 694574
rect 225822 694338 261266 694574
rect 261502 694338 261586 694574
rect 261822 694338 297266 694574
rect 297502 694338 297586 694574
rect 297822 694338 333266 694574
rect 333502 694338 333586 694574
rect 333822 694338 369266 694574
rect 369502 694338 369586 694574
rect 369822 694338 405266 694574
rect 405502 694338 405586 694574
rect 405822 694338 441266 694574
rect 441502 694338 441586 694574
rect 441822 694338 477266 694574
rect 477502 694338 477586 694574
rect 477822 694338 513266 694574
rect 513502 694338 513586 694574
rect 513822 694338 549266 694574
rect 549502 694338 549586 694574
rect 549822 694338 587262 694574
rect 587498 694338 587582 694574
rect 587818 694338 592650 694574
rect -8726 694306 592650 694338
rect -8726 691174 592650 691206
rect -8726 690938 -2934 691174
rect -2698 690938 -2614 691174
rect -2378 690938 5546 691174
rect 5782 690938 5866 691174
rect 6102 690938 41546 691174
rect 41782 690938 41866 691174
rect 42102 690938 77546 691174
rect 77782 690938 77866 691174
rect 78102 690938 113546 691174
rect 113782 690938 113866 691174
rect 114102 690938 149546 691174
rect 149782 690938 149866 691174
rect 150102 690938 185546 691174
rect 185782 690938 185866 691174
rect 186102 690938 221546 691174
rect 221782 690938 221866 691174
rect 222102 690938 257546 691174
rect 257782 690938 257866 691174
rect 258102 690938 293546 691174
rect 293782 690938 293866 691174
rect 294102 690938 329546 691174
rect 329782 690938 329866 691174
rect 330102 690938 365546 691174
rect 365782 690938 365866 691174
rect 366102 690938 401546 691174
rect 401782 690938 401866 691174
rect 402102 690938 437546 691174
rect 437782 690938 437866 691174
rect 438102 690938 473546 691174
rect 473782 690938 473866 691174
rect 474102 690938 509546 691174
rect 509782 690938 509866 691174
rect 510102 690938 545546 691174
rect 545782 690938 545866 691174
rect 546102 690938 581546 691174
rect 581782 690938 581866 691174
rect 582102 690938 586302 691174
rect 586538 690938 586622 691174
rect 586858 690938 592650 691174
rect -8726 690854 592650 690938
rect -8726 690618 -2934 690854
rect -2698 690618 -2614 690854
rect -2378 690618 5546 690854
rect 5782 690618 5866 690854
rect 6102 690618 41546 690854
rect 41782 690618 41866 690854
rect 42102 690618 77546 690854
rect 77782 690618 77866 690854
rect 78102 690618 113546 690854
rect 113782 690618 113866 690854
rect 114102 690618 149546 690854
rect 149782 690618 149866 690854
rect 150102 690618 185546 690854
rect 185782 690618 185866 690854
rect 186102 690618 221546 690854
rect 221782 690618 221866 690854
rect 222102 690618 257546 690854
rect 257782 690618 257866 690854
rect 258102 690618 293546 690854
rect 293782 690618 293866 690854
rect 294102 690618 329546 690854
rect 329782 690618 329866 690854
rect 330102 690618 365546 690854
rect 365782 690618 365866 690854
rect 366102 690618 401546 690854
rect 401782 690618 401866 690854
rect 402102 690618 437546 690854
rect 437782 690618 437866 690854
rect 438102 690618 473546 690854
rect 473782 690618 473866 690854
rect 474102 690618 509546 690854
rect 509782 690618 509866 690854
rect 510102 690618 545546 690854
rect 545782 690618 545866 690854
rect 546102 690618 581546 690854
rect 581782 690618 581866 690854
rect 582102 690618 586302 690854
rect 586538 690618 586622 690854
rect 586858 690618 592650 690854
rect -8726 690586 592650 690618
rect -8726 687454 592650 687486
rect -8726 687218 -1974 687454
rect -1738 687218 -1654 687454
rect -1418 687218 1826 687454
rect 2062 687218 2146 687454
rect 2382 687218 37826 687454
rect 38062 687218 38146 687454
rect 38382 687218 73826 687454
rect 74062 687218 74146 687454
rect 74382 687218 109826 687454
rect 110062 687218 110146 687454
rect 110382 687218 145826 687454
rect 146062 687218 146146 687454
rect 146382 687218 181826 687454
rect 182062 687218 182146 687454
rect 182382 687218 217826 687454
rect 218062 687218 218146 687454
rect 218382 687218 253826 687454
rect 254062 687218 254146 687454
rect 254382 687218 289826 687454
rect 290062 687218 290146 687454
rect 290382 687218 325826 687454
rect 326062 687218 326146 687454
rect 326382 687218 361826 687454
rect 362062 687218 362146 687454
rect 362382 687218 397826 687454
rect 398062 687218 398146 687454
rect 398382 687218 433826 687454
rect 434062 687218 434146 687454
rect 434382 687218 469826 687454
rect 470062 687218 470146 687454
rect 470382 687218 505826 687454
rect 506062 687218 506146 687454
rect 506382 687218 541826 687454
rect 542062 687218 542146 687454
rect 542382 687218 577826 687454
rect 578062 687218 578146 687454
rect 578382 687218 585342 687454
rect 585578 687218 585662 687454
rect 585898 687218 592650 687454
rect -8726 687134 592650 687218
rect -8726 686898 -1974 687134
rect -1738 686898 -1654 687134
rect -1418 686898 1826 687134
rect 2062 686898 2146 687134
rect 2382 686898 37826 687134
rect 38062 686898 38146 687134
rect 38382 686898 73826 687134
rect 74062 686898 74146 687134
rect 74382 686898 109826 687134
rect 110062 686898 110146 687134
rect 110382 686898 145826 687134
rect 146062 686898 146146 687134
rect 146382 686898 181826 687134
rect 182062 686898 182146 687134
rect 182382 686898 217826 687134
rect 218062 686898 218146 687134
rect 218382 686898 253826 687134
rect 254062 686898 254146 687134
rect 254382 686898 289826 687134
rect 290062 686898 290146 687134
rect 290382 686898 325826 687134
rect 326062 686898 326146 687134
rect 326382 686898 361826 687134
rect 362062 686898 362146 687134
rect 362382 686898 397826 687134
rect 398062 686898 398146 687134
rect 398382 686898 433826 687134
rect 434062 686898 434146 687134
rect 434382 686898 469826 687134
rect 470062 686898 470146 687134
rect 470382 686898 505826 687134
rect 506062 686898 506146 687134
rect 506382 686898 541826 687134
rect 542062 686898 542146 687134
rect 542382 686898 577826 687134
rect 578062 686898 578146 687134
rect 578382 686898 585342 687134
rect 585578 686898 585662 687134
rect 585898 686898 592650 687134
rect -8726 686866 592650 686898
rect -8726 677494 592650 677526
rect -8726 677258 -8694 677494
rect -8458 677258 -8374 677494
rect -8138 677258 27866 677494
rect 28102 677258 28186 677494
rect 28422 677258 63866 677494
rect 64102 677258 64186 677494
rect 64422 677258 99866 677494
rect 100102 677258 100186 677494
rect 100422 677258 135866 677494
rect 136102 677258 136186 677494
rect 136422 677258 171866 677494
rect 172102 677258 172186 677494
rect 172422 677258 207866 677494
rect 208102 677258 208186 677494
rect 208422 677258 243866 677494
rect 244102 677258 244186 677494
rect 244422 677258 279866 677494
rect 280102 677258 280186 677494
rect 280422 677258 315866 677494
rect 316102 677258 316186 677494
rect 316422 677258 351866 677494
rect 352102 677258 352186 677494
rect 352422 677258 387866 677494
rect 388102 677258 388186 677494
rect 388422 677258 423866 677494
rect 424102 677258 424186 677494
rect 424422 677258 459866 677494
rect 460102 677258 460186 677494
rect 460422 677258 495866 677494
rect 496102 677258 496186 677494
rect 496422 677258 531866 677494
rect 532102 677258 532186 677494
rect 532422 677258 567866 677494
rect 568102 677258 568186 677494
rect 568422 677258 592062 677494
rect 592298 677258 592382 677494
rect 592618 677258 592650 677494
rect -8726 677174 592650 677258
rect -8726 676938 -8694 677174
rect -8458 676938 -8374 677174
rect -8138 676938 27866 677174
rect 28102 676938 28186 677174
rect 28422 676938 63866 677174
rect 64102 676938 64186 677174
rect 64422 676938 99866 677174
rect 100102 676938 100186 677174
rect 100422 676938 135866 677174
rect 136102 676938 136186 677174
rect 136422 676938 171866 677174
rect 172102 676938 172186 677174
rect 172422 676938 207866 677174
rect 208102 676938 208186 677174
rect 208422 676938 243866 677174
rect 244102 676938 244186 677174
rect 244422 676938 279866 677174
rect 280102 676938 280186 677174
rect 280422 676938 315866 677174
rect 316102 676938 316186 677174
rect 316422 676938 351866 677174
rect 352102 676938 352186 677174
rect 352422 676938 387866 677174
rect 388102 676938 388186 677174
rect 388422 676938 423866 677174
rect 424102 676938 424186 677174
rect 424422 676938 459866 677174
rect 460102 676938 460186 677174
rect 460422 676938 495866 677174
rect 496102 676938 496186 677174
rect 496422 676938 531866 677174
rect 532102 676938 532186 677174
rect 532422 676938 567866 677174
rect 568102 676938 568186 677174
rect 568422 676938 592062 677174
rect 592298 676938 592382 677174
rect 592618 676938 592650 677174
rect -8726 676906 592650 676938
rect -8726 673774 592650 673806
rect -8726 673538 -7734 673774
rect -7498 673538 -7414 673774
rect -7178 673538 24146 673774
rect 24382 673538 24466 673774
rect 24702 673538 60146 673774
rect 60382 673538 60466 673774
rect 60702 673538 96146 673774
rect 96382 673538 96466 673774
rect 96702 673538 132146 673774
rect 132382 673538 132466 673774
rect 132702 673538 168146 673774
rect 168382 673538 168466 673774
rect 168702 673538 204146 673774
rect 204382 673538 204466 673774
rect 204702 673538 240146 673774
rect 240382 673538 240466 673774
rect 240702 673538 276146 673774
rect 276382 673538 276466 673774
rect 276702 673538 312146 673774
rect 312382 673538 312466 673774
rect 312702 673538 348146 673774
rect 348382 673538 348466 673774
rect 348702 673538 384146 673774
rect 384382 673538 384466 673774
rect 384702 673538 420146 673774
rect 420382 673538 420466 673774
rect 420702 673538 456146 673774
rect 456382 673538 456466 673774
rect 456702 673538 492146 673774
rect 492382 673538 492466 673774
rect 492702 673538 528146 673774
rect 528382 673538 528466 673774
rect 528702 673538 564146 673774
rect 564382 673538 564466 673774
rect 564702 673538 591102 673774
rect 591338 673538 591422 673774
rect 591658 673538 592650 673774
rect -8726 673454 592650 673538
rect -8726 673218 -7734 673454
rect -7498 673218 -7414 673454
rect -7178 673218 24146 673454
rect 24382 673218 24466 673454
rect 24702 673218 60146 673454
rect 60382 673218 60466 673454
rect 60702 673218 96146 673454
rect 96382 673218 96466 673454
rect 96702 673218 132146 673454
rect 132382 673218 132466 673454
rect 132702 673218 168146 673454
rect 168382 673218 168466 673454
rect 168702 673218 204146 673454
rect 204382 673218 204466 673454
rect 204702 673218 240146 673454
rect 240382 673218 240466 673454
rect 240702 673218 276146 673454
rect 276382 673218 276466 673454
rect 276702 673218 312146 673454
rect 312382 673218 312466 673454
rect 312702 673218 348146 673454
rect 348382 673218 348466 673454
rect 348702 673218 384146 673454
rect 384382 673218 384466 673454
rect 384702 673218 420146 673454
rect 420382 673218 420466 673454
rect 420702 673218 456146 673454
rect 456382 673218 456466 673454
rect 456702 673218 492146 673454
rect 492382 673218 492466 673454
rect 492702 673218 528146 673454
rect 528382 673218 528466 673454
rect 528702 673218 564146 673454
rect 564382 673218 564466 673454
rect 564702 673218 591102 673454
rect 591338 673218 591422 673454
rect 591658 673218 592650 673454
rect -8726 673186 592650 673218
rect -8726 670054 592650 670086
rect -8726 669818 -6774 670054
rect -6538 669818 -6454 670054
rect -6218 669818 20426 670054
rect 20662 669818 20746 670054
rect 20982 669818 56426 670054
rect 56662 669818 56746 670054
rect 56982 669818 92426 670054
rect 92662 669818 92746 670054
rect 92982 669818 128426 670054
rect 128662 669818 128746 670054
rect 128982 669818 164426 670054
rect 164662 669818 164746 670054
rect 164982 669818 200426 670054
rect 200662 669818 200746 670054
rect 200982 669818 236426 670054
rect 236662 669818 236746 670054
rect 236982 669818 272426 670054
rect 272662 669818 272746 670054
rect 272982 669818 308426 670054
rect 308662 669818 308746 670054
rect 308982 669818 344426 670054
rect 344662 669818 344746 670054
rect 344982 669818 380426 670054
rect 380662 669818 380746 670054
rect 380982 669818 416426 670054
rect 416662 669818 416746 670054
rect 416982 669818 452426 670054
rect 452662 669818 452746 670054
rect 452982 669818 488426 670054
rect 488662 669818 488746 670054
rect 488982 669818 524426 670054
rect 524662 669818 524746 670054
rect 524982 669818 560426 670054
rect 560662 669818 560746 670054
rect 560982 669818 590142 670054
rect 590378 669818 590462 670054
rect 590698 669818 592650 670054
rect -8726 669734 592650 669818
rect -8726 669498 -6774 669734
rect -6538 669498 -6454 669734
rect -6218 669498 20426 669734
rect 20662 669498 20746 669734
rect 20982 669498 56426 669734
rect 56662 669498 56746 669734
rect 56982 669498 92426 669734
rect 92662 669498 92746 669734
rect 92982 669498 128426 669734
rect 128662 669498 128746 669734
rect 128982 669498 164426 669734
rect 164662 669498 164746 669734
rect 164982 669498 200426 669734
rect 200662 669498 200746 669734
rect 200982 669498 236426 669734
rect 236662 669498 236746 669734
rect 236982 669498 272426 669734
rect 272662 669498 272746 669734
rect 272982 669498 308426 669734
rect 308662 669498 308746 669734
rect 308982 669498 344426 669734
rect 344662 669498 344746 669734
rect 344982 669498 380426 669734
rect 380662 669498 380746 669734
rect 380982 669498 416426 669734
rect 416662 669498 416746 669734
rect 416982 669498 452426 669734
rect 452662 669498 452746 669734
rect 452982 669498 488426 669734
rect 488662 669498 488746 669734
rect 488982 669498 524426 669734
rect 524662 669498 524746 669734
rect 524982 669498 560426 669734
rect 560662 669498 560746 669734
rect 560982 669498 590142 669734
rect 590378 669498 590462 669734
rect 590698 669498 592650 669734
rect -8726 669466 592650 669498
rect -8726 666334 592650 666366
rect -8726 666098 -5814 666334
rect -5578 666098 -5494 666334
rect -5258 666098 16706 666334
rect 16942 666098 17026 666334
rect 17262 666098 52706 666334
rect 52942 666098 53026 666334
rect 53262 666098 88706 666334
rect 88942 666098 89026 666334
rect 89262 666098 124706 666334
rect 124942 666098 125026 666334
rect 125262 666098 160706 666334
rect 160942 666098 161026 666334
rect 161262 666098 196706 666334
rect 196942 666098 197026 666334
rect 197262 666098 232706 666334
rect 232942 666098 233026 666334
rect 233262 666098 268706 666334
rect 268942 666098 269026 666334
rect 269262 666098 304706 666334
rect 304942 666098 305026 666334
rect 305262 666098 340706 666334
rect 340942 666098 341026 666334
rect 341262 666098 376706 666334
rect 376942 666098 377026 666334
rect 377262 666098 412706 666334
rect 412942 666098 413026 666334
rect 413262 666098 448706 666334
rect 448942 666098 449026 666334
rect 449262 666098 484706 666334
rect 484942 666098 485026 666334
rect 485262 666098 520706 666334
rect 520942 666098 521026 666334
rect 521262 666098 556706 666334
rect 556942 666098 557026 666334
rect 557262 666098 589182 666334
rect 589418 666098 589502 666334
rect 589738 666098 592650 666334
rect -8726 666014 592650 666098
rect -8726 665778 -5814 666014
rect -5578 665778 -5494 666014
rect -5258 665778 16706 666014
rect 16942 665778 17026 666014
rect 17262 665778 52706 666014
rect 52942 665778 53026 666014
rect 53262 665778 88706 666014
rect 88942 665778 89026 666014
rect 89262 665778 124706 666014
rect 124942 665778 125026 666014
rect 125262 665778 160706 666014
rect 160942 665778 161026 666014
rect 161262 665778 196706 666014
rect 196942 665778 197026 666014
rect 197262 665778 232706 666014
rect 232942 665778 233026 666014
rect 233262 665778 268706 666014
rect 268942 665778 269026 666014
rect 269262 665778 304706 666014
rect 304942 665778 305026 666014
rect 305262 665778 340706 666014
rect 340942 665778 341026 666014
rect 341262 665778 376706 666014
rect 376942 665778 377026 666014
rect 377262 665778 412706 666014
rect 412942 665778 413026 666014
rect 413262 665778 448706 666014
rect 448942 665778 449026 666014
rect 449262 665778 484706 666014
rect 484942 665778 485026 666014
rect 485262 665778 520706 666014
rect 520942 665778 521026 666014
rect 521262 665778 556706 666014
rect 556942 665778 557026 666014
rect 557262 665778 589182 666014
rect 589418 665778 589502 666014
rect 589738 665778 592650 666014
rect -8726 665746 592650 665778
rect -8726 662614 592650 662646
rect -8726 662378 -4854 662614
rect -4618 662378 -4534 662614
rect -4298 662378 12986 662614
rect 13222 662378 13306 662614
rect 13542 662378 48986 662614
rect 49222 662378 49306 662614
rect 49542 662378 84986 662614
rect 85222 662378 85306 662614
rect 85542 662378 120986 662614
rect 121222 662378 121306 662614
rect 121542 662378 156986 662614
rect 157222 662378 157306 662614
rect 157542 662378 192986 662614
rect 193222 662378 193306 662614
rect 193542 662378 228986 662614
rect 229222 662378 229306 662614
rect 229542 662378 264986 662614
rect 265222 662378 265306 662614
rect 265542 662378 300986 662614
rect 301222 662378 301306 662614
rect 301542 662378 336986 662614
rect 337222 662378 337306 662614
rect 337542 662378 372986 662614
rect 373222 662378 373306 662614
rect 373542 662378 408986 662614
rect 409222 662378 409306 662614
rect 409542 662378 444986 662614
rect 445222 662378 445306 662614
rect 445542 662378 480986 662614
rect 481222 662378 481306 662614
rect 481542 662378 516986 662614
rect 517222 662378 517306 662614
rect 517542 662378 552986 662614
rect 553222 662378 553306 662614
rect 553542 662378 588222 662614
rect 588458 662378 588542 662614
rect 588778 662378 592650 662614
rect -8726 662294 592650 662378
rect -8726 662058 -4854 662294
rect -4618 662058 -4534 662294
rect -4298 662058 12986 662294
rect 13222 662058 13306 662294
rect 13542 662058 48986 662294
rect 49222 662058 49306 662294
rect 49542 662058 84986 662294
rect 85222 662058 85306 662294
rect 85542 662058 120986 662294
rect 121222 662058 121306 662294
rect 121542 662058 156986 662294
rect 157222 662058 157306 662294
rect 157542 662058 192986 662294
rect 193222 662058 193306 662294
rect 193542 662058 228986 662294
rect 229222 662058 229306 662294
rect 229542 662058 264986 662294
rect 265222 662058 265306 662294
rect 265542 662058 300986 662294
rect 301222 662058 301306 662294
rect 301542 662058 336986 662294
rect 337222 662058 337306 662294
rect 337542 662058 372986 662294
rect 373222 662058 373306 662294
rect 373542 662058 408986 662294
rect 409222 662058 409306 662294
rect 409542 662058 444986 662294
rect 445222 662058 445306 662294
rect 445542 662058 480986 662294
rect 481222 662058 481306 662294
rect 481542 662058 516986 662294
rect 517222 662058 517306 662294
rect 517542 662058 552986 662294
rect 553222 662058 553306 662294
rect 553542 662058 588222 662294
rect 588458 662058 588542 662294
rect 588778 662058 592650 662294
rect -8726 662026 592650 662058
rect -8726 658894 592650 658926
rect -8726 658658 -3894 658894
rect -3658 658658 -3574 658894
rect -3338 658658 9266 658894
rect 9502 658658 9586 658894
rect 9822 658658 45266 658894
rect 45502 658658 45586 658894
rect 45822 658658 81266 658894
rect 81502 658658 81586 658894
rect 81822 658658 117266 658894
rect 117502 658658 117586 658894
rect 117822 658658 153266 658894
rect 153502 658658 153586 658894
rect 153822 658658 189266 658894
rect 189502 658658 189586 658894
rect 189822 658658 225266 658894
rect 225502 658658 225586 658894
rect 225822 658658 261266 658894
rect 261502 658658 261586 658894
rect 261822 658658 297266 658894
rect 297502 658658 297586 658894
rect 297822 658658 333266 658894
rect 333502 658658 333586 658894
rect 333822 658658 369266 658894
rect 369502 658658 369586 658894
rect 369822 658658 405266 658894
rect 405502 658658 405586 658894
rect 405822 658658 441266 658894
rect 441502 658658 441586 658894
rect 441822 658658 477266 658894
rect 477502 658658 477586 658894
rect 477822 658658 513266 658894
rect 513502 658658 513586 658894
rect 513822 658658 549266 658894
rect 549502 658658 549586 658894
rect 549822 658658 587262 658894
rect 587498 658658 587582 658894
rect 587818 658658 592650 658894
rect -8726 658574 592650 658658
rect -8726 658338 -3894 658574
rect -3658 658338 -3574 658574
rect -3338 658338 9266 658574
rect 9502 658338 9586 658574
rect 9822 658338 45266 658574
rect 45502 658338 45586 658574
rect 45822 658338 81266 658574
rect 81502 658338 81586 658574
rect 81822 658338 117266 658574
rect 117502 658338 117586 658574
rect 117822 658338 153266 658574
rect 153502 658338 153586 658574
rect 153822 658338 189266 658574
rect 189502 658338 189586 658574
rect 189822 658338 225266 658574
rect 225502 658338 225586 658574
rect 225822 658338 261266 658574
rect 261502 658338 261586 658574
rect 261822 658338 297266 658574
rect 297502 658338 297586 658574
rect 297822 658338 333266 658574
rect 333502 658338 333586 658574
rect 333822 658338 369266 658574
rect 369502 658338 369586 658574
rect 369822 658338 405266 658574
rect 405502 658338 405586 658574
rect 405822 658338 441266 658574
rect 441502 658338 441586 658574
rect 441822 658338 477266 658574
rect 477502 658338 477586 658574
rect 477822 658338 513266 658574
rect 513502 658338 513586 658574
rect 513822 658338 549266 658574
rect 549502 658338 549586 658574
rect 549822 658338 587262 658574
rect 587498 658338 587582 658574
rect 587818 658338 592650 658574
rect -8726 658306 592650 658338
rect -8726 655174 592650 655206
rect -8726 654938 -2934 655174
rect -2698 654938 -2614 655174
rect -2378 654938 5546 655174
rect 5782 654938 5866 655174
rect 6102 654938 41546 655174
rect 41782 654938 41866 655174
rect 42102 654938 77546 655174
rect 77782 654938 77866 655174
rect 78102 654938 113546 655174
rect 113782 654938 113866 655174
rect 114102 654938 149546 655174
rect 149782 654938 149866 655174
rect 150102 654938 185546 655174
rect 185782 654938 185866 655174
rect 186102 654938 221546 655174
rect 221782 654938 221866 655174
rect 222102 654938 257546 655174
rect 257782 654938 257866 655174
rect 258102 654938 293546 655174
rect 293782 654938 293866 655174
rect 294102 654938 329546 655174
rect 329782 654938 329866 655174
rect 330102 654938 365546 655174
rect 365782 654938 365866 655174
rect 366102 654938 401546 655174
rect 401782 654938 401866 655174
rect 402102 654938 437546 655174
rect 437782 654938 437866 655174
rect 438102 654938 473546 655174
rect 473782 654938 473866 655174
rect 474102 654938 509546 655174
rect 509782 654938 509866 655174
rect 510102 654938 545546 655174
rect 545782 654938 545866 655174
rect 546102 654938 581546 655174
rect 581782 654938 581866 655174
rect 582102 654938 586302 655174
rect 586538 654938 586622 655174
rect 586858 654938 592650 655174
rect -8726 654854 592650 654938
rect -8726 654618 -2934 654854
rect -2698 654618 -2614 654854
rect -2378 654618 5546 654854
rect 5782 654618 5866 654854
rect 6102 654618 41546 654854
rect 41782 654618 41866 654854
rect 42102 654618 77546 654854
rect 77782 654618 77866 654854
rect 78102 654618 113546 654854
rect 113782 654618 113866 654854
rect 114102 654618 149546 654854
rect 149782 654618 149866 654854
rect 150102 654618 185546 654854
rect 185782 654618 185866 654854
rect 186102 654618 221546 654854
rect 221782 654618 221866 654854
rect 222102 654618 257546 654854
rect 257782 654618 257866 654854
rect 258102 654618 293546 654854
rect 293782 654618 293866 654854
rect 294102 654618 329546 654854
rect 329782 654618 329866 654854
rect 330102 654618 365546 654854
rect 365782 654618 365866 654854
rect 366102 654618 401546 654854
rect 401782 654618 401866 654854
rect 402102 654618 437546 654854
rect 437782 654618 437866 654854
rect 438102 654618 473546 654854
rect 473782 654618 473866 654854
rect 474102 654618 509546 654854
rect 509782 654618 509866 654854
rect 510102 654618 545546 654854
rect 545782 654618 545866 654854
rect 546102 654618 581546 654854
rect 581782 654618 581866 654854
rect 582102 654618 586302 654854
rect 586538 654618 586622 654854
rect 586858 654618 592650 654854
rect -8726 654586 592650 654618
rect -8726 651454 592650 651486
rect -8726 651218 -1974 651454
rect -1738 651218 -1654 651454
rect -1418 651218 1826 651454
rect 2062 651218 2146 651454
rect 2382 651218 37826 651454
rect 38062 651218 38146 651454
rect 38382 651218 73826 651454
rect 74062 651218 74146 651454
rect 74382 651218 109826 651454
rect 110062 651218 110146 651454
rect 110382 651218 145826 651454
rect 146062 651218 146146 651454
rect 146382 651218 181826 651454
rect 182062 651218 182146 651454
rect 182382 651218 217826 651454
rect 218062 651218 218146 651454
rect 218382 651218 253826 651454
rect 254062 651218 254146 651454
rect 254382 651218 289826 651454
rect 290062 651218 290146 651454
rect 290382 651218 325826 651454
rect 326062 651218 326146 651454
rect 326382 651218 361826 651454
rect 362062 651218 362146 651454
rect 362382 651218 397826 651454
rect 398062 651218 398146 651454
rect 398382 651218 433826 651454
rect 434062 651218 434146 651454
rect 434382 651218 469826 651454
rect 470062 651218 470146 651454
rect 470382 651218 505826 651454
rect 506062 651218 506146 651454
rect 506382 651218 541826 651454
rect 542062 651218 542146 651454
rect 542382 651218 577826 651454
rect 578062 651218 578146 651454
rect 578382 651218 585342 651454
rect 585578 651218 585662 651454
rect 585898 651218 592650 651454
rect -8726 651134 592650 651218
rect -8726 650898 -1974 651134
rect -1738 650898 -1654 651134
rect -1418 650898 1826 651134
rect 2062 650898 2146 651134
rect 2382 650898 37826 651134
rect 38062 650898 38146 651134
rect 38382 650898 73826 651134
rect 74062 650898 74146 651134
rect 74382 650898 109826 651134
rect 110062 650898 110146 651134
rect 110382 650898 145826 651134
rect 146062 650898 146146 651134
rect 146382 650898 181826 651134
rect 182062 650898 182146 651134
rect 182382 650898 217826 651134
rect 218062 650898 218146 651134
rect 218382 650898 253826 651134
rect 254062 650898 254146 651134
rect 254382 650898 289826 651134
rect 290062 650898 290146 651134
rect 290382 650898 325826 651134
rect 326062 650898 326146 651134
rect 326382 650898 361826 651134
rect 362062 650898 362146 651134
rect 362382 650898 397826 651134
rect 398062 650898 398146 651134
rect 398382 650898 433826 651134
rect 434062 650898 434146 651134
rect 434382 650898 469826 651134
rect 470062 650898 470146 651134
rect 470382 650898 505826 651134
rect 506062 650898 506146 651134
rect 506382 650898 541826 651134
rect 542062 650898 542146 651134
rect 542382 650898 577826 651134
rect 578062 650898 578146 651134
rect 578382 650898 585342 651134
rect 585578 650898 585662 651134
rect 585898 650898 592650 651134
rect -8726 650866 592650 650898
rect -8726 641494 592650 641526
rect -8726 641258 -8694 641494
rect -8458 641258 -8374 641494
rect -8138 641258 27866 641494
rect 28102 641258 28186 641494
rect 28422 641258 63866 641494
rect 64102 641258 64186 641494
rect 64422 641258 99866 641494
rect 100102 641258 100186 641494
rect 100422 641258 135866 641494
rect 136102 641258 136186 641494
rect 136422 641258 171866 641494
rect 172102 641258 172186 641494
rect 172422 641258 207866 641494
rect 208102 641258 208186 641494
rect 208422 641258 243866 641494
rect 244102 641258 244186 641494
rect 244422 641258 567866 641494
rect 568102 641258 568186 641494
rect 568422 641258 592062 641494
rect 592298 641258 592382 641494
rect 592618 641258 592650 641494
rect -8726 641174 592650 641258
rect -8726 640938 -8694 641174
rect -8458 640938 -8374 641174
rect -8138 640938 27866 641174
rect 28102 640938 28186 641174
rect 28422 640938 63866 641174
rect 64102 640938 64186 641174
rect 64422 640938 99866 641174
rect 100102 640938 100186 641174
rect 100422 640938 135866 641174
rect 136102 640938 136186 641174
rect 136422 640938 171866 641174
rect 172102 640938 172186 641174
rect 172422 640938 207866 641174
rect 208102 640938 208186 641174
rect 208422 640938 243866 641174
rect 244102 640938 244186 641174
rect 244422 640938 567866 641174
rect 568102 640938 568186 641174
rect 568422 640938 592062 641174
rect 592298 640938 592382 641174
rect 592618 640938 592650 641174
rect -8726 640906 592650 640938
rect -8726 637774 592650 637806
rect -8726 637538 -7734 637774
rect -7498 637538 -7414 637774
rect -7178 637538 24146 637774
rect 24382 637538 24466 637774
rect 24702 637538 60146 637774
rect 60382 637538 60466 637774
rect 60702 637538 96146 637774
rect 96382 637538 96466 637774
rect 96702 637538 132146 637774
rect 132382 637538 132466 637774
rect 132702 637538 168146 637774
rect 168382 637538 168466 637774
rect 168702 637538 204146 637774
rect 204382 637538 204466 637774
rect 204702 637538 240146 637774
rect 240382 637538 240466 637774
rect 240702 637538 564146 637774
rect 564382 637538 564466 637774
rect 564702 637538 591102 637774
rect 591338 637538 591422 637774
rect 591658 637538 592650 637774
rect -8726 637454 592650 637538
rect -8726 637218 -7734 637454
rect -7498 637218 -7414 637454
rect -7178 637218 24146 637454
rect 24382 637218 24466 637454
rect 24702 637218 60146 637454
rect 60382 637218 60466 637454
rect 60702 637218 96146 637454
rect 96382 637218 96466 637454
rect 96702 637218 132146 637454
rect 132382 637218 132466 637454
rect 132702 637218 168146 637454
rect 168382 637218 168466 637454
rect 168702 637218 204146 637454
rect 204382 637218 204466 637454
rect 204702 637218 240146 637454
rect 240382 637218 240466 637454
rect 240702 637218 564146 637454
rect 564382 637218 564466 637454
rect 564702 637218 591102 637454
rect 591338 637218 591422 637454
rect 591658 637218 592650 637454
rect -8726 637186 592650 637218
rect -8726 634054 592650 634086
rect -8726 633818 -6774 634054
rect -6538 633818 -6454 634054
rect -6218 633818 20426 634054
rect 20662 633818 20746 634054
rect 20982 633818 56426 634054
rect 56662 633818 56746 634054
rect 56982 633818 92426 634054
rect 92662 633818 92746 634054
rect 92982 633818 128426 634054
rect 128662 633818 128746 634054
rect 128982 633818 164426 634054
rect 164662 633818 164746 634054
rect 164982 633818 200426 634054
rect 200662 633818 200746 634054
rect 200982 633818 236426 634054
rect 236662 633818 236746 634054
rect 236982 633818 560426 634054
rect 560662 633818 560746 634054
rect 560982 633818 590142 634054
rect 590378 633818 590462 634054
rect 590698 633818 592650 634054
rect -8726 633734 592650 633818
rect -8726 633498 -6774 633734
rect -6538 633498 -6454 633734
rect -6218 633498 20426 633734
rect 20662 633498 20746 633734
rect 20982 633498 56426 633734
rect 56662 633498 56746 633734
rect 56982 633498 92426 633734
rect 92662 633498 92746 633734
rect 92982 633498 128426 633734
rect 128662 633498 128746 633734
rect 128982 633498 164426 633734
rect 164662 633498 164746 633734
rect 164982 633498 200426 633734
rect 200662 633498 200746 633734
rect 200982 633498 236426 633734
rect 236662 633498 236746 633734
rect 236982 633498 560426 633734
rect 560662 633498 560746 633734
rect 560982 633498 590142 633734
rect 590378 633498 590462 633734
rect 590698 633498 592650 633734
rect -8726 633466 592650 633498
rect -8726 630334 592650 630366
rect -8726 630098 -5814 630334
rect -5578 630098 -5494 630334
rect -5258 630098 16706 630334
rect 16942 630098 17026 630334
rect 17262 630098 52706 630334
rect 52942 630098 53026 630334
rect 53262 630098 88706 630334
rect 88942 630098 89026 630334
rect 89262 630098 124706 630334
rect 124942 630098 125026 630334
rect 125262 630098 160706 630334
rect 160942 630098 161026 630334
rect 161262 630098 196706 630334
rect 196942 630098 197026 630334
rect 197262 630098 232706 630334
rect 232942 630098 233026 630334
rect 233262 630098 556706 630334
rect 556942 630098 557026 630334
rect 557262 630098 589182 630334
rect 589418 630098 589502 630334
rect 589738 630098 592650 630334
rect -8726 630014 592650 630098
rect -8726 629778 -5814 630014
rect -5578 629778 -5494 630014
rect -5258 629778 16706 630014
rect 16942 629778 17026 630014
rect 17262 629778 52706 630014
rect 52942 629778 53026 630014
rect 53262 629778 88706 630014
rect 88942 629778 89026 630014
rect 89262 629778 124706 630014
rect 124942 629778 125026 630014
rect 125262 629778 160706 630014
rect 160942 629778 161026 630014
rect 161262 629778 196706 630014
rect 196942 629778 197026 630014
rect 197262 629778 232706 630014
rect 232942 629778 233026 630014
rect 233262 629778 556706 630014
rect 556942 629778 557026 630014
rect 557262 629778 589182 630014
rect 589418 629778 589502 630014
rect 589738 629778 592650 630014
rect -8726 629746 592650 629778
rect -8726 626614 592650 626646
rect -8726 626378 -4854 626614
rect -4618 626378 -4534 626614
rect -4298 626378 12986 626614
rect 13222 626378 13306 626614
rect 13542 626378 48986 626614
rect 49222 626378 49306 626614
rect 49542 626378 84986 626614
rect 85222 626378 85306 626614
rect 85542 626378 120986 626614
rect 121222 626378 121306 626614
rect 121542 626378 156986 626614
rect 157222 626378 157306 626614
rect 157542 626378 192986 626614
rect 193222 626378 193306 626614
rect 193542 626378 228986 626614
rect 229222 626378 229306 626614
rect 229542 626378 552986 626614
rect 553222 626378 553306 626614
rect 553542 626378 588222 626614
rect 588458 626378 588542 626614
rect 588778 626378 592650 626614
rect -8726 626294 592650 626378
rect -8726 626058 -4854 626294
rect -4618 626058 -4534 626294
rect -4298 626058 12986 626294
rect 13222 626058 13306 626294
rect 13542 626058 48986 626294
rect 49222 626058 49306 626294
rect 49542 626058 84986 626294
rect 85222 626058 85306 626294
rect 85542 626058 120986 626294
rect 121222 626058 121306 626294
rect 121542 626058 156986 626294
rect 157222 626058 157306 626294
rect 157542 626058 192986 626294
rect 193222 626058 193306 626294
rect 193542 626058 228986 626294
rect 229222 626058 229306 626294
rect 229542 626058 552986 626294
rect 553222 626058 553306 626294
rect 553542 626058 588222 626294
rect 588458 626058 588542 626294
rect 588778 626058 592650 626294
rect -8726 626026 592650 626058
rect -8726 622894 592650 622926
rect -8726 622658 -3894 622894
rect -3658 622658 -3574 622894
rect -3338 622658 9266 622894
rect 9502 622658 9586 622894
rect 9822 622658 45266 622894
rect 45502 622658 45586 622894
rect 45822 622658 81266 622894
rect 81502 622658 81586 622894
rect 81822 622658 117266 622894
rect 117502 622658 117586 622894
rect 117822 622658 153266 622894
rect 153502 622658 153586 622894
rect 153822 622658 189266 622894
rect 189502 622658 189586 622894
rect 189822 622658 225266 622894
rect 225502 622658 225586 622894
rect 225822 622658 587262 622894
rect 587498 622658 587582 622894
rect 587818 622658 592650 622894
rect -8726 622574 592650 622658
rect -8726 622338 -3894 622574
rect -3658 622338 -3574 622574
rect -3338 622338 9266 622574
rect 9502 622338 9586 622574
rect 9822 622338 45266 622574
rect 45502 622338 45586 622574
rect 45822 622338 81266 622574
rect 81502 622338 81586 622574
rect 81822 622338 117266 622574
rect 117502 622338 117586 622574
rect 117822 622338 153266 622574
rect 153502 622338 153586 622574
rect 153822 622338 189266 622574
rect 189502 622338 189586 622574
rect 189822 622338 225266 622574
rect 225502 622338 225586 622574
rect 225822 622338 587262 622574
rect 587498 622338 587582 622574
rect 587818 622338 592650 622574
rect -8726 622306 592650 622338
rect -8726 619174 592650 619206
rect -8726 618938 -2934 619174
rect -2698 618938 -2614 619174
rect -2378 618938 5546 619174
rect 5782 618938 5866 619174
rect 6102 618938 41546 619174
rect 41782 618938 41866 619174
rect 42102 618938 77546 619174
rect 77782 618938 77866 619174
rect 78102 618938 113546 619174
rect 113782 618938 113866 619174
rect 114102 618938 149546 619174
rect 149782 618938 149866 619174
rect 150102 618938 185546 619174
rect 185782 618938 185866 619174
rect 186102 618938 221546 619174
rect 221782 618938 221866 619174
rect 222102 618938 273210 619174
rect 273446 618938 303930 619174
rect 304166 618938 334650 619174
rect 334886 618938 365370 619174
rect 365606 618938 396090 619174
rect 396326 618938 426810 619174
rect 427046 618938 457530 619174
rect 457766 618938 488250 619174
rect 488486 618938 518970 619174
rect 519206 618938 545546 619174
rect 545782 618938 545866 619174
rect 546102 618938 549690 619174
rect 549926 618938 581546 619174
rect 581782 618938 581866 619174
rect 582102 618938 586302 619174
rect 586538 618938 586622 619174
rect 586858 618938 592650 619174
rect -8726 618854 592650 618938
rect -8726 618618 -2934 618854
rect -2698 618618 -2614 618854
rect -2378 618618 5546 618854
rect 5782 618618 5866 618854
rect 6102 618618 41546 618854
rect 41782 618618 41866 618854
rect 42102 618618 77546 618854
rect 77782 618618 77866 618854
rect 78102 618618 113546 618854
rect 113782 618618 113866 618854
rect 114102 618618 149546 618854
rect 149782 618618 149866 618854
rect 150102 618618 185546 618854
rect 185782 618618 185866 618854
rect 186102 618618 221546 618854
rect 221782 618618 221866 618854
rect 222102 618618 273210 618854
rect 273446 618618 303930 618854
rect 304166 618618 334650 618854
rect 334886 618618 365370 618854
rect 365606 618618 396090 618854
rect 396326 618618 426810 618854
rect 427046 618618 457530 618854
rect 457766 618618 488250 618854
rect 488486 618618 518970 618854
rect 519206 618618 545546 618854
rect 545782 618618 545866 618854
rect 546102 618618 549690 618854
rect 549926 618618 581546 618854
rect 581782 618618 581866 618854
rect 582102 618618 586302 618854
rect 586538 618618 586622 618854
rect 586858 618618 592650 618854
rect -8726 618586 592650 618618
rect -8726 615454 592650 615486
rect -8726 615218 -1974 615454
rect -1738 615218 -1654 615454
rect -1418 615218 1826 615454
rect 2062 615218 2146 615454
rect 2382 615218 37826 615454
rect 38062 615218 38146 615454
rect 38382 615218 73826 615454
rect 74062 615218 74146 615454
rect 74382 615218 109826 615454
rect 110062 615218 110146 615454
rect 110382 615218 145826 615454
rect 146062 615218 146146 615454
rect 146382 615218 181826 615454
rect 182062 615218 182146 615454
rect 182382 615218 217826 615454
rect 218062 615218 218146 615454
rect 218382 615218 253826 615454
rect 254062 615218 254146 615454
rect 254382 615218 257850 615454
rect 258086 615218 288570 615454
rect 288806 615218 319290 615454
rect 319526 615218 350010 615454
rect 350246 615218 380730 615454
rect 380966 615218 411450 615454
rect 411686 615218 442170 615454
rect 442406 615218 472890 615454
rect 473126 615218 503610 615454
rect 503846 615218 534330 615454
rect 534566 615218 541826 615454
rect 542062 615218 542146 615454
rect 542382 615218 565050 615454
rect 565286 615218 577826 615454
rect 578062 615218 578146 615454
rect 578382 615218 585342 615454
rect 585578 615218 585662 615454
rect 585898 615218 592650 615454
rect -8726 615134 592650 615218
rect -8726 614898 -1974 615134
rect -1738 614898 -1654 615134
rect -1418 614898 1826 615134
rect 2062 614898 2146 615134
rect 2382 614898 37826 615134
rect 38062 614898 38146 615134
rect 38382 614898 73826 615134
rect 74062 614898 74146 615134
rect 74382 614898 109826 615134
rect 110062 614898 110146 615134
rect 110382 614898 145826 615134
rect 146062 614898 146146 615134
rect 146382 614898 181826 615134
rect 182062 614898 182146 615134
rect 182382 614898 217826 615134
rect 218062 614898 218146 615134
rect 218382 614898 253826 615134
rect 254062 614898 254146 615134
rect 254382 614898 257850 615134
rect 258086 614898 288570 615134
rect 288806 614898 319290 615134
rect 319526 614898 350010 615134
rect 350246 614898 380730 615134
rect 380966 614898 411450 615134
rect 411686 614898 442170 615134
rect 442406 614898 472890 615134
rect 473126 614898 503610 615134
rect 503846 614898 534330 615134
rect 534566 614898 541826 615134
rect 542062 614898 542146 615134
rect 542382 614898 565050 615134
rect 565286 614898 577826 615134
rect 578062 614898 578146 615134
rect 578382 614898 585342 615134
rect 585578 614898 585662 615134
rect 585898 614898 592650 615134
rect -8726 614866 592650 614898
rect -8726 605494 592650 605526
rect -8726 605258 -8694 605494
rect -8458 605258 -8374 605494
rect -8138 605258 27866 605494
rect 28102 605258 28186 605494
rect 28422 605258 63866 605494
rect 64102 605258 64186 605494
rect 64422 605258 99866 605494
rect 100102 605258 100186 605494
rect 100422 605258 135866 605494
rect 136102 605258 136186 605494
rect 136422 605258 171866 605494
rect 172102 605258 172186 605494
rect 172422 605258 207866 605494
rect 208102 605258 208186 605494
rect 208422 605258 243866 605494
rect 244102 605258 244186 605494
rect 244422 605258 567866 605494
rect 568102 605258 568186 605494
rect 568422 605258 592062 605494
rect 592298 605258 592382 605494
rect 592618 605258 592650 605494
rect -8726 605174 592650 605258
rect -8726 604938 -8694 605174
rect -8458 604938 -8374 605174
rect -8138 604938 27866 605174
rect 28102 604938 28186 605174
rect 28422 604938 63866 605174
rect 64102 604938 64186 605174
rect 64422 604938 99866 605174
rect 100102 604938 100186 605174
rect 100422 604938 135866 605174
rect 136102 604938 136186 605174
rect 136422 604938 171866 605174
rect 172102 604938 172186 605174
rect 172422 604938 207866 605174
rect 208102 604938 208186 605174
rect 208422 604938 243866 605174
rect 244102 604938 244186 605174
rect 244422 604938 567866 605174
rect 568102 604938 568186 605174
rect 568422 604938 592062 605174
rect 592298 604938 592382 605174
rect 592618 604938 592650 605174
rect -8726 604906 592650 604938
rect -8726 601774 592650 601806
rect -8726 601538 -7734 601774
rect -7498 601538 -7414 601774
rect -7178 601538 24146 601774
rect 24382 601538 24466 601774
rect 24702 601538 60146 601774
rect 60382 601538 60466 601774
rect 60702 601538 96146 601774
rect 96382 601538 96466 601774
rect 96702 601538 132146 601774
rect 132382 601538 132466 601774
rect 132702 601538 168146 601774
rect 168382 601538 168466 601774
rect 168702 601538 204146 601774
rect 204382 601538 204466 601774
rect 204702 601538 240146 601774
rect 240382 601538 240466 601774
rect 240702 601538 564146 601774
rect 564382 601538 564466 601774
rect 564702 601538 591102 601774
rect 591338 601538 591422 601774
rect 591658 601538 592650 601774
rect -8726 601454 592650 601538
rect -8726 601218 -7734 601454
rect -7498 601218 -7414 601454
rect -7178 601218 24146 601454
rect 24382 601218 24466 601454
rect 24702 601218 60146 601454
rect 60382 601218 60466 601454
rect 60702 601218 96146 601454
rect 96382 601218 96466 601454
rect 96702 601218 132146 601454
rect 132382 601218 132466 601454
rect 132702 601218 168146 601454
rect 168382 601218 168466 601454
rect 168702 601218 204146 601454
rect 204382 601218 204466 601454
rect 204702 601218 240146 601454
rect 240382 601218 240466 601454
rect 240702 601218 564146 601454
rect 564382 601218 564466 601454
rect 564702 601218 591102 601454
rect 591338 601218 591422 601454
rect 591658 601218 592650 601454
rect -8726 601186 592650 601218
rect -8726 598054 592650 598086
rect -8726 597818 -6774 598054
rect -6538 597818 -6454 598054
rect -6218 597818 20426 598054
rect 20662 597818 20746 598054
rect 20982 597818 56426 598054
rect 56662 597818 56746 598054
rect 56982 597818 92426 598054
rect 92662 597818 92746 598054
rect 92982 597818 128426 598054
rect 128662 597818 128746 598054
rect 128982 597818 164426 598054
rect 164662 597818 164746 598054
rect 164982 597818 200426 598054
rect 200662 597818 200746 598054
rect 200982 597818 236426 598054
rect 236662 597818 236746 598054
rect 236982 597818 560426 598054
rect 560662 597818 560746 598054
rect 560982 597818 590142 598054
rect 590378 597818 590462 598054
rect 590698 597818 592650 598054
rect -8726 597734 592650 597818
rect -8726 597498 -6774 597734
rect -6538 597498 -6454 597734
rect -6218 597498 20426 597734
rect 20662 597498 20746 597734
rect 20982 597498 56426 597734
rect 56662 597498 56746 597734
rect 56982 597498 92426 597734
rect 92662 597498 92746 597734
rect 92982 597498 128426 597734
rect 128662 597498 128746 597734
rect 128982 597498 164426 597734
rect 164662 597498 164746 597734
rect 164982 597498 200426 597734
rect 200662 597498 200746 597734
rect 200982 597498 236426 597734
rect 236662 597498 236746 597734
rect 236982 597498 560426 597734
rect 560662 597498 560746 597734
rect 560982 597498 590142 597734
rect 590378 597498 590462 597734
rect 590698 597498 592650 597734
rect -8726 597466 592650 597498
rect -8726 594334 592650 594366
rect -8726 594098 -5814 594334
rect -5578 594098 -5494 594334
rect -5258 594098 16706 594334
rect 16942 594098 17026 594334
rect 17262 594098 52706 594334
rect 52942 594098 53026 594334
rect 53262 594098 124706 594334
rect 124942 594098 125026 594334
rect 125262 594098 160706 594334
rect 160942 594098 161026 594334
rect 161262 594098 196706 594334
rect 196942 594098 197026 594334
rect 197262 594098 232706 594334
rect 232942 594098 233026 594334
rect 233262 594098 556706 594334
rect 556942 594098 557026 594334
rect 557262 594098 589182 594334
rect 589418 594098 589502 594334
rect 589738 594098 592650 594334
rect -8726 594014 592650 594098
rect -8726 593778 -5814 594014
rect -5578 593778 -5494 594014
rect -5258 593778 16706 594014
rect 16942 593778 17026 594014
rect 17262 593778 52706 594014
rect 52942 593778 53026 594014
rect 53262 593778 124706 594014
rect 124942 593778 125026 594014
rect 125262 593778 160706 594014
rect 160942 593778 161026 594014
rect 161262 593778 196706 594014
rect 196942 593778 197026 594014
rect 197262 593778 232706 594014
rect 232942 593778 233026 594014
rect 233262 593778 556706 594014
rect 556942 593778 557026 594014
rect 557262 593778 589182 594014
rect 589418 593778 589502 594014
rect 589738 593778 592650 594014
rect -8726 593746 592650 593778
rect -8726 590614 592650 590646
rect -8726 590378 -4854 590614
rect -4618 590378 -4534 590614
rect -4298 590378 12986 590614
rect 13222 590378 13306 590614
rect 13542 590378 120986 590614
rect 121222 590378 121306 590614
rect 121542 590378 156986 590614
rect 157222 590378 157306 590614
rect 157542 590378 192986 590614
rect 193222 590378 193306 590614
rect 193542 590378 228986 590614
rect 229222 590378 229306 590614
rect 229542 590378 552986 590614
rect 553222 590378 553306 590614
rect 553542 590378 588222 590614
rect 588458 590378 588542 590614
rect 588778 590378 592650 590614
rect -8726 590294 592650 590378
rect -8726 590058 -4854 590294
rect -4618 590058 -4534 590294
rect -4298 590058 12986 590294
rect 13222 590058 13306 590294
rect 13542 590058 120986 590294
rect 121222 590058 121306 590294
rect 121542 590058 156986 590294
rect 157222 590058 157306 590294
rect 157542 590058 192986 590294
rect 193222 590058 193306 590294
rect 193542 590058 228986 590294
rect 229222 590058 229306 590294
rect 229542 590058 552986 590294
rect 553222 590058 553306 590294
rect 553542 590058 588222 590294
rect 588458 590058 588542 590294
rect 588778 590058 592650 590294
rect -8726 590026 592650 590058
rect -8726 586894 592650 586926
rect -8726 586658 -3894 586894
rect -3658 586658 -3574 586894
rect -3338 586658 9266 586894
rect 9502 586658 9586 586894
rect 9822 586658 45266 586894
rect 45502 586658 45586 586894
rect 45822 586658 117266 586894
rect 117502 586658 117586 586894
rect 117822 586658 153266 586894
rect 153502 586658 153586 586894
rect 153822 586658 189266 586894
rect 189502 586658 189586 586894
rect 189822 586658 225266 586894
rect 225502 586658 225586 586894
rect 225822 586658 587262 586894
rect 587498 586658 587582 586894
rect 587818 586658 592650 586894
rect -8726 586574 592650 586658
rect -8726 586338 -3894 586574
rect -3658 586338 -3574 586574
rect -3338 586338 9266 586574
rect 9502 586338 9586 586574
rect 9822 586338 45266 586574
rect 45502 586338 45586 586574
rect 45822 586338 117266 586574
rect 117502 586338 117586 586574
rect 117822 586338 153266 586574
rect 153502 586338 153586 586574
rect 153822 586338 189266 586574
rect 189502 586338 189586 586574
rect 189822 586338 225266 586574
rect 225502 586338 225586 586574
rect 225822 586338 587262 586574
rect 587498 586338 587582 586574
rect 587818 586338 592650 586574
rect -8726 586306 592650 586338
rect -8726 583174 592650 583206
rect -8726 582938 -2934 583174
rect -2698 582938 -2614 583174
rect -2378 582938 5546 583174
rect 5782 582938 5866 583174
rect 6102 582938 41546 583174
rect 41782 582938 41866 583174
rect 42102 582938 49610 583174
rect 49846 582938 80330 583174
rect 80566 582938 113546 583174
rect 113782 582938 113866 583174
rect 114102 582938 149546 583174
rect 149782 582938 149866 583174
rect 150102 582938 185546 583174
rect 185782 582938 185866 583174
rect 186102 582938 221546 583174
rect 221782 582938 221866 583174
rect 222102 582938 273210 583174
rect 273446 582938 303930 583174
rect 304166 582938 334650 583174
rect 334886 582938 365370 583174
rect 365606 582938 396090 583174
rect 396326 582938 426810 583174
rect 427046 582938 457530 583174
rect 457766 582938 488250 583174
rect 488486 582938 518970 583174
rect 519206 582938 545546 583174
rect 545782 582938 545866 583174
rect 546102 582938 549690 583174
rect 549926 582938 581546 583174
rect 581782 582938 581866 583174
rect 582102 582938 586302 583174
rect 586538 582938 586622 583174
rect 586858 582938 592650 583174
rect -8726 582854 592650 582938
rect -8726 582618 -2934 582854
rect -2698 582618 -2614 582854
rect -2378 582618 5546 582854
rect 5782 582618 5866 582854
rect 6102 582618 41546 582854
rect 41782 582618 41866 582854
rect 42102 582618 49610 582854
rect 49846 582618 80330 582854
rect 80566 582618 113546 582854
rect 113782 582618 113866 582854
rect 114102 582618 149546 582854
rect 149782 582618 149866 582854
rect 150102 582618 185546 582854
rect 185782 582618 185866 582854
rect 186102 582618 221546 582854
rect 221782 582618 221866 582854
rect 222102 582618 273210 582854
rect 273446 582618 303930 582854
rect 304166 582618 334650 582854
rect 334886 582618 365370 582854
rect 365606 582618 396090 582854
rect 396326 582618 426810 582854
rect 427046 582618 457530 582854
rect 457766 582618 488250 582854
rect 488486 582618 518970 582854
rect 519206 582618 545546 582854
rect 545782 582618 545866 582854
rect 546102 582618 549690 582854
rect 549926 582618 581546 582854
rect 581782 582618 581866 582854
rect 582102 582618 586302 582854
rect 586538 582618 586622 582854
rect 586858 582618 592650 582854
rect -8726 582586 592650 582618
rect -8726 579454 592650 579486
rect -8726 579218 -1974 579454
rect -1738 579218 -1654 579454
rect -1418 579218 1826 579454
rect 2062 579218 2146 579454
rect 2382 579218 34250 579454
rect 34486 579218 37826 579454
rect 38062 579218 38146 579454
rect 38382 579218 64970 579454
rect 65206 579218 95690 579454
rect 95926 579218 109826 579454
rect 110062 579218 110146 579454
rect 110382 579218 145826 579454
rect 146062 579218 146146 579454
rect 146382 579218 181826 579454
rect 182062 579218 182146 579454
rect 182382 579218 217826 579454
rect 218062 579218 218146 579454
rect 218382 579218 253826 579454
rect 254062 579218 254146 579454
rect 254382 579218 257850 579454
rect 258086 579218 288570 579454
rect 288806 579218 319290 579454
rect 319526 579218 350010 579454
rect 350246 579218 380730 579454
rect 380966 579218 411450 579454
rect 411686 579218 442170 579454
rect 442406 579218 472890 579454
rect 473126 579218 503610 579454
rect 503846 579218 534330 579454
rect 534566 579218 541826 579454
rect 542062 579218 542146 579454
rect 542382 579218 565050 579454
rect 565286 579218 577826 579454
rect 578062 579218 578146 579454
rect 578382 579218 585342 579454
rect 585578 579218 585662 579454
rect 585898 579218 592650 579454
rect -8726 579134 592650 579218
rect -8726 578898 -1974 579134
rect -1738 578898 -1654 579134
rect -1418 578898 1826 579134
rect 2062 578898 2146 579134
rect 2382 578898 34250 579134
rect 34486 578898 37826 579134
rect 38062 578898 38146 579134
rect 38382 578898 64970 579134
rect 65206 578898 95690 579134
rect 95926 578898 109826 579134
rect 110062 578898 110146 579134
rect 110382 578898 145826 579134
rect 146062 578898 146146 579134
rect 146382 578898 181826 579134
rect 182062 578898 182146 579134
rect 182382 578898 217826 579134
rect 218062 578898 218146 579134
rect 218382 578898 253826 579134
rect 254062 578898 254146 579134
rect 254382 578898 257850 579134
rect 258086 578898 288570 579134
rect 288806 578898 319290 579134
rect 319526 578898 350010 579134
rect 350246 578898 380730 579134
rect 380966 578898 411450 579134
rect 411686 578898 442170 579134
rect 442406 578898 472890 579134
rect 473126 578898 503610 579134
rect 503846 578898 534330 579134
rect 534566 578898 541826 579134
rect 542062 578898 542146 579134
rect 542382 578898 565050 579134
rect 565286 578898 577826 579134
rect 578062 578898 578146 579134
rect 578382 578898 585342 579134
rect 585578 578898 585662 579134
rect 585898 578898 592650 579134
rect -8726 578866 592650 578898
rect -8726 569494 592650 569526
rect -8726 569258 -8694 569494
rect -8458 569258 -8374 569494
rect -8138 569258 27866 569494
rect 28102 569258 28186 569494
rect 28422 569258 135866 569494
rect 136102 569258 136186 569494
rect 136422 569258 171866 569494
rect 172102 569258 172186 569494
rect 172422 569258 207866 569494
rect 208102 569258 208186 569494
rect 208422 569258 243866 569494
rect 244102 569258 244186 569494
rect 244422 569258 567866 569494
rect 568102 569258 568186 569494
rect 568422 569258 592062 569494
rect 592298 569258 592382 569494
rect 592618 569258 592650 569494
rect -8726 569174 592650 569258
rect -8726 568938 -8694 569174
rect -8458 568938 -8374 569174
rect -8138 568938 27866 569174
rect 28102 568938 28186 569174
rect 28422 568938 135866 569174
rect 136102 568938 136186 569174
rect 136422 568938 171866 569174
rect 172102 568938 172186 569174
rect 172422 568938 207866 569174
rect 208102 568938 208186 569174
rect 208422 568938 243866 569174
rect 244102 568938 244186 569174
rect 244422 568938 567866 569174
rect 568102 568938 568186 569174
rect 568422 568938 592062 569174
rect 592298 568938 592382 569174
rect 592618 568938 592650 569174
rect -8726 568906 592650 568938
rect -8726 565774 592650 565806
rect -8726 565538 -7734 565774
rect -7498 565538 -7414 565774
rect -7178 565538 24146 565774
rect 24382 565538 24466 565774
rect 24702 565538 60146 565774
rect 60382 565538 60466 565774
rect 60702 565538 132146 565774
rect 132382 565538 132466 565774
rect 132702 565538 168146 565774
rect 168382 565538 168466 565774
rect 168702 565538 204146 565774
rect 204382 565538 204466 565774
rect 204702 565538 240146 565774
rect 240382 565538 240466 565774
rect 240702 565538 564146 565774
rect 564382 565538 564466 565774
rect 564702 565538 591102 565774
rect 591338 565538 591422 565774
rect 591658 565538 592650 565774
rect -8726 565454 592650 565538
rect -8726 565218 -7734 565454
rect -7498 565218 -7414 565454
rect -7178 565218 24146 565454
rect 24382 565218 24466 565454
rect 24702 565218 60146 565454
rect 60382 565218 60466 565454
rect 60702 565218 132146 565454
rect 132382 565218 132466 565454
rect 132702 565218 168146 565454
rect 168382 565218 168466 565454
rect 168702 565218 204146 565454
rect 204382 565218 204466 565454
rect 204702 565218 240146 565454
rect 240382 565218 240466 565454
rect 240702 565218 564146 565454
rect 564382 565218 564466 565454
rect 564702 565218 591102 565454
rect 591338 565218 591422 565454
rect 591658 565218 592650 565454
rect -8726 565186 592650 565218
rect -8726 562054 592650 562086
rect -8726 561818 -6774 562054
rect -6538 561818 -6454 562054
rect -6218 561818 20426 562054
rect 20662 561818 20746 562054
rect 20982 561818 56426 562054
rect 56662 561818 56746 562054
rect 56982 561818 128426 562054
rect 128662 561818 128746 562054
rect 128982 561818 164426 562054
rect 164662 561818 164746 562054
rect 164982 561818 200426 562054
rect 200662 561818 200746 562054
rect 200982 561818 236426 562054
rect 236662 561818 236746 562054
rect 236982 561818 560426 562054
rect 560662 561818 560746 562054
rect 560982 561818 590142 562054
rect 590378 561818 590462 562054
rect 590698 561818 592650 562054
rect -8726 561734 592650 561818
rect -8726 561498 -6774 561734
rect -6538 561498 -6454 561734
rect -6218 561498 20426 561734
rect 20662 561498 20746 561734
rect 20982 561498 56426 561734
rect 56662 561498 56746 561734
rect 56982 561498 128426 561734
rect 128662 561498 128746 561734
rect 128982 561498 164426 561734
rect 164662 561498 164746 561734
rect 164982 561498 200426 561734
rect 200662 561498 200746 561734
rect 200982 561498 236426 561734
rect 236662 561498 236746 561734
rect 236982 561498 560426 561734
rect 560662 561498 560746 561734
rect 560982 561498 590142 561734
rect 590378 561498 590462 561734
rect 590698 561498 592650 561734
rect -8726 561466 592650 561498
rect -8726 558334 592650 558366
rect -8726 558098 -5814 558334
rect -5578 558098 -5494 558334
rect -5258 558098 16706 558334
rect 16942 558098 17026 558334
rect 17262 558098 52706 558334
rect 52942 558098 53026 558334
rect 53262 558098 124706 558334
rect 124942 558098 125026 558334
rect 125262 558098 160706 558334
rect 160942 558098 161026 558334
rect 161262 558098 196706 558334
rect 196942 558098 197026 558334
rect 197262 558098 232706 558334
rect 232942 558098 233026 558334
rect 233262 558098 556706 558334
rect 556942 558098 557026 558334
rect 557262 558098 589182 558334
rect 589418 558098 589502 558334
rect 589738 558098 592650 558334
rect -8726 558014 592650 558098
rect -8726 557778 -5814 558014
rect -5578 557778 -5494 558014
rect -5258 557778 16706 558014
rect 16942 557778 17026 558014
rect 17262 557778 52706 558014
rect 52942 557778 53026 558014
rect 53262 557778 124706 558014
rect 124942 557778 125026 558014
rect 125262 557778 160706 558014
rect 160942 557778 161026 558014
rect 161262 557778 196706 558014
rect 196942 557778 197026 558014
rect 197262 557778 232706 558014
rect 232942 557778 233026 558014
rect 233262 557778 556706 558014
rect 556942 557778 557026 558014
rect 557262 557778 589182 558014
rect 589418 557778 589502 558014
rect 589738 557778 592650 558014
rect -8726 557746 592650 557778
rect -8726 554614 592650 554646
rect -8726 554378 -4854 554614
rect -4618 554378 -4534 554614
rect -4298 554378 12986 554614
rect 13222 554378 13306 554614
rect 13542 554378 120986 554614
rect 121222 554378 121306 554614
rect 121542 554378 156986 554614
rect 157222 554378 157306 554614
rect 157542 554378 192986 554614
rect 193222 554378 193306 554614
rect 193542 554378 228986 554614
rect 229222 554378 229306 554614
rect 229542 554378 552986 554614
rect 553222 554378 553306 554614
rect 553542 554378 588222 554614
rect 588458 554378 588542 554614
rect 588778 554378 592650 554614
rect -8726 554294 592650 554378
rect -8726 554058 -4854 554294
rect -4618 554058 -4534 554294
rect -4298 554058 12986 554294
rect 13222 554058 13306 554294
rect 13542 554058 120986 554294
rect 121222 554058 121306 554294
rect 121542 554058 156986 554294
rect 157222 554058 157306 554294
rect 157542 554058 192986 554294
rect 193222 554058 193306 554294
rect 193542 554058 228986 554294
rect 229222 554058 229306 554294
rect 229542 554058 552986 554294
rect 553222 554058 553306 554294
rect 553542 554058 588222 554294
rect 588458 554058 588542 554294
rect 588778 554058 592650 554294
rect -8726 554026 592650 554058
rect -8726 550894 592650 550926
rect -8726 550658 -3894 550894
rect -3658 550658 -3574 550894
rect -3338 550658 9266 550894
rect 9502 550658 9586 550894
rect 9822 550658 45266 550894
rect 45502 550658 45586 550894
rect 45822 550658 117266 550894
rect 117502 550658 117586 550894
rect 117822 550658 153266 550894
rect 153502 550658 153586 550894
rect 153822 550658 189266 550894
rect 189502 550658 189586 550894
rect 189822 550658 225266 550894
rect 225502 550658 225586 550894
rect 225822 550658 587262 550894
rect 587498 550658 587582 550894
rect 587818 550658 592650 550894
rect -8726 550574 592650 550658
rect -8726 550338 -3894 550574
rect -3658 550338 -3574 550574
rect -3338 550338 9266 550574
rect 9502 550338 9586 550574
rect 9822 550338 45266 550574
rect 45502 550338 45586 550574
rect 45822 550338 117266 550574
rect 117502 550338 117586 550574
rect 117822 550338 153266 550574
rect 153502 550338 153586 550574
rect 153822 550338 189266 550574
rect 189502 550338 189586 550574
rect 189822 550338 225266 550574
rect 225502 550338 225586 550574
rect 225822 550338 587262 550574
rect 587498 550338 587582 550574
rect 587818 550338 592650 550574
rect -8726 550306 592650 550338
rect -8726 547174 592650 547206
rect -8726 546938 -2934 547174
rect -2698 546938 -2614 547174
rect -2378 546938 5546 547174
rect 5782 546938 5866 547174
rect 6102 546938 41546 547174
rect 41782 546938 41866 547174
rect 42102 546938 49610 547174
rect 49846 546938 80330 547174
rect 80566 546938 113546 547174
rect 113782 546938 113866 547174
rect 114102 546938 149546 547174
rect 149782 546938 149866 547174
rect 150102 546938 185546 547174
rect 185782 546938 185866 547174
rect 186102 546938 221546 547174
rect 221782 546938 221866 547174
rect 222102 546938 273210 547174
rect 273446 546938 303930 547174
rect 304166 546938 334650 547174
rect 334886 546938 365370 547174
rect 365606 546938 396090 547174
rect 396326 546938 426810 547174
rect 427046 546938 457530 547174
rect 457766 546938 488250 547174
rect 488486 546938 518970 547174
rect 519206 546938 545546 547174
rect 545782 546938 545866 547174
rect 546102 546938 549690 547174
rect 549926 546938 581546 547174
rect 581782 546938 581866 547174
rect 582102 546938 586302 547174
rect 586538 546938 586622 547174
rect 586858 546938 592650 547174
rect -8726 546854 592650 546938
rect -8726 546618 -2934 546854
rect -2698 546618 -2614 546854
rect -2378 546618 5546 546854
rect 5782 546618 5866 546854
rect 6102 546618 41546 546854
rect 41782 546618 41866 546854
rect 42102 546618 49610 546854
rect 49846 546618 80330 546854
rect 80566 546618 113546 546854
rect 113782 546618 113866 546854
rect 114102 546618 149546 546854
rect 149782 546618 149866 546854
rect 150102 546618 185546 546854
rect 185782 546618 185866 546854
rect 186102 546618 221546 546854
rect 221782 546618 221866 546854
rect 222102 546618 273210 546854
rect 273446 546618 303930 546854
rect 304166 546618 334650 546854
rect 334886 546618 365370 546854
rect 365606 546618 396090 546854
rect 396326 546618 426810 546854
rect 427046 546618 457530 546854
rect 457766 546618 488250 546854
rect 488486 546618 518970 546854
rect 519206 546618 545546 546854
rect 545782 546618 545866 546854
rect 546102 546618 549690 546854
rect 549926 546618 581546 546854
rect 581782 546618 581866 546854
rect 582102 546618 586302 546854
rect 586538 546618 586622 546854
rect 586858 546618 592650 546854
rect -8726 546586 592650 546618
rect -8726 543454 592650 543486
rect -8726 543218 -1974 543454
rect -1738 543218 -1654 543454
rect -1418 543218 1826 543454
rect 2062 543218 2146 543454
rect 2382 543218 34250 543454
rect 34486 543218 37826 543454
rect 38062 543218 38146 543454
rect 38382 543218 64970 543454
rect 65206 543218 95690 543454
rect 95926 543218 109826 543454
rect 110062 543218 110146 543454
rect 110382 543218 145826 543454
rect 146062 543218 146146 543454
rect 146382 543218 181826 543454
rect 182062 543218 182146 543454
rect 182382 543218 217826 543454
rect 218062 543218 218146 543454
rect 218382 543218 253826 543454
rect 254062 543218 254146 543454
rect 254382 543218 257850 543454
rect 258086 543218 288570 543454
rect 288806 543218 319290 543454
rect 319526 543218 350010 543454
rect 350246 543218 380730 543454
rect 380966 543218 411450 543454
rect 411686 543218 442170 543454
rect 442406 543218 472890 543454
rect 473126 543218 503610 543454
rect 503846 543218 534330 543454
rect 534566 543218 541826 543454
rect 542062 543218 542146 543454
rect 542382 543218 565050 543454
rect 565286 543218 577826 543454
rect 578062 543218 578146 543454
rect 578382 543218 585342 543454
rect 585578 543218 585662 543454
rect 585898 543218 592650 543454
rect -8726 543134 592650 543218
rect -8726 542898 -1974 543134
rect -1738 542898 -1654 543134
rect -1418 542898 1826 543134
rect 2062 542898 2146 543134
rect 2382 542898 34250 543134
rect 34486 542898 37826 543134
rect 38062 542898 38146 543134
rect 38382 542898 64970 543134
rect 65206 542898 95690 543134
rect 95926 542898 109826 543134
rect 110062 542898 110146 543134
rect 110382 542898 145826 543134
rect 146062 542898 146146 543134
rect 146382 542898 181826 543134
rect 182062 542898 182146 543134
rect 182382 542898 217826 543134
rect 218062 542898 218146 543134
rect 218382 542898 253826 543134
rect 254062 542898 254146 543134
rect 254382 542898 257850 543134
rect 258086 542898 288570 543134
rect 288806 542898 319290 543134
rect 319526 542898 350010 543134
rect 350246 542898 380730 543134
rect 380966 542898 411450 543134
rect 411686 542898 442170 543134
rect 442406 542898 472890 543134
rect 473126 542898 503610 543134
rect 503846 542898 534330 543134
rect 534566 542898 541826 543134
rect 542062 542898 542146 543134
rect 542382 542898 565050 543134
rect 565286 542898 577826 543134
rect 578062 542898 578146 543134
rect 578382 542898 585342 543134
rect 585578 542898 585662 543134
rect 585898 542898 592650 543134
rect -8726 542866 592650 542898
rect -8726 533494 592650 533526
rect -8726 533258 -8694 533494
rect -8458 533258 -8374 533494
rect -8138 533258 27866 533494
rect 28102 533258 28186 533494
rect 28422 533258 135866 533494
rect 136102 533258 136186 533494
rect 136422 533258 171866 533494
rect 172102 533258 172186 533494
rect 172422 533258 207866 533494
rect 208102 533258 208186 533494
rect 208422 533258 243866 533494
rect 244102 533258 244186 533494
rect 244422 533258 567866 533494
rect 568102 533258 568186 533494
rect 568422 533258 592062 533494
rect 592298 533258 592382 533494
rect 592618 533258 592650 533494
rect -8726 533174 592650 533258
rect -8726 532938 -8694 533174
rect -8458 532938 -8374 533174
rect -8138 532938 27866 533174
rect 28102 532938 28186 533174
rect 28422 532938 135866 533174
rect 136102 532938 136186 533174
rect 136422 532938 171866 533174
rect 172102 532938 172186 533174
rect 172422 532938 207866 533174
rect 208102 532938 208186 533174
rect 208422 532938 243866 533174
rect 244102 532938 244186 533174
rect 244422 532938 567866 533174
rect 568102 532938 568186 533174
rect 568422 532938 592062 533174
rect 592298 532938 592382 533174
rect 592618 532938 592650 533174
rect -8726 532906 592650 532938
rect -8726 529774 592650 529806
rect -8726 529538 -7734 529774
rect -7498 529538 -7414 529774
rect -7178 529538 24146 529774
rect 24382 529538 24466 529774
rect 24702 529538 60146 529774
rect 60382 529538 60466 529774
rect 60702 529538 132146 529774
rect 132382 529538 132466 529774
rect 132702 529538 168146 529774
rect 168382 529538 168466 529774
rect 168702 529538 204146 529774
rect 204382 529538 204466 529774
rect 204702 529538 240146 529774
rect 240382 529538 240466 529774
rect 240702 529538 276146 529774
rect 276382 529538 276466 529774
rect 276702 529538 312146 529774
rect 312382 529538 312466 529774
rect 312702 529538 348146 529774
rect 348382 529538 348466 529774
rect 348702 529538 384146 529774
rect 384382 529538 384466 529774
rect 384702 529538 420146 529774
rect 420382 529538 420466 529774
rect 420702 529538 456146 529774
rect 456382 529538 456466 529774
rect 456702 529538 492146 529774
rect 492382 529538 492466 529774
rect 492702 529538 528146 529774
rect 528382 529538 528466 529774
rect 528702 529538 564146 529774
rect 564382 529538 564466 529774
rect 564702 529538 591102 529774
rect 591338 529538 591422 529774
rect 591658 529538 592650 529774
rect -8726 529454 592650 529538
rect -8726 529218 -7734 529454
rect -7498 529218 -7414 529454
rect -7178 529218 24146 529454
rect 24382 529218 24466 529454
rect 24702 529218 60146 529454
rect 60382 529218 60466 529454
rect 60702 529218 132146 529454
rect 132382 529218 132466 529454
rect 132702 529218 168146 529454
rect 168382 529218 168466 529454
rect 168702 529218 204146 529454
rect 204382 529218 204466 529454
rect 204702 529218 240146 529454
rect 240382 529218 240466 529454
rect 240702 529218 276146 529454
rect 276382 529218 276466 529454
rect 276702 529218 312146 529454
rect 312382 529218 312466 529454
rect 312702 529218 348146 529454
rect 348382 529218 348466 529454
rect 348702 529218 384146 529454
rect 384382 529218 384466 529454
rect 384702 529218 420146 529454
rect 420382 529218 420466 529454
rect 420702 529218 456146 529454
rect 456382 529218 456466 529454
rect 456702 529218 492146 529454
rect 492382 529218 492466 529454
rect 492702 529218 528146 529454
rect 528382 529218 528466 529454
rect 528702 529218 564146 529454
rect 564382 529218 564466 529454
rect 564702 529218 591102 529454
rect 591338 529218 591422 529454
rect 591658 529218 592650 529454
rect -8726 529186 592650 529218
rect -8726 526054 592650 526086
rect -8726 525818 -6774 526054
rect -6538 525818 -6454 526054
rect -6218 525818 20426 526054
rect 20662 525818 20746 526054
rect 20982 525818 56426 526054
rect 56662 525818 56746 526054
rect 56982 525818 128426 526054
rect 128662 525818 128746 526054
rect 128982 525818 164426 526054
rect 164662 525818 164746 526054
rect 164982 525818 200426 526054
rect 200662 525818 200746 526054
rect 200982 525818 236426 526054
rect 236662 525818 236746 526054
rect 236982 525818 560426 526054
rect 560662 525818 560746 526054
rect 560982 525818 590142 526054
rect 590378 525818 590462 526054
rect 590698 525818 592650 526054
rect -8726 525734 592650 525818
rect -8726 525498 -6774 525734
rect -6538 525498 -6454 525734
rect -6218 525498 20426 525734
rect 20662 525498 20746 525734
rect 20982 525498 56426 525734
rect 56662 525498 56746 525734
rect 56982 525498 128426 525734
rect 128662 525498 128746 525734
rect 128982 525498 164426 525734
rect 164662 525498 164746 525734
rect 164982 525498 200426 525734
rect 200662 525498 200746 525734
rect 200982 525498 236426 525734
rect 236662 525498 236746 525734
rect 236982 525498 560426 525734
rect 560662 525498 560746 525734
rect 560982 525498 590142 525734
rect 590378 525498 590462 525734
rect 590698 525498 592650 525734
rect -8726 525466 592650 525498
rect -8726 522334 592650 522366
rect -8726 522098 -5814 522334
rect -5578 522098 -5494 522334
rect -5258 522098 16706 522334
rect 16942 522098 17026 522334
rect 17262 522098 52706 522334
rect 52942 522098 53026 522334
rect 53262 522098 124706 522334
rect 124942 522098 125026 522334
rect 125262 522098 160706 522334
rect 160942 522098 161026 522334
rect 161262 522098 196706 522334
rect 196942 522098 197026 522334
rect 197262 522098 232706 522334
rect 232942 522098 233026 522334
rect 233262 522098 556706 522334
rect 556942 522098 557026 522334
rect 557262 522098 589182 522334
rect 589418 522098 589502 522334
rect 589738 522098 592650 522334
rect -8726 522014 592650 522098
rect -8726 521778 -5814 522014
rect -5578 521778 -5494 522014
rect -5258 521778 16706 522014
rect 16942 521778 17026 522014
rect 17262 521778 52706 522014
rect 52942 521778 53026 522014
rect 53262 521778 124706 522014
rect 124942 521778 125026 522014
rect 125262 521778 160706 522014
rect 160942 521778 161026 522014
rect 161262 521778 196706 522014
rect 196942 521778 197026 522014
rect 197262 521778 232706 522014
rect 232942 521778 233026 522014
rect 233262 521778 556706 522014
rect 556942 521778 557026 522014
rect 557262 521778 589182 522014
rect 589418 521778 589502 522014
rect 589738 521778 592650 522014
rect -8726 521746 592650 521778
rect -8726 518614 592650 518646
rect -8726 518378 -4854 518614
rect -4618 518378 -4534 518614
rect -4298 518378 12986 518614
rect 13222 518378 13306 518614
rect 13542 518378 120986 518614
rect 121222 518378 121306 518614
rect 121542 518378 156986 518614
rect 157222 518378 157306 518614
rect 157542 518378 192986 518614
rect 193222 518378 193306 518614
rect 193542 518378 228986 518614
rect 229222 518378 229306 518614
rect 229542 518378 552986 518614
rect 553222 518378 553306 518614
rect 553542 518378 588222 518614
rect 588458 518378 588542 518614
rect 588778 518378 592650 518614
rect -8726 518294 592650 518378
rect -8726 518058 -4854 518294
rect -4618 518058 -4534 518294
rect -4298 518058 12986 518294
rect 13222 518058 13306 518294
rect 13542 518058 120986 518294
rect 121222 518058 121306 518294
rect 121542 518058 156986 518294
rect 157222 518058 157306 518294
rect 157542 518058 192986 518294
rect 193222 518058 193306 518294
rect 193542 518058 228986 518294
rect 229222 518058 229306 518294
rect 229542 518058 552986 518294
rect 553222 518058 553306 518294
rect 553542 518058 588222 518294
rect 588458 518058 588542 518294
rect 588778 518058 592650 518294
rect -8726 518026 592650 518058
rect -8726 514894 592650 514926
rect -8726 514658 -3894 514894
rect -3658 514658 -3574 514894
rect -3338 514658 9266 514894
rect 9502 514658 9586 514894
rect 9822 514658 45266 514894
rect 45502 514658 45586 514894
rect 45822 514658 117266 514894
rect 117502 514658 117586 514894
rect 117822 514658 153266 514894
rect 153502 514658 153586 514894
rect 153822 514658 189266 514894
rect 189502 514658 189586 514894
rect 189822 514658 225266 514894
rect 225502 514658 225586 514894
rect 225822 514658 587262 514894
rect 587498 514658 587582 514894
rect 587818 514658 592650 514894
rect -8726 514574 592650 514658
rect -8726 514338 -3894 514574
rect -3658 514338 -3574 514574
rect -3338 514338 9266 514574
rect 9502 514338 9586 514574
rect 9822 514338 45266 514574
rect 45502 514338 45586 514574
rect 45822 514338 117266 514574
rect 117502 514338 117586 514574
rect 117822 514338 153266 514574
rect 153502 514338 153586 514574
rect 153822 514338 189266 514574
rect 189502 514338 189586 514574
rect 189822 514338 225266 514574
rect 225502 514338 225586 514574
rect 225822 514338 587262 514574
rect 587498 514338 587582 514574
rect 587818 514338 592650 514574
rect -8726 514306 592650 514338
rect -8726 511174 592650 511206
rect -8726 510938 -2934 511174
rect -2698 510938 -2614 511174
rect -2378 510938 5546 511174
rect 5782 510938 5866 511174
rect 6102 510938 41546 511174
rect 41782 510938 41866 511174
rect 42102 510938 49610 511174
rect 49846 510938 80330 511174
rect 80566 510938 113546 511174
rect 113782 510938 113866 511174
rect 114102 510938 149546 511174
rect 149782 510938 149866 511174
rect 150102 510938 185546 511174
rect 185782 510938 185866 511174
rect 186102 510938 221546 511174
rect 221782 510938 221866 511174
rect 222102 510938 545546 511174
rect 545782 510938 545866 511174
rect 546102 510938 581546 511174
rect 581782 510938 581866 511174
rect 582102 510938 586302 511174
rect 586538 510938 586622 511174
rect 586858 510938 592650 511174
rect -8726 510854 592650 510938
rect -8726 510618 -2934 510854
rect -2698 510618 -2614 510854
rect -2378 510618 5546 510854
rect 5782 510618 5866 510854
rect 6102 510618 41546 510854
rect 41782 510618 41866 510854
rect 42102 510618 49610 510854
rect 49846 510618 80330 510854
rect 80566 510618 113546 510854
rect 113782 510618 113866 510854
rect 114102 510618 149546 510854
rect 149782 510618 149866 510854
rect 150102 510618 185546 510854
rect 185782 510618 185866 510854
rect 186102 510618 221546 510854
rect 221782 510618 221866 510854
rect 222102 510618 545546 510854
rect 545782 510618 545866 510854
rect 546102 510618 581546 510854
rect 581782 510618 581866 510854
rect 582102 510618 586302 510854
rect 586538 510618 586622 510854
rect 586858 510618 592650 510854
rect -8726 510586 592650 510618
rect -8726 507454 592650 507486
rect -8726 507218 -1974 507454
rect -1738 507218 -1654 507454
rect -1418 507218 1826 507454
rect 2062 507218 2146 507454
rect 2382 507218 34250 507454
rect 34486 507218 37826 507454
rect 38062 507218 38146 507454
rect 38382 507218 64970 507454
rect 65206 507218 95690 507454
rect 95926 507218 109826 507454
rect 110062 507218 110146 507454
rect 110382 507218 145826 507454
rect 146062 507218 146146 507454
rect 146382 507218 181826 507454
rect 182062 507218 182146 507454
rect 182382 507218 217826 507454
rect 218062 507218 218146 507454
rect 218382 507218 253826 507454
rect 254062 507218 254146 507454
rect 254382 507218 541826 507454
rect 542062 507218 542146 507454
rect 542382 507218 577826 507454
rect 578062 507218 578146 507454
rect 578382 507218 585342 507454
rect 585578 507218 585662 507454
rect 585898 507218 592650 507454
rect -8726 507134 592650 507218
rect -8726 506898 -1974 507134
rect -1738 506898 -1654 507134
rect -1418 506898 1826 507134
rect 2062 506898 2146 507134
rect 2382 506898 34250 507134
rect 34486 506898 37826 507134
rect 38062 506898 38146 507134
rect 38382 506898 64970 507134
rect 65206 506898 95690 507134
rect 95926 506898 109826 507134
rect 110062 506898 110146 507134
rect 110382 506898 145826 507134
rect 146062 506898 146146 507134
rect 146382 506898 181826 507134
rect 182062 506898 182146 507134
rect 182382 506898 217826 507134
rect 218062 506898 218146 507134
rect 218382 506898 253826 507134
rect 254062 506898 254146 507134
rect 254382 506898 541826 507134
rect 542062 506898 542146 507134
rect 542382 506898 577826 507134
rect 578062 506898 578146 507134
rect 578382 506898 585342 507134
rect 585578 506898 585662 507134
rect 585898 506898 592650 507134
rect -8726 506866 592650 506898
rect -8726 497494 592650 497526
rect -8726 497258 -8694 497494
rect -8458 497258 -8374 497494
rect -8138 497258 27866 497494
rect 28102 497258 28186 497494
rect 28422 497258 135866 497494
rect 136102 497258 136186 497494
rect 136422 497258 171866 497494
rect 172102 497258 172186 497494
rect 172422 497258 207866 497494
rect 208102 497258 208186 497494
rect 208422 497258 243866 497494
rect 244102 497258 244186 497494
rect 244422 497258 567866 497494
rect 568102 497258 568186 497494
rect 568422 497258 592062 497494
rect 592298 497258 592382 497494
rect 592618 497258 592650 497494
rect -8726 497174 592650 497258
rect -8726 496938 -8694 497174
rect -8458 496938 -8374 497174
rect -8138 496938 27866 497174
rect 28102 496938 28186 497174
rect 28422 496938 135866 497174
rect 136102 496938 136186 497174
rect 136422 496938 171866 497174
rect 172102 496938 172186 497174
rect 172422 496938 207866 497174
rect 208102 496938 208186 497174
rect 208422 496938 243866 497174
rect 244102 496938 244186 497174
rect 244422 496938 567866 497174
rect 568102 496938 568186 497174
rect 568422 496938 592062 497174
rect 592298 496938 592382 497174
rect 592618 496938 592650 497174
rect -8726 496906 592650 496938
rect -8726 493774 592650 493806
rect -8726 493538 -7734 493774
rect -7498 493538 -7414 493774
rect -7178 493538 24146 493774
rect 24382 493538 24466 493774
rect 24702 493538 60146 493774
rect 60382 493538 60466 493774
rect 60702 493538 132146 493774
rect 132382 493538 132466 493774
rect 132702 493538 168146 493774
rect 168382 493538 168466 493774
rect 168702 493538 204146 493774
rect 204382 493538 204466 493774
rect 204702 493538 240146 493774
rect 240382 493538 240466 493774
rect 240702 493538 564146 493774
rect 564382 493538 564466 493774
rect 564702 493538 591102 493774
rect 591338 493538 591422 493774
rect 591658 493538 592650 493774
rect -8726 493454 592650 493538
rect -8726 493218 -7734 493454
rect -7498 493218 -7414 493454
rect -7178 493218 24146 493454
rect 24382 493218 24466 493454
rect 24702 493218 60146 493454
rect 60382 493218 60466 493454
rect 60702 493218 132146 493454
rect 132382 493218 132466 493454
rect 132702 493218 168146 493454
rect 168382 493218 168466 493454
rect 168702 493218 204146 493454
rect 204382 493218 204466 493454
rect 204702 493218 240146 493454
rect 240382 493218 240466 493454
rect 240702 493218 564146 493454
rect 564382 493218 564466 493454
rect 564702 493218 591102 493454
rect 591338 493218 591422 493454
rect 591658 493218 592650 493454
rect -8726 493186 592650 493218
rect -8726 490054 592650 490086
rect -8726 489818 -6774 490054
rect -6538 489818 -6454 490054
rect -6218 489818 20426 490054
rect 20662 489818 20746 490054
rect 20982 489818 56426 490054
rect 56662 489818 56746 490054
rect 56982 489818 128426 490054
rect 128662 489818 128746 490054
rect 128982 489818 164426 490054
rect 164662 489818 164746 490054
rect 164982 489818 200426 490054
rect 200662 489818 200746 490054
rect 200982 489818 236426 490054
rect 236662 489818 236746 490054
rect 236982 489818 560426 490054
rect 560662 489818 560746 490054
rect 560982 489818 590142 490054
rect 590378 489818 590462 490054
rect 590698 489818 592650 490054
rect -8726 489734 592650 489818
rect -8726 489498 -6774 489734
rect -6538 489498 -6454 489734
rect -6218 489498 20426 489734
rect 20662 489498 20746 489734
rect 20982 489498 56426 489734
rect 56662 489498 56746 489734
rect 56982 489498 128426 489734
rect 128662 489498 128746 489734
rect 128982 489498 164426 489734
rect 164662 489498 164746 489734
rect 164982 489498 200426 489734
rect 200662 489498 200746 489734
rect 200982 489498 236426 489734
rect 236662 489498 236746 489734
rect 236982 489498 560426 489734
rect 560662 489498 560746 489734
rect 560982 489498 590142 489734
rect 590378 489498 590462 489734
rect 590698 489498 592650 489734
rect -8726 489466 592650 489498
rect -8726 486334 592650 486366
rect -8726 486098 -5814 486334
rect -5578 486098 -5494 486334
rect -5258 486098 16706 486334
rect 16942 486098 17026 486334
rect 17262 486098 52706 486334
rect 52942 486098 53026 486334
rect 53262 486098 124706 486334
rect 124942 486098 125026 486334
rect 125262 486098 160706 486334
rect 160942 486098 161026 486334
rect 161262 486098 196706 486334
rect 196942 486098 197026 486334
rect 197262 486098 232706 486334
rect 232942 486098 233026 486334
rect 233262 486098 556706 486334
rect 556942 486098 557026 486334
rect 557262 486098 589182 486334
rect 589418 486098 589502 486334
rect 589738 486098 592650 486334
rect -8726 486014 592650 486098
rect -8726 485778 -5814 486014
rect -5578 485778 -5494 486014
rect -5258 485778 16706 486014
rect 16942 485778 17026 486014
rect 17262 485778 52706 486014
rect 52942 485778 53026 486014
rect 53262 485778 124706 486014
rect 124942 485778 125026 486014
rect 125262 485778 160706 486014
rect 160942 485778 161026 486014
rect 161262 485778 196706 486014
rect 196942 485778 197026 486014
rect 197262 485778 232706 486014
rect 232942 485778 233026 486014
rect 233262 485778 556706 486014
rect 556942 485778 557026 486014
rect 557262 485778 589182 486014
rect 589418 485778 589502 486014
rect 589738 485778 592650 486014
rect -8726 485746 592650 485778
rect -8726 482614 592650 482646
rect -8726 482378 -4854 482614
rect -4618 482378 -4534 482614
rect -4298 482378 12986 482614
rect 13222 482378 13306 482614
rect 13542 482378 120986 482614
rect 121222 482378 121306 482614
rect 121542 482378 156986 482614
rect 157222 482378 157306 482614
rect 157542 482378 192986 482614
rect 193222 482378 193306 482614
rect 193542 482378 228986 482614
rect 229222 482378 229306 482614
rect 229542 482378 552986 482614
rect 553222 482378 553306 482614
rect 553542 482378 588222 482614
rect 588458 482378 588542 482614
rect 588778 482378 592650 482614
rect -8726 482294 592650 482378
rect -8726 482058 -4854 482294
rect -4618 482058 -4534 482294
rect -4298 482058 12986 482294
rect 13222 482058 13306 482294
rect 13542 482058 120986 482294
rect 121222 482058 121306 482294
rect 121542 482058 156986 482294
rect 157222 482058 157306 482294
rect 157542 482058 192986 482294
rect 193222 482058 193306 482294
rect 193542 482058 228986 482294
rect 229222 482058 229306 482294
rect 229542 482058 552986 482294
rect 553222 482058 553306 482294
rect 553542 482058 588222 482294
rect 588458 482058 588542 482294
rect 588778 482058 592650 482294
rect -8726 482026 592650 482058
rect -8726 478894 592650 478926
rect -8726 478658 -3894 478894
rect -3658 478658 -3574 478894
rect -3338 478658 9266 478894
rect 9502 478658 9586 478894
rect 9822 478658 45266 478894
rect 45502 478658 45586 478894
rect 45822 478658 117266 478894
rect 117502 478658 117586 478894
rect 117822 478658 153266 478894
rect 153502 478658 153586 478894
rect 153822 478658 189266 478894
rect 189502 478658 189586 478894
rect 189822 478658 225266 478894
rect 225502 478658 225586 478894
rect 225822 478658 587262 478894
rect 587498 478658 587582 478894
rect 587818 478658 592650 478894
rect -8726 478574 592650 478658
rect -8726 478338 -3894 478574
rect -3658 478338 -3574 478574
rect -3338 478338 9266 478574
rect 9502 478338 9586 478574
rect 9822 478338 45266 478574
rect 45502 478338 45586 478574
rect 45822 478338 117266 478574
rect 117502 478338 117586 478574
rect 117822 478338 153266 478574
rect 153502 478338 153586 478574
rect 153822 478338 189266 478574
rect 189502 478338 189586 478574
rect 189822 478338 225266 478574
rect 225502 478338 225586 478574
rect 225822 478338 587262 478574
rect 587498 478338 587582 478574
rect 587818 478338 592650 478574
rect -8726 478306 592650 478338
rect -8726 475174 592650 475206
rect -8726 474938 -2934 475174
rect -2698 474938 -2614 475174
rect -2378 474938 5546 475174
rect 5782 474938 5866 475174
rect 6102 474938 41546 475174
rect 41782 474938 41866 475174
rect 42102 474938 49610 475174
rect 49846 474938 80330 475174
rect 80566 474938 113546 475174
rect 113782 474938 113866 475174
rect 114102 474938 149546 475174
rect 149782 474938 149866 475174
rect 150102 474938 185546 475174
rect 185782 474938 185866 475174
rect 186102 474938 221546 475174
rect 221782 474938 221866 475174
rect 222102 474938 273210 475174
rect 273446 474938 303930 475174
rect 304166 474938 334650 475174
rect 334886 474938 365370 475174
rect 365606 474938 396090 475174
rect 396326 474938 426810 475174
rect 427046 474938 457530 475174
rect 457766 474938 488250 475174
rect 488486 474938 518970 475174
rect 519206 474938 545546 475174
rect 545782 474938 545866 475174
rect 546102 474938 549690 475174
rect 549926 474938 581546 475174
rect 581782 474938 581866 475174
rect 582102 474938 586302 475174
rect 586538 474938 586622 475174
rect 586858 474938 592650 475174
rect -8726 474854 592650 474938
rect -8726 474618 -2934 474854
rect -2698 474618 -2614 474854
rect -2378 474618 5546 474854
rect 5782 474618 5866 474854
rect 6102 474618 41546 474854
rect 41782 474618 41866 474854
rect 42102 474618 49610 474854
rect 49846 474618 80330 474854
rect 80566 474618 113546 474854
rect 113782 474618 113866 474854
rect 114102 474618 149546 474854
rect 149782 474618 149866 474854
rect 150102 474618 185546 474854
rect 185782 474618 185866 474854
rect 186102 474618 221546 474854
rect 221782 474618 221866 474854
rect 222102 474618 273210 474854
rect 273446 474618 303930 474854
rect 304166 474618 334650 474854
rect 334886 474618 365370 474854
rect 365606 474618 396090 474854
rect 396326 474618 426810 474854
rect 427046 474618 457530 474854
rect 457766 474618 488250 474854
rect 488486 474618 518970 474854
rect 519206 474618 545546 474854
rect 545782 474618 545866 474854
rect 546102 474618 549690 474854
rect 549926 474618 581546 474854
rect 581782 474618 581866 474854
rect 582102 474618 586302 474854
rect 586538 474618 586622 474854
rect 586858 474618 592650 474854
rect -8726 474586 592650 474618
rect -8726 471454 592650 471486
rect -8726 471218 -1974 471454
rect -1738 471218 -1654 471454
rect -1418 471218 1826 471454
rect 2062 471218 2146 471454
rect 2382 471218 34250 471454
rect 34486 471218 37826 471454
rect 38062 471218 38146 471454
rect 38382 471218 64970 471454
rect 65206 471218 95690 471454
rect 95926 471218 109826 471454
rect 110062 471218 110146 471454
rect 110382 471218 145826 471454
rect 146062 471218 146146 471454
rect 146382 471218 181826 471454
rect 182062 471218 182146 471454
rect 182382 471218 217826 471454
rect 218062 471218 218146 471454
rect 218382 471218 253826 471454
rect 254062 471218 254146 471454
rect 254382 471218 257850 471454
rect 258086 471218 288570 471454
rect 288806 471218 319290 471454
rect 319526 471218 350010 471454
rect 350246 471218 380730 471454
rect 380966 471218 411450 471454
rect 411686 471218 442170 471454
rect 442406 471218 472890 471454
rect 473126 471218 503610 471454
rect 503846 471218 534330 471454
rect 534566 471218 541826 471454
rect 542062 471218 542146 471454
rect 542382 471218 565050 471454
rect 565286 471218 577826 471454
rect 578062 471218 578146 471454
rect 578382 471218 585342 471454
rect 585578 471218 585662 471454
rect 585898 471218 592650 471454
rect -8726 471134 592650 471218
rect -8726 470898 -1974 471134
rect -1738 470898 -1654 471134
rect -1418 470898 1826 471134
rect 2062 470898 2146 471134
rect 2382 470898 34250 471134
rect 34486 470898 37826 471134
rect 38062 470898 38146 471134
rect 38382 470898 64970 471134
rect 65206 470898 95690 471134
rect 95926 470898 109826 471134
rect 110062 470898 110146 471134
rect 110382 470898 145826 471134
rect 146062 470898 146146 471134
rect 146382 470898 181826 471134
rect 182062 470898 182146 471134
rect 182382 470898 217826 471134
rect 218062 470898 218146 471134
rect 218382 470898 253826 471134
rect 254062 470898 254146 471134
rect 254382 470898 257850 471134
rect 258086 470898 288570 471134
rect 288806 470898 319290 471134
rect 319526 470898 350010 471134
rect 350246 470898 380730 471134
rect 380966 470898 411450 471134
rect 411686 470898 442170 471134
rect 442406 470898 472890 471134
rect 473126 470898 503610 471134
rect 503846 470898 534330 471134
rect 534566 470898 541826 471134
rect 542062 470898 542146 471134
rect 542382 470898 565050 471134
rect 565286 470898 577826 471134
rect 578062 470898 578146 471134
rect 578382 470898 585342 471134
rect 585578 470898 585662 471134
rect 585898 470898 592650 471134
rect -8726 470866 592650 470898
rect -8726 461494 592650 461526
rect -8726 461258 -8694 461494
rect -8458 461258 -8374 461494
rect -8138 461258 27866 461494
rect 28102 461258 28186 461494
rect 28422 461258 135866 461494
rect 136102 461258 136186 461494
rect 136422 461258 171866 461494
rect 172102 461258 172186 461494
rect 172422 461258 207866 461494
rect 208102 461258 208186 461494
rect 208422 461258 243866 461494
rect 244102 461258 244186 461494
rect 244422 461258 567866 461494
rect 568102 461258 568186 461494
rect 568422 461258 592062 461494
rect 592298 461258 592382 461494
rect 592618 461258 592650 461494
rect -8726 461174 592650 461258
rect -8726 460938 -8694 461174
rect -8458 460938 -8374 461174
rect -8138 460938 27866 461174
rect 28102 460938 28186 461174
rect 28422 460938 135866 461174
rect 136102 460938 136186 461174
rect 136422 460938 171866 461174
rect 172102 460938 172186 461174
rect 172422 460938 207866 461174
rect 208102 460938 208186 461174
rect 208422 460938 243866 461174
rect 244102 460938 244186 461174
rect 244422 460938 567866 461174
rect 568102 460938 568186 461174
rect 568422 460938 592062 461174
rect 592298 460938 592382 461174
rect 592618 460938 592650 461174
rect -8726 460906 592650 460938
rect -8726 457774 592650 457806
rect -8726 457538 -7734 457774
rect -7498 457538 -7414 457774
rect -7178 457538 24146 457774
rect 24382 457538 24466 457774
rect 24702 457538 60146 457774
rect 60382 457538 60466 457774
rect 60702 457538 132146 457774
rect 132382 457538 132466 457774
rect 132702 457538 168146 457774
rect 168382 457538 168466 457774
rect 168702 457538 204146 457774
rect 204382 457538 204466 457774
rect 204702 457538 240146 457774
rect 240382 457538 240466 457774
rect 240702 457538 564146 457774
rect 564382 457538 564466 457774
rect 564702 457538 591102 457774
rect 591338 457538 591422 457774
rect 591658 457538 592650 457774
rect -8726 457454 592650 457538
rect -8726 457218 -7734 457454
rect -7498 457218 -7414 457454
rect -7178 457218 24146 457454
rect 24382 457218 24466 457454
rect 24702 457218 60146 457454
rect 60382 457218 60466 457454
rect 60702 457218 132146 457454
rect 132382 457218 132466 457454
rect 132702 457218 168146 457454
rect 168382 457218 168466 457454
rect 168702 457218 204146 457454
rect 204382 457218 204466 457454
rect 204702 457218 240146 457454
rect 240382 457218 240466 457454
rect 240702 457218 564146 457454
rect 564382 457218 564466 457454
rect 564702 457218 591102 457454
rect 591338 457218 591422 457454
rect 591658 457218 592650 457454
rect -8726 457186 592650 457218
rect -8726 454054 592650 454086
rect -8726 453818 -6774 454054
rect -6538 453818 -6454 454054
rect -6218 453818 20426 454054
rect 20662 453818 20746 454054
rect 20982 453818 56426 454054
rect 56662 453818 56746 454054
rect 56982 453818 128426 454054
rect 128662 453818 128746 454054
rect 128982 453818 164426 454054
rect 164662 453818 164746 454054
rect 164982 453818 200426 454054
rect 200662 453818 200746 454054
rect 200982 453818 236426 454054
rect 236662 453818 236746 454054
rect 236982 453818 560426 454054
rect 560662 453818 560746 454054
rect 560982 453818 590142 454054
rect 590378 453818 590462 454054
rect 590698 453818 592650 454054
rect -8726 453734 592650 453818
rect -8726 453498 -6774 453734
rect -6538 453498 -6454 453734
rect -6218 453498 20426 453734
rect 20662 453498 20746 453734
rect 20982 453498 56426 453734
rect 56662 453498 56746 453734
rect 56982 453498 128426 453734
rect 128662 453498 128746 453734
rect 128982 453498 164426 453734
rect 164662 453498 164746 453734
rect 164982 453498 200426 453734
rect 200662 453498 200746 453734
rect 200982 453498 236426 453734
rect 236662 453498 236746 453734
rect 236982 453498 560426 453734
rect 560662 453498 560746 453734
rect 560982 453498 590142 453734
rect 590378 453498 590462 453734
rect 590698 453498 592650 453734
rect -8726 453466 592650 453498
rect -8726 450334 592650 450366
rect -8726 450098 -5814 450334
rect -5578 450098 -5494 450334
rect -5258 450098 16706 450334
rect 16942 450098 17026 450334
rect 17262 450098 52706 450334
rect 52942 450098 53026 450334
rect 53262 450098 124706 450334
rect 124942 450098 125026 450334
rect 125262 450098 160706 450334
rect 160942 450098 161026 450334
rect 161262 450098 196706 450334
rect 196942 450098 197026 450334
rect 197262 450098 232706 450334
rect 232942 450098 233026 450334
rect 233262 450098 556706 450334
rect 556942 450098 557026 450334
rect 557262 450098 589182 450334
rect 589418 450098 589502 450334
rect 589738 450098 592650 450334
rect -8726 450014 592650 450098
rect -8726 449778 -5814 450014
rect -5578 449778 -5494 450014
rect -5258 449778 16706 450014
rect 16942 449778 17026 450014
rect 17262 449778 52706 450014
rect 52942 449778 53026 450014
rect 53262 449778 124706 450014
rect 124942 449778 125026 450014
rect 125262 449778 160706 450014
rect 160942 449778 161026 450014
rect 161262 449778 196706 450014
rect 196942 449778 197026 450014
rect 197262 449778 232706 450014
rect 232942 449778 233026 450014
rect 233262 449778 556706 450014
rect 556942 449778 557026 450014
rect 557262 449778 589182 450014
rect 589418 449778 589502 450014
rect 589738 449778 592650 450014
rect -8726 449746 592650 449778
rect -8726 446614 592650 446646
rect -8726 446378 -4854 446614
rect -4618 446378 -4534 446614
rect -4298 446378 12986 446614
rect 13222 446378 13306 446614
rect 13542 446378 84986 446614
rect 85222 446378 85306 446614
rect 85542 446378 120986 446614
rect 121222 446378 121306 446614
rect 121542 446378 156986 446614
rect 157222 446378 157306 446614
rect 157542 446378 192986 446614
rect 193222 446378 193306 446614
rect 193542 446378 228986 446614
rect 229222 446378 229306 446614
rect 229542 446378 552986 446614
rect 553222 446378 553306 446614
rect 553542 446378 588222 446614
rect 588458 446378 588542 446614
rect 588778 446378 592650 446614
rect -8726 446294 592650 446378
rect -8726 446058 -4854 446294
rect -4618 446058 -4534 446294
rect -4298 446058 12986 446294
rect 13222 446058 13306 446294
rect 13542 446058 84986 446294
rect 85222 446058 85306 446294
rect 85542 446058 120986 446294
rect 121222 446058 121306 446294
rect 121542 446058 156986 446294
rect 157222 446058 157306 446294
rect 157542 446058 192986 446294
rect 193222 446058 193306 446294
rect 193542 446058 228986 446294
rect 229222 446058 229306 446294
rect 229542 446058 552986 446294
rect 553222 446058 553306 446294
rect 553542 446058 588222 446294
rect 588458 446058 588542 446294
rect 588778 446058 592650 446294
rect -8726 446026 592650 446058
rect -8726 442894 592650 442926
rect -8726 442658 -3894 442894
rect -3658 442658 -3574 442894
rect -3338 442658 9266 442894
rect 9502 442658 9586 442894
rect 9822 442658 45266 442894
rect 45502 442658 45586 442894
rect 45822 442658 81266 442894
rect 81502 442658 81586 442894
rect 81822 442658 117266 442894
rect 117502 442658 117586 442894
rect 117822 442658 153266 442894
rect 153502 442658 153586 442894
rect 153822 442658 189266 442894
rect 189502 442658 189586 442894
rect 189822 442658 225266 442894
rect 225502 442658 225586 442894
rect 225822 442658 587262 442894
rect 587498 442658 587582 442894
rect 587818 442658 592650 442894
rect -8726 442574 592650 442658
rect -8726 442338 -3894 442574
rect -3658 442338 -3574 442574
rect -3338 442338 9266 442574
rect 9502 442338 9586 442574
rect 9822 442338 45266 442574
rect 45502 442338 45586 442574
rect 45822 442338 81266 442574
rect 81502 442338 81586 442574
rect 81822 442338 117266 442574
rect 117502 442338 117586 442574
rect 117822 442338 153266 442574
rect 153502 442338 153586 442574
rect 153822 442338 189266 442574
rect 189502 442338 189586 442574
rect 189822 442338 225266 442574
rect 225502 442338 225586 442574
rect 225822 442338 587262 442574
rect 587498 442338 587582 442574
rect 587818 442338 592650 442574
rect -8726 442306 592650 442338
rect -8726 439174 592650 439206
rect -8726 438938 -2934 439174
rect -2698 438938 -2614 439174
rect -2378 438938 5546 439174
rect 5782 438938 5866 439174
rect 6102 438938 41546 439174
rect 41782 438938 41866 439174
rect 42102 438938 77546 439174
rect 77782 438938 77866 439174
rect 78102 438938 113546 439174
rect 113782 438938 113866 439174
rect 114102 438938 149546 439174
rect 149782 438938 149866 439174
rect 150102 438938 185546 439174
rect 185782 438938 185866 439174
rect 186102 438938 221546 439174
rect 221782 438938 221866 439174
rect 222102 438938 273210 439174
rect 273446 438938 303930 439174
rect 304166 438938 334650 439174
rect 334886 438938 365370 439174
rect 365606 438938 396090 439174
rect 396326 438938 426810 439174
rect 427046 438938 457530 439174
rect 457766 438938 488250 439174
rect 488486 438938 518970 439174
rect 519206 438938 545546 439174
rect 545782 438938 545866 439174
rect 546102 438938 549690 439174
rect 549926 438938 581546 439174
rect 581782 438938 581866 439174
rect 582102 438938 586302 439174
rect 586538 438938 586622 439174
rect 586858 438938 592650 439174
rect -8726 438854 592650 438938
rect -8726 438618 -2934 438854
rect -2698 438618 -2614 438854
rect -2378 438618 5546 438854
rect 5782 438618 5866 438854
rect 6102 438618 41546 438854
rect 41782 438618 41866 438854
rect 42102 438618 77546 438854
rect 77782 438618 77866 438854
rect 78102 438618 113546 438854
rect 113782 438618 113866 438854
rect 114102 438618 149546 438854
rect 149782 438618 149866 438854
rect 150102 438618 185546 438854
rect 185782 438618 185866 438854
rect 186102 438618 221546 438854
rect 221782 438618 221866 438854
rect 222102 438618 273210 438854
rect 273446 438618 303930 438854
rect 304166 438618 334650 438854
rect 334886 438618 365370 438854
rect 365606 438618 396090 438854
rect 396326 438618 426810 438854
rect 427046 438618 457530 438854
rect 457766 438618 488250 438854
rect 488486 438618 518970 438854
rect 519206 438618 545546 438854
rect 545782 438618 545866 438854
rect 546102 438618 549690 438854
rect 549926 438618 581546 438854
rect 581782 438618 581866 438854
rect 582102 438618 586302 438854
rect 586538 438618 586622 438854
rect 586858 438618 592650 438854
rect -8726 438586 592650 438618
rect -8726 435454 592650 435486
rect -8726 435218 -1974 435454
rect -1738 435218 -1654 435454
rect -1418 435218 1826 435454
rect 2062 435218 2146 435454
rect 2382 435218 37826 435454
rect 38062 435218 38146 435454
rect 38382 435218 73826 435454
rect 74062 435218 74146 435454
rect 74382 435218 109826 435454
rect 110062 435218 110146 435454
rect 110382 435218 145826 435454
rect 146062 435218 146146 435454
rect 146382 435218 181826 435454
rect 182062 435218 182146 435454
rect 182382 435218 217826 435454
rect 218062 435218 218146 435454
rect 218382 435218 253826 435454
rect 254062 435218 254146 435454
rect 254382 435218 257850 435454
rect 258086 435218 288570 435454
rect 288806 435218 319290 435454
rect 319526 435218 350010 435454
rect 350246 435218 380730 435454
rect 380966 435218 411450 435454
rect 411686 435218 442170 435454
rect 442406 435218 472890 435454
rect 473126 435218 503610 435454
rect 503846 435218 534330 435454
rect 534566 435218 541826 435454
rect 542062 435218 542146 435454
rect 542382 435218 565050 435454
rect 565286 435218 577826 435454
rect 578062 435218 578146 435454
rect 578382 435218 585342 435454
rect 585578 435218 585662 435454
rect 585898 435218 592650 435454
rect -8726 435134 592650 435218
rect -8726 434898 -1974 435134
rect -1738 434898 -1654 435134
rect -1418 434898 1826 435134
rect 2062 434898 2146 435134
rect 2382 434898 37826 435134
rect 38062 434898 38146 435134
rect 38382 434898 73826 435134
rect 74062 434898 74146 435134
rect 74382 434898 109826 435134
rect 110062 434898 110146 435134
rect 110382 434898 145826 435134
rect 146062 434898 146146 435134
rect 146382 434898 181826 435134
rect 182062 434898 182146 435134
rect 182382 434898 217826 435134
rect 218062 434898 218146 435134
rect 218382 434898 253826 435134
rect 254062 434898 254146 435134
rect 254382 434898 257850 435134
rect 258086 434898 288570 435134
rect 288806 434898 319290 435134
rect 319526 434898 350010 435134
rect 350246 434898 380730 435134
rect 380966 434898 411450 435134
rect 411686 434898 442170 435134
rect 442406 434898 472890 435134
rect 473126 434898 503610 435134
rect 503846 434898 534330 435134
rect 534566 434898 541826 435134
rect 542062 434898 542146 435134
rect 542382 434898 565050 435134
rect 565286 434898 577826 435134
rect 578062 434898 578146 435134
rect 578382 434898 585342 435134
rect 585578 434898 585662 435134
rect 585898 434898 592650 435134
rect -8726 434866 592650 434898
rect -8726 425494 592650 425526
rect -8726 425258 -8694 425494
rect -8458 425258 -8374 425494
rect -8138 425258 27866 425494
rect 28102 425258 28186 425494
rect 28422 425258 63866 425494
rect 64102 425258 64186 425494
rect 64422 425258 99866 425494
rect 100102 425258 100186 425494
rect 100422 425258 135866 425494
rect 136102 425258 136186 425494
rect 136422 425258 171866 425494
rect 172102 425258 172186 425494
rect 172422 425258 243866 425494
rect 244102 425258 244186 425494
rect 244422 425258 567866 425494
rect 568102 425258 568186 425494
rect 568422 425258 592062 425494
rect 592298 425258 592382 425494
rect 592618 425258 592650 425494
rect -8726 425174 592650 425258
rect -8726 424938 -8694 425174
rect -8458 424938 -8374 425174
rect -8138 424938 27866 425174
rect 28102 424938 28186 425174
rect 28422 424938 63866 425174
rect 64102 424938 64186 425174
rect 64422 424938 99866 425174
rect 100102 424938 100186 425174
rect 100422 424938 135866 425174
rect 136102 424938 136186 425174
rect 136422 424938 171866 425174
rect 172102 424938 172186 425174
rect 172422 424938 243866 425174
rect 244102 424938 244186 425174
rect 244422 424938 567866 425174
rect 568102 424938 568186 425174
rect 568422 424938 592062 425174
rect 592298 424938 592382 425174
rect 592618 424938 592650 425174
rect -8726 424906 592650 424938
rect -8726 421774 592650 421806
rect -8726 421538 -7734 421774
rect -7498 421538 -7414 421774
rect -7178 421538 24146 421774
rect 24382 421538 24466 421774
rect 24702 421538 60146 421774
rect 60382 421538 60466 421774
rect 60702 421538 96146 421774
rect 96382 421538 96466 421774
rect 96702 421538 132146 421774
rect 132382 421538 132466 421774
rect 132702 421538 240146 421774
rect 240382 421538 240466 421774
rect 240702 421538 564146 421774
rect 564382 421538 564466 421774
rect 564702 421538 591102 421774
rect 591338 421538 591422 421774
rect 591658 421538 592650 421774
rect -8726 421454 592650 421538
rect -8726 421218 -7734 421454
rect -7498 421218 -7414 421454
rect -7178 421218 24146 421454
rect 24382 421218 24466 421454
rect 24702 421218 60146 421454
rect 60382 421218 60466 421454
rect 60702 421218 96146 421454
rect 96382 421218 96466 421454
rect 96702 421218 132146 421454
rect 132382 421218 132466 421454
rect 132702 421218 240146 421454
rect 240382 421218 240466 421454
rect 240702 421218 564146 421454
rect 564382 421218 564466 421454
rect 564702 421218 591102 421454
rect 591338 421218 591422 421454
rect 591658 421218 592650 421454
rect -8726 421186 592650 421218
rect -8726 418054 592650 418086
rect -8726 417818 -6774 418054
rect -6538 417818 -6454 418054
rect -6218 417818 20426 418054
rect 20662 417818 20746 418054
rect 20982 417818 56426 418054
rect 56662 417818 56746 418054
rect 56982 417818 92426 418054
rect 92662 417818 92746 418054
rect 92982 417818 128426 418054
rect 128662 417818 128746 418054
rect 128982 417818 236426 418054
rect 236662 417818 236746 418054
rect 236982 417818 560426 418054
rect 560662 417818 560746 418054
rect 560982 417818 590142 418054
rect 590378 417818 590462 418054
rect 590698 417818 592650 418054
rect -8726 417734 592650 417818
rect -8726 417498 -6774 417734
rect -6538 417498 -6454 417734
rect -6218 417498 20426 417734
rect 20662 417498 20746 417734
rect 20982 417498 56426 417734
rect 56662 417498 56746 417734
rect 56982 417498 92426 417734
rect 92662 417498 92746 417734
rect 92982 417498 128426 417734
rect 128662 417498 128746 417734
rect 128982 417498 236426 417734
rect 236662 417498 236746 417734
rect 236982 417498 560426 417734
rect 560662 417498 560746 417734
rect 560982 417498 590142 417734
rect 590378 417498 590462 417734
rect 590698 417498 592650 417734
rect -8726 417466 592650 417498
rect -8726 414334 592650 414366
rect -8726 414098 -5814 414334
rect -5578 414098 -5494 414334
rect -5258 414098 16706 414334
rect 16942 414098 17026 414334
rect 17262 414098 52706 414334
rect 52942 414098 53026 414334
rect 53262 414098 88706 414334
rect 88942 414098 89026 414334
rect 89262 414098 124706 414334
rect 124942 414098 125026 414334
rect 125262 414098 232706 414334
rect 232942 414098 233026 414334
rect 233262 414098 556706 414334
rect 556942 414098 557026 414334
rect 557262 414098 589182 414334
rect 589418 414098 589502 414334
rect 589738 414098 592650 414334
rect -8726 414014 592650 414098
rect -8726 413778 -5814 414014
rect -5578 413778 -5494 414014
rect -5258 413778 16706 414014
rect 16942 413778 17026 414014
rect 17262 413778 52706 414014
rect 52942 413778 53026 414014
rect 53262 413778 88706 414014
rect 88942 413778 89026 414014
rect 89262 413778 124706 414014
rect 124942 413778 125026 414014
rect 125262 413778 232706 414014
rect 232942 413778 233026 414014
rect 233262 413778 556706 414014
rect 556942 413778 557026 414014
rect 557262 413778 589182 414014
rect 589418 413778 589502 414014
rect 589738 413778 592650 414014
rect -8726 413746 592650 413778
rect -8726 410614 592650 410646
rect -8726 410378 -4854 410614
rect -4618 410378 -4534 410614
rect -4298 410378 12986 410614
rect 13222 410378 13306 410614
rect 13542 410378 48986 410614
rect 49222 410378 49306 410614
rect 49542 410378 84986 410614
rect 85222 410378 85306 410614
rect 85542 410378 120986 410614
rect 121222 410378 121306 410614
rect 121542 410378 228986 410614
rect 229222 410378 229306 410614
rect 229542 410378 552986 410614
rect 553222 410378 553306 410614
rect 553542 410378 588222 410614
rect 588458 410378 588542 410614
rect 588778 410378 592650 410614
rect -8726 410294 592650 410378
rect -8726 410058 -4854 410294
rect -4618 410058 -4534 410294
rect -4298 410058 12986 410294
rect 13222 410058 13306 410294
rect 13542 410058 48986 410294
rect 49222 410058 49306 410294
rect 49542 410058 84986 410294
rect 85222 410058 85306 410294
rect 85542 410058 120986 410294
rect 121222 410058 121306 410294
rect 121542 410058 228986 410294
rect 229222 410058 229306 410294
rect 229542 410058 552986 410294
rect 553222 410058 553306 410294
rect 553542 410058 588222 410294
rect 588458 410058 588542 410294
rect 588778 410058 592650 410294
rect -8726 410026 592650 410058
rect -8726 406894 592650 406926
rect -8726 406658 -3894 406894
rect -3658 406658 -3574 406894
rect -3338 406658 9266 406894
rect 9502 406658 9586 406894
rect 9822 406658 45266 406894
rect 45502 406658 45586 406894
rect 45822 406658 81266 406894
rect 81502 406658 81586 406894
rect 81822 406658 117266 406894
rect 117502 406658 117586 406894
rect 117822 406658 153266 406894
rect 153502 406658 153586 406894
rect 153822 406658 225266 406894
rect 225502 406658 225586 406894
rect 225822 406658 587262 406894
rect 587498 406658 587582 406894
rect 587818 406658 592650 406894
rect -8726 406574 592650 406658
rect -8726 406338 -3894 406574
rect -3658 406338 -3574 406574
rect -3338 406338 9266 406574
rect 9502 406338 9586 406574
rect 9822 406338 45266 406574
rect 45502 406338 45586 406574
rect 45822 406338 81266 406574
rect 81502 406338 81586 406574
rect 81822 406338 117266 406574
rect 117502 406338 117586 406574
rect 117822 406338 153266 406574
rect 153502 406338 153586 406574
rect 153822 406338 225266 406574
rect 225502 406338 225586 406574
rect 225822 406338 587262 406574
rect 587498 406338 587582 406574
rect 587818 406338 592650 406574
rect -8726 406306 592650 406338
rect -8726 403174 592650 403206
rect -8726 402938 -2934 403174
rect -2698 402938 -2614 403174
rect -2378 402938 5546 403174
rect 5782 402938 5866 403174
rect 6102 402938 41546 403174
rect 41782 402938 41866 403174
rect 42102 402938 77546 403174
rect 77782 402938 77866 403174
rect 78102 402938 113546 403174
rect 113782 402938 113866 403174
rect 114102 402938 149546 403174
rect 149782 402938 149866 403174
rect 150102 402938 177610 403174
rect 177846 402938 208330 403174
rect 208566 402938 221546 403174
rect 221782 402938 221866 403174
rect 222102 402938 273210 403174
rect 273446 402938 303930 403174
rect 304166 402938 334650 403174
rect 334886 402938 365370 403174
rect 365606 402938 396090 403174
rect 396326 402938 426810 403174
rect 427046 402938 457530 403174
rect 457766 402938 488250 403174
rect 488486 402938 518970 403174
rect 519206 402938 545546 403174
rect 545782 402938 545866 403174
rect 546102 402938 549690 403174
rect 549926 402938 581546 403174
rect 581782 402938 581866 403174
rect 582102 402938 586302 403174
rect 586538 402938 586622 403174
rect 586858 402938 592650 403174
rect -8726 402854 592650 402938
rect -8726 402618 -2934 402854
rect -2698 402618 -2614 402854
rect -2378 402618 5546 402854
rect 5782 402618 5866 402854
rect 6102 402618 41546 402854
rect 41782 402618 41866 402854
rect 42102 402618 77546 402854
rect 77782 402618 77866 402854
rect 78102 402618 113546 402854
rect 113782 402618 113866 402854
rect 114102 402618 149546 402854
rect 149782 402618 149866 402854
rect 150102 402618 177610 402854
rect 177846 402618 208330 402854
rect 208566 402618 221546 402854
rect 221782 402618 221866 402854
rect 222102 402618 273210 402854
rect 273446 402618 303930 402854
rect 304166 402618 334650 402854
rect 334886 402618 365370 402854
rect 365606 402618 396090 402854
rect 396326 402618 426810 402854
rect 427046 402618 457530 402854
rect 457766 402618 488250 402854
rect 488486 402618 518970 402854
rect 519206 402618 545546 402854
rect 545782 402618 545866 402854
rect 546102 402618 549690 402854
rect 549926 402618 581546 402854
rect 581782 402618 581866 402854
rect 582102 402618 586302 402854
rect 586538 402618 586622 402854
rect 586858 402618 592650 402854
rect -8726 402586 592650 402618
rect -8726 399454 592650 399486
rect -8726 399218 -1974 399454
rect -1738 399218 -1654 399454
rect -1418 399218 1826 399454
rect 2062 399218 2146 399454
rect 2382 399218 37826 399454
rect 38062 399218 38146 399454
rect 38382 399218 73826 399454
rect 74062 399218 74146 399454
rect 74382 399218 109826 399454
rect 110062 399218 110146 399454
rect 110382 399218 145826 399454
rect 146062 399218 146146 399454
rect 146382 399218 162250 399454
rect 162486 399218 192970 399454
rect 193206 399218 217826 399454
rect 218062 399218 218146 399454
rect 218382 399218 253826 399454
rect 254062 399218 254146 399454
rect 254382 399218 257850 399454
rect 258086 399218 288570 399454
rect 288806 399218 319290 399454
rect 319526 399218 350010 399454
rect 350246 399218 380730 399454
rect 380966 399218 411450 399454
rect 411686 399218 442170 399454
rect 442406 399218 472890 399454
rect 473126 399218 503610 399454
rect 503846 399218 534330 399454
rect 534566 399218 541826 399454
rect 542062 399218 542146 399454
rect 542382 399218 565050 399454
rect 565286 399218 577826 399454
rect 578062 399218 578146 399454
rect 578382 399218 585342 399454
rect 585578 399218 585662 399454
rect 585898 399218 592650 399454
rect -8726 399134 592650 399218
rect -8726 398898 -1974 399134
rect -1738 398898 -1654 399134
rect -1418 398898 1826 399134
rect 2062 398898 2146 399134
rect 2382 398898 37826 399134
rect 38062 398898 38146 399134
rect 38382 398898 73826 399134
rect 74062 398898 74146 399134
rect 74382 398898 109826 399134
rect 110062 398898 110146 399134
rect 110382 398898 145826 399134
rect 146062 398898 146146 399134
rect 146382 398898 162250 399134
rect 162486 398898 192970 399134
rect 193206 398898 217826 399134
rect 218062 398898 218146 399134
rect 218382 398898 253826 399134
rect 254062 398898 254146 399134
rect 254382 398898 257850 399134
rect 258086 398898 288570 399134
rect 288806 398898 319290 399134
rect 319526 398898 350010 399134
rect 350246 398898 380730 399134
rect 380966 398898 411450 399134
rect 411686 398898 442170 399134
rect 442406 398898 472890 399134
rect 473126 398898 503610 399134
rect 503846 398898 534330 399134
rect 534566 398898 541826 399134
rect 542062 398898 542146 399134
rect 542382 398898 565050 399134
rect 565286 398898 577826 399134
rect 578062 398898 578146 399134
rect 578382 398898 585342 399134
rect 585578 398898 585662 399134
rect 585898 398898 592650 399134
rect -8726 398866 592650 398898
rect -8726 389494 592650 389526
rect -8726 389258 -8694 389494
rect -8458 389258 -8374 389494
rect -8138 389258 27866 389494
rect 28102 389258 28186 389494
rect 28422 389258 63866 389494
rect 64102 389258 64186 389494
rect 64422 389258 99866 389494
rect 100102 389258 100186 389494
rect 100422 389258 135866 389494
rect 136102 389258 136186 389494
rect 136422 389258 243866 389494
rect 244102 389258 244186 389494
rect 244422 389258 567866 389494
rect 568102 389258 568186 389494
rect 568422 389258 592062 389494
rect 592298 389258 592382 389494
rect 592618 389258 592650 389494
rect -8726 389174 592650 389258
rect -8726 388938 -8694 389174
rect -8458 388938 -8374 389174
rect -8138 388938 27866 389174
rect 28102 388938 28186 389174
rect 28422 388938 63866 389174
rect 64102 388938 64186 389174
rect 64422 388938 99866 389174
rect 100102 388938 100186 389174
rect 100422 388938 135866 389174
rect 136102 388938 136186 389174
rect 136422 388938 243866 389174
rect 244102 388938 244186 389174
rect 244422 388938 567866 389174
rect 568102 388938 568186 389174
rect 568422 388938 592062 389174
rect 592298 388938 592382 389174
rect 592618 388938 592650 389174
rect -8726 388906 592650 388938
rect -8726 385774 592650 385806
rect -8726 385538 -7734 385774
rect -7498 385538 -7414 385774
rect -7178 385538 24146 385774
rect 24382 385538 24466 385774
rect 24702 385538 60146 385774
rect 60382 385538 60466 385774
rect 60702 385538 96146 385774
rect 96382 385538 96466 385774
rect 96702 385538 132146 385774
rect 132382 385538 132466 385774
rect 132702 385538 240146 385774
rect 240382 385538 240466 385774
rect 240702 385538 564146 385774
rect 564382 385538 564466 385774
rect 564702 385538 591102 385774
rect 591338 385538 591422 385774
rect 591658 385538 592650 385774
rect -8726 385454 592650 385538
rect -8726 385218 -7734 385454
rect -7498 385218 -7414 385454
rect -7178 385218 24146 385454
rect 24382 385218 24466 385454
rect 24702 385218 60146 385454
rect 60382 385218 60466 385454
rect 60702 385218 96146 385454
rect 96382 385218 96466 385454
rect 96702 385218 132146 385454
rect 132382 385218 132466 385454
rect 132702 385218 240146 385454
rect 240382 385218 240466 385454
rect 240702 385218 564146 385454
rect 564382 385218 564466 385454
rect 564702 385218 591102 385454
rect 591338 385218 591422 385454
rect 591658 385218 592650 385454
rect -8726 385186 592650 385218
rect -8726 382054 592650 382086
rect -8726 381818 -6774 382054
rect -6538 381818 -6454 382054
rect -6218 381818 20426 382054
rect 20662 381818 20746 382054
rect 20982 381818 56426 382054
rect 56662 381818 56746 382054
rect 56982 381818 92426 382054
rect 92662 381818 92746 382054
rect 92982 381818 128426 382054
rect 128662 381818 128746 382054
rect 128982 381818 236426 382054
rect 236662 381818 236746 382054
rect 236982 381818 560426 382054
rect 560662 381818 560746 382054
rect 560982 381818 590142 382054
rect 590378 381818 590462 382054
rect 590698 381818 592650 382054
rect -8726 381734 592650 381818
rect -8726 381498 -6774 381734
rect -6538 381498 -6454 381734
rect -6218 381498 20426 381734
rect 20662 381498 20746 381734
rect 20982 381498 56426 381734
rect 56662 381498 56746 381734
rect 56982 381498 92426 381734
rect 92662 381498 92746 381734
rect 92982 381498 128426 381734
rect 128662 381498 128746 381734
rect 128982 381498 236426 381734
rect 236662 381498 236746 381734
rect 236982 381498 560426 381734
rect 560662 381498 560746 381734
rect 560982 381498 590142 381734
rect 590378 381498 590462 381734
rect 590698 381498 592650 381734
rect -8726 381466 592650 381498
rect -8726 378334 592650 378366
rect -8726 378098 -5814 378334
rect -5578 378098 -5494 378334
rect -5258 378098 16706 378334
rect 16942 378098 17026 378334
rect 17262 378098 52706 378334
rect 52942 378098 53026 378334
rect 53262 378098 88706 378334
rect 88942 378098 89026 378334
rect 89262 378098 124706 378334
rect 124942 378098 125026 378334
rect 125262 378098 232706 378334
rect 232942 378098 233026 378334
rect 233262 378098 268706 378334
rect 268942 378098 269026 378334
rect 269262 378098 304706 378334
rect 304942 378098 305026 378334
rect 305262 378098 340706 378334
rect 340942 378098 341026 378334
rect 341262 378098 376706 378334
rect 376942 378098 377026 378334
rect 377262 378098 412706 378334
rect 412942 378098 413026 378334
rect 413262 378098 448706 378334
rect 448942 378098 449026 378334
rect 449262 378098 484706 378334
rect 484942 378098 485026 378334
rect 485262 378098 520706 378334
rect 520942 378098 521026 378334
rect 521262 378098 556706 378334
rect 556942 378098 557026 378334
rect 557262 378098 589182 378334
rect 589418 378098 589502 378334
rect 589738 378098 592650 378334
rect -8726 378014 592650 378098
rect -8726 377778 -5814 378014
rect -5578 377778 -5494 378014
rect -5258 377778 16706 378014
rect 16942 377778 17026 378014
rect 17262 377778 52706 378014
rect 52942 377778 53026 378014
rect 53262 377778 88706 378014
rect 88942 377778 89026 378014
rect 89262 377778 124706 378014
rect 124942 377778 125026 378014
rect 125262 377778 232706 378014
rect 232942 377778 233026 378014
rect 233262 377778 268706 378014
rect 268942 377778 269026 378014
rect 269262 377778 304706 378014
rect 304942 377778 305026 378014
rect 305262 377778 340706 378014
rect 340942 377778 341026 378014
rect 341262 377778 376706 378014
rect 376942 377778 377026 378014
rect 377262 377778 412706 378014
rect 412942 377778 413026 378014
rect 413262 377778 448706 378014
rect 448942 377778 449026 378014
rect 449262 377778 484706 378014
rect 484942 377778 485026 378014
rect 485262 377778 520706 378014
rect 520942 377778 521026 378014
rect 521262 377778 556706 378014
rect 556942 377778 557026 378014
rect 557262 377778 589182 378014
rect 589418 377778 589502 378014
rect 589738 377778 592650 378014
rect -8726 377746 592650 377778
rect -8726 374614 592650 374646
rect -8726 374378 -4854 374614
rect -4618 374378 -4534 374614
rect -4298 374378 12986 374614
rect 13222 374378 13306 374614
rect 13542 374378 48986 374614
rect 49222 374378 49306 374614
rect 49542 374378 84986 374614
rect 85222 374378 85306 374614
rect 85542 374378 120986 374614
rect 121222 374378 121306 374614
rect 121542 374378 228986 374614
rect 229222 374378 229306 374614
rect 229542 374378 264986 374614
rect 265222 374378 265306 374614
rect 265542 374378 300986 374614
rect 301222 374378 301306 374614
rect 301542 374378 336986 374614
rect 337222 374378 337306 374614
rect 337542 374378 372986 374614
rect 373222 374378 373306 374614
rect 373542 374378 408986 374614
rect 409222 374378 409306 374614
rect 409542 374378 444986 374614
rect 445222 374378 445306 374614
rect 445542 374378 480986 374614
rect 481222 374378 481306 374614
rect 481542 374378 516986 374614
rect 517222 374378 517306 374614
rect 517542 374378 552986 374614
rect 553222 374378 553306 374614
rect 553542 374378 588222 374614
rect 588458 374378 588542 374614
rect 588778 374378 592650 374614
rect -8726 374294 592650 374378
rect -8726 374058 -4854 374294
rect -4618 374058 -4534 374294
rect -4298 374058 12986 374294
rect 13222 374058 13306 374294
rect 13542 374058 48986 374294
rect 49222 374058 49306 374294
rect 49542 374058 84986 374294
rect 85222 374058 85306 374294
rect 85542 374058 120986 374294
rect 121222 374058 121306 374294
rect 121542 374058 228986 374294
rect 229222 374058 229306 374294
rect 229542 374058 264986 374294
rect 265222 374058 265306 374294
rect 265542 374058 300986 374294
rect 301222 374058 301306 374294
rect 301542 374058 336986 374294
rect 337222 374058 337306 374294
rect 337542 374058 372986 374294
rect 373222 374058 373306 374294
rect 373542 374058 408986 374294
rect 409222 374058 409306 374294
rect 409542 374058 444986 374294
rect 445222 374058 445306 374294
rect 445542 374058 480986 374294
rect 481222 374058 481306 374294
rect 481542 374058 516986 374294
rect 517222 374058 517306 374294
rect 517542 374058 552986 374294
rect 553222 374058 553306 374294
rect 553542 374058 588222 374294
rect 588458 374058 588542 374294
rect 588778 374058 592650 374294
rect -8726 374026 592650 374058
rect -8726 370894 592650 370926
rect -8726 370658 -3894 370894
rect -3658 370658 -3574 370894
rect -3338 370658 9266 370894
rect 9502 370658 9586 370894
rect 9822 370658 45266 370894
rect 45502 370658 45586 370894
rect 45822 370658 81266 370894
rect 81502 370658 81586 370894
rect 81822 370658 117266 370894
rect 117502 370658 117586 370894
rect 117822 370658 153266 370894
rect 153502 370658 153586 370894
rect 153822 370658 225266 370894
rect 225502 370658 225586 370894
rect 225822 370658 261266 370894
rect 261502 370658 261586 370894
rect 261822 370658 297266 370894
rect 297502 370658 297586 370894
rect 297822 370658 333266 370894
rect 333502 370658 333586 370894
rect 333822 370658 369266 370894
rect 369502 370658 369586 370894
rect 369822 370658 405266 370894
rect 405502 370658 405586 370894
rect 405822 370658 441266 370894
rect 441502 370658 441586 370894
rect 441822 370658 477266 370894
rect 477502 370658 477586 370894
rect 477822 370658 513266 370894
rect 513502 370658 513586 370894
rect 513822 370658 549266 370894
rect 549502 370658 549586 370894
rect 549822 370658 587262 370894
rect 587498 370658 587582 370894
rect 587818 370658 592650 370894
rect -8726 370574 592650 370658
rect -8726 370338 -3894 370574
rect -3658 370338 -3574 370574
rect -3338 370338 9266 370574
rect 9502 370338 9586 370574
rect 9822 370338 45266 370574
rect 45502 370338 45586 370574
rect 45822 370338 81266 370574
rect 81502 370338 81586 370574
rect 81822 370338 117266 370574
rect 117502 370338 117586 370574
rect 117822 370338 153266 370574
rect 153502 370338 153586 370574
rect 153822 370338 225266 370574
rect 225502 370338 225586 370574
rect 225822 370338 261266 370574
rect 261502 370338 261586 370574
rect 261822 370338 297266 370574
rect 297502 370338 297586 370574
rect 297822 370338 333266 370574
rect 333502 370338 333586 370574
rect 333822 370338 369266 370574
rect 369502 370338 369586 370574
rect 369822 370338 405266 370574
rect 405502 370338 405586 370574
rect 405822 370338 441266 370574
rect 441502 370338 441586 370574
rect 441822 370338 477266 370574
rect 477502 370338 477586 370574
rect 477822 370338 513266 370574
rect 513502 370338 513586 370574
rect 513822 370338 549266 370574
rect 549502 370338 549586 370574
rect 549822 370338 587262 370574
rect 587498 370338 587582 370574
rect 587818 370338 592650 370574
rect -8726 370306 592650 370338
rect -8726 367174 592650 367206
rect -8726 366938 -2934 367174
rect -2698 366938 -2614 367174
rect -2378 366938 5546 367174
rect 5782 366938 5866 367174
rect 6102 366938 41546 367174
rect 41782 366938 41866 367174
rect 42102 366938 77546 367174
rect 77782 366938 77866 367174
rect 78102 366938 113546 367174
rect 113782 366938 113866 367174
rect 114102 366938 149546 367174
rect 149782 366938 149866 367174
rect 150102 366938 177610 367174
rect 177846 366938 208330 367174
rect 208566 366938 221546 367174
rect 221782 366938 221866 367174
rect 222102 366938 257546 367174
rect 257782 366938 257866 367174
rect 258102 366938 293546 367174
rect 293782 366938 293866 367174
rect 294102 366938 329546 367174
rect 329782 366938 329866 367174
rect 330102 366938 365546 367174
rect 365782 366938 365866 367174
rect 366102 366938 401546 367174
rect 401782 366938 401866 367174
rect 402102 366938 437546 367174
rect 437782 366938 437866 367174
rect 438102 366938 473546 367174
rect 473782 366938 473866 367174
rect 474102 366938 509546 367174
rect 509782 366938 509866 367174
rect 510102 366938 545546 367174
rect 545782 366938 545866 367174
rect 546102 366938 581546 367174
rect 581782 366938 581866 367174
rect 582102 366938 586302 367174
rect 586538 366938 586622 367174
rect 586858 366938 592650 367174
rect -8726 366854 592650 366938
rect -8726 366618 -2934 366854
rect -2698 366618 -2614 366854
rect -2378 366618 5546 366854
rect 5782 366618 5866 366854
rect 6102 366618 41546 366854
rect 41782 366618 41866 366854
rect 42102 366618 77546 366854
rect 77782 366618 77866 366854
rect 78102 366618 113546 366854
rect 113782 366618 113866 366854
rect 114102 366618 149546 366854
rect 149782 366618 149866 366854
rect 150102 366618 177610 366854
rect 177846 366618 208330 366854
rect 208566 366618 221546 366854
rect 221782 366618 221866 366854
rect 222102 366618 257546 366854
rect 257782 366618 257866 366854
rect 258102 366618 293546 366854
rect 293782 366618 293866 366854
rect 294102 366618 329546 366854
rect 329782 366618 329866 366854
rect 330102 366618 365546 366854
rect 365782 366618 365866 366854
rect 366102 366618 401546 366854
rect 401782 366618 401866 366854
rect 402102 366618 437546 366854
rect 437782 366618 437866 366854
rect 438102 366618 473546 366854
rect 473782 366618 473866 366854
rect 474102 366618 509546 366854
rect 509782 366618 509866 366854
rect 510102 366618 545546 366854
rect 545782 366618 545866 366854
rect 546102 366618 581546 366854
rect 581782 366618 581866 366854
rect 582102 366618 586302 366854
rect 586538 366618 586622 366854
rect 586858 366618 592650 366854
rect -8726 366586 592650 366618
rect -8726 363454 592650 363486
rect -8726 363218 -1974 363454
rect -1738 363218 -1654 363454
rect -1418 363218 1826 363454
rect 2062 363218 2146 363454
rect 2382 363218 37826 363454
rect 38062 363218 38146 363454
rect 38382 363218 73826 363454
rect 74062 363218 74146 363454
rect 74382 363218 109826 363454
rect 110062 363218 110146 363454
rect 110382 363218 145826 363454
rect 146062 363218 146146 363454
rect 146382 363218 162250 363454
rect 162486 363218 192970 363454
rect 193206 363218 217826 363454
rect 218062 363218 218146 363454
rect 218382 363218 253826 363454
rect 254062 363218 254146 363454
rect 254382 363218 289826 363454
rect 290062 363218 290146 363454
rect 290382 363218 325826 363454
rect 326062 363218 326146 363454
rect 326382 363218 361826 363454
rect 362062 363218 362146 363454
rect 362382 363218 397826 363454
rect 398062 363218 398146 363454
rect 398382 363218 433826 363454
rect 434062 363218 434146 363454
rect 434382 363218 469826 363454
rect 470062 363218 470146 363454
rect 470382 363218 505826 363454
rect 506062 363218 506146 363454
rect 506382 363218 541826 363454
rect 542062 363218 542146 363454
rect 542382 363218 577826 363454
rect 578062 363218 578146 363454
rect 578382 363218 585342 363454
rect 585578 363218 585662 363454
rect 585898 363218 592650 363454
rect -8726 363134 592650 363218
rect -8726 362898 -1974 363134
rect -1738 362898 -1654 363134
rect -1418 362898 1826 363134
rect 2062 362898 2146 363134
rect 2382 362898 37826 363134
rect 38062 362898 38146 363134
rect 38382 362898 73826 363134
rect 74062 362898 74146 363134
rect 74382 362898 109826 363134
rect 110062 362898 110146 363134
rect 110382 362898 145826 363134
rect 146062 362898 146146 363134
rect 146382 362898 162250 363134
rect 162486 362898 192970 363134
rect 193206 362898 217826 363134
rect 218062 362898 218146 363134
rect 218382 362898 253826 363134
rect 254062 362898 254146 363134
rect 254382 362898 289826 363134
rect 290062 362898 290146 363134
rect 290382 362898 325826 363134
rect 326062 362898 326146 363134
rect 326382 362898 361826 363134
rect 362062 362898 362146 363134
rect 362382 362898 397826 363134
rect 398062 362898 398146 363134
rect 398382 362898 433826 363134
rect 434062 362898 434146 363134
rect 434382 362898 469826 363134
rect 470062 362898 470146 363134
rect 470382 362898 505826 363134
rect 506062 362898 506146 363134
rect 506382 362898 541826 363134
rect 542062 362898 542146 363134
rect 542382 362898 577826 363134
rect 578062 362898 578146 363134
rect 578382 362898 585342 363134
rect 585578 362898 585662 363134
rect 585898 362898 592650 363134
rect -8726 362866 592650 362898
rect -8726 353494 592650 353526
rect -8726 353258 -8694 353494
rect -8458 353258 -8374 353494
rect -8138 353258 27866 353494
rect 28102 353258 28186 353494
rect 28422 353258 63866 353494
rect 64102 353258 64186 353494
rect 64422 353258 99866 353494
rect 100102 353258 100186 353494
rect 100422 353258 135866 353494
rect 136102 353258 136186 353494
rect 136422 353258 243866 353494
rect 244102 353258 244186 353494
rect 244422 353258 567866 353494
rect 568102 353258 568186 353494
rect 568422 353258 592062 353494
rect 592298 353258 592382 353494
rect 592618 353258 592650 353494
rect -8726 353174 592650 353258
rect -8726 352938 -8694 353174
rect -8458 352938 -8374 353174
rect -8138 352938 27866 353174
rect 28102 352938 28186 353174
rect 28422 352938 63866 353174
rect 64102 352938 64186 353174
rect 64422 352938 99866 353174
rect 100102 352938 100186 353174
rect 100422 352938 135866 353174
rect 136102 352938 136186 353174
rect 136422 352938 243866 353174
rect 244102 352938 244186 353174
rect 244422 352938 567866 353174
rect 568102 352938 568186 353174
rect 568422 352938 592062 353174
rect 592298 352938 592382 353174
rect 592618 352938 592650 353174
rect -8726 352906 592650 352938
rect -8726 349774 592650 349806
rect -8726 349538 -7734 349774
rect -7498 349538 -7414 349774
rect -7178 349538 24146 349774
rect 24382 349538 24466 349774
rect 24702 349538 60146 349774
rect 60382 349538 60466 349774
rect 60702 349538 96146 349774
rect 96382 349538 96466 349774
rect 96702 349538 132146 349774
rect 132382 349538 132466 349774
rect 132702 349538 240146 349774
rect 240382 349538 240466 349774
rect 240702 349538 564146 349774
rect 564382 349538 564466 349774
rect 564702 349538 591102 349774
rect 591338 349538 591422 349774
rect 591658 349538 592650 349774
rect -8726 349454 592650 349538
rect -8726 349218 -7734 349454
rect -7498 349218 -7414 349454
rect -7178 349218 24146 349454
rect 24382 349218 24466 349454
rect 24702 349218 60146 349454
rect 60382 349218 60466 349454
rect 60702 349218 96146 349454
rect 96382 349218 96466 349454
rect 96702 349218 132146 349454
rect 132382 349218 132466 349454
rect 132702 349218 240146 349454
rect 240382 349218 240466 349454
rect 240702 349218 564146 349454
rect 564382 349218 564466 349454
rect 564702 349218 591102 349454
rect 591338 349218 591422 349454
rect 591658 349218 592650 349454
rect -8726 349186 592650 349218
rect -8726 346054 592650 346086
rect -8726 345818 -6774 346054
rect -6538 345818 -6454 346054
rect -6218 345818 20426 346054
rect 20662 345818 20746 346054
rect 20982 345818 56426 346054
rect 56662 345818 56746 346054
rect 56982 345818 92426 346054
rect 92662 345818 92746 346054
rect 92982 345818 128426 346054
rect 128662 345818 128746 346054
rect 128982 345818 236426 346054
rect 236662 345818 236746 346054
rect 236982 345818 560426 346054
rect 560662 345818 560746 346054
rect 560982 345818 590142 346054
rect 590378 345818 590462 346054
rect 590698 345818 592650 346054
rect -8726 345734 592650 345818
rect -8726 345498 -6774 345734
rect -6538 345498 -6454 345734
rect -6218 345498 20426 345734
rect 20662 345498 20746 345734
rect 20982 345498 56426 345734
rect 56662 345498 56746 345734
rect 56982 345498 92426 345734
rect 92662 345498 92746 345734
rect 92982 345498 128426 345734
rect 128662 345498 128746 345734
rect 128982 345498 236426 345734
rect 236662 345498 236746 345734
rect 236982 345498 560426 345734
rect 560662 345498 560746 345734
rect 560982 345498 590142 345734
rect 590378 345498 590462 345734
rect 590698 345498 592650 345734
rect -8726 345466 592650 345498
rect -8726 342334 592650 342366
rect -8726 342098 -5814 342334
rect -5578 342098 -5494 342334
rect -5258 342098 16706 342334
rect 16942 342098 17026 342334
rect 17262 342098 52706 342334
rect 52942 342098 53026 342334
rect 53262 342098 88706 342334
rect 88942 342098 89026 342334
rect 89262 342098 124706 342334
rect 124942 342098 125026 342334
rect 125262 342098 232706 342334
rect 232942 342098 233026 342334
rect 233262 342098 268706 342334
rect 268942 342098 269026 342334
rect 269262 342098 304706 342334
rect 304942 342098 305026 342334
rect 305262 342098 340706 342334
rect 340942 342098 341026 342334
rect 341262 342098 376706 342334
rect 376942 342098 377026 342334
rect 377262 342098 412706 342334
rect 412942 342098 413026 342334
rect 413262 342098 448706 342334
rect 448942 342098 449026 342334
rect 449262 342098 484706 342334
rect 484942 342098 485026 342334
rect 485262 342098 520706 342334
rect 520942 342098 521026 342334
rect 521262 342098 556706 342334
rect 556942 342098 557026 342334
rect 557262 342098 589182 342334
rect 589418 342098 589502 342334
rect 589738 342098 592650 342334
rect -8726 342014 592650 342098
rect -8726 341778 -5814 342014
rect -5578 341778 -5494 342014
rect -5258 341778 16706 342014
rect 16942 341778 17026 342014
rect 17262 341778 52706 342014
rect 52942 341778 53026 342014
rect 53262 341778 88706 342014
rect 88942 341778 89026 342014
rect 89262 341778 124706 342014
rect 124942 341778 125026 342014
rect 125262 341778 232706 342014
rect 232942 341778 233026 342014
rect 233262 341778 268706 342014
rect 268942 341778 269026 342014
rect 269262 341778 304706 342014
rect 304942 341778 305026 342014
rect 305262 341778 340706 342014
rect 340942 341778 341026 342014
rect 341262 341778 376706 342014
rect 376942 341778 377026 342014
rect 377262 341778 412706 342014
rect 412942 341778 413026 342014
rect 413262 341778 448706 342014
rect 448942 341778 449026 342014
rect 449262 341778 484706 342014
rect 484942 341778 485026 342014
rect 485262 341778 520706 342014
rect 520942 341778 521026 342014
rect 521262 341778 556706 342014
rect 556942 341778 557026 342014
rect 557262 341778 589182 342014
rect 589418 341778 589502 342014
rect 589738 341778 592650 342014
rect -8726 341746 592650 341778
rect -8726 338614 592650 338646
rect -8726 338378 -4854 338614
rect -4618 338378 -4534 338614
rect -4298 338378 12986 338614
rect 13222 338378 13306 338614
rect 13542 338378 48986 338614
rect 49222 338378 49306 338614
rect 49542 338378 84986 338614
rect 85222 338378 85306 338614
rect 85542 338378 120986 338614
rect 121222 338378 121306 338614
rect 121542 338378 228986 338614
rect 229222 338378 229306 338614
rect 229542 338378 264986 338614
rect 265222 338378 265306 338614
rect 265542 338378 300986 338614
rect 301222 338378 301306 338614
rect 301542 338378 336986 338614
rect 337222 338378 337306 338614
rect 337542 338378 372986 338614
rect 373222 338378 373306 338614
rect 373542 338378 408986 338614
rect 409222 338378 409306 338614
rect 409542 338378 444986 338614
rect 445222 338378 445306 338614
rect 445542 338378 480986 338614
rect 481222 338378 481306 338614
rect 481542 338378 516986 338614
rect 517222 338378 517306 338614
rect 517542 338378 552986 338614
rect 553222 338378 553306 338614
rect 553542 338378 588222 338614
rect 588458 338378 588542 338614
rect 588778 338378 592650 338614
rect -8726 338294 592650 338378
rect -8726 338058 -4854 338294
rect -4618 338058 -4534 338294
rect -4298 338058 12986 338294
rect 13222 338058 13306 338294
rect 13542 338058 48986 338294
rect 49222 338058 49306 338294
rect 49542 338058 84986 338294
rect 85222 338058 85306 338294
rect 85542 338058 120986 338294
rect 121222 338058 121306 338294
rect 121542 338058 228986 338294
rect 229222 338058 229306 338294
rect 229542 338058 264986 338294
rect 265222 338058 265306 338294
rect 265542 338058 300986 338294
rect 301222 338058 301306 338294
rect 301542 338058 336986 338294
rect 337222 338058 337306 338294
rect 337542 338058 372986 338294
rect 373222 338058 373306 338294
rect 373542 338058 408986 338294
rect 409222 338058 409306 338294
rect 409542 338058 444986 338294
rect 445222 338058 445306 338294
rect 445542 338058 480986 338294
rect 481222 338058 481306 338294
rect 481542 338058 516986 338294
rect 517222 338058 517306 338294
rect 517542 338058 552986 338294
rect 553222 338058 553306 338294
rect 553542 338058 588222 338294
rect 588458 338058 588542 338294
rect 588778 338058 592650 338294
rect -8726 338026 592650 338058
rect -8726 334894 592650 334926
rect -8726 334658 -3894 334894
rect -3658 334658 -3574 334894
rect -3338 334658 9266 334894
rect 9502 334658 9586 334894
rect 9822 334658 45266 334894
rect 45502 334658 45586 334894
rect 45822 334658 81266 334894
rect 81502 334658 81586 334894
rect 81822 334658 117266 334894
rect 117502 334658 117586 334894
rect 117822 334658 153266 334894
rect 153502 334658 153586 334894
rect 153822 334658 225266 334894
rect 225502 334658 225586 334894
rect 225822 334658 261266 334894
rect 261502 334658 261586 334894
rect 261822 334658 297266 334894
rect 297502 334658 297586 334894
rect 297822 334658 333266 334894
rect 333502 334658 333586 334894
rect 333822 334658 369266 334894
rect 369502 334658 369586 334894
rect 369822 334658 405266 334894
rect 405502 334658 405586 334894
rect 405822 334658 441266 334894
rect 441502 334658 441586 334894
rect 441822 334658 477266 334894
rect 477502 334658 477586 334894
rect 477822 334658 513266 334894
rect 513502 334658 513586 334894
rect 513822 334658 549266 334894
rect 549502 334658 549586 334894
rect 549822 334658 587262 334894
rect 587498 334658 587582 334894
rect 587818 334658 592650 334894
rect -8726 334574 592650 334658
rect -8726 334338 -3894 334574
rect -3658 334338 -3574 334574
rect -3338 334338 9266 334574
rect 9502 334338 9586 334574
rect 9822 334338 45266 334574
rect 45502 334338 45586 334574
rect 45822 334338 81266 334574
rect 81502 334338 81586 334574
rect 81822 334338 117266 334574
rect 117502 334338 117586 334574
rect 117822 334338 153266 334574
rect 153502 334338 153586 334574
rect 153822 334338 225266 334574
rect 225502 334338 225586 334574
rect 225822 334338 261266 334574
rect 261502 334338 261586 334574
rect 261822 334338 297266 334574
rect 297502 334338 297586 334574
rect 297822 334338 333266 334574
rect 333502 334338 333586 334574
rect 333822 334338 369266 334574
rect 369502 334338 369586 334574
rect 369822 334338 405266 334574
rect 405502 334338 405586 334574
rect 405822 334338 441266 334574
rect 441502 334338 441586 334574
rect 441822 334338 477266 334574
rect 477502 334338 477586 334574
rect 477822 334338 513266 334574
rect 513502 334338 513586 334574
rect 513822 334338 549266 334574
rect 549502 334338 549586 334574
rect 549822 334338 587262 334574
rect 587498 334338 587582 334574
rect 587818 334338 592650 334574
rect -8726 334306 592650 334338
rect -8726 331174 592650 331206
rect -8726 330938 -2934 331174
rect -2698 330938 -2614 331174
rect -2378 330938 5546 331174
rect 5782 330938 5866 331174
rect 6102 330938 41546 331174
rect 41782 330938 41866 331174
rect 42102 330938 77546 331174
rect 77782 330938 77866 331174
rect 78102 330938 113546 331174
rect 113782 330938 113866 331174
rect 114102 330938 149546 331174
rect 149782 330938 149866 331174
rect 150102 330938 177610 331174
rect 177846 330938 208330 331174
rect 208566 330938 221546 331174
rect 221782 330938 221866 331174
rect 222102 330938 257546 331174
rect 257782 330938 257866 331174
rect 258102 330938 293546 331174
rect 293782 330938 293866 331174
rect 294102 330938 329546 331174
rect 329782 330938 329866 331174
rect 330102 330938 365546 331174
rect 365782 330938 365866 331174
rect 366102 330938 401546 331174
rect 401782 330938 401866 331174
rect 402102 330938 437546 331174
rect 437782 330938 437866 331174
rect 438102 330938 473546 331174
rect 473782 330938 473866 331174
rect 474102 330938 509546 331174
rect 509782 330938 509866 331174
rect 510102 330938 545546 331174
rect 545782 330938 545866 331174
rect 546102 330938 581546 331174
rect 581782 330938 581866 331174
rect 582102 330938 586302 331174
rect 586538 330938 586622 331174
rect 586858 330938 592650 331174
rect -8726 330854 592650 330938
rect -8726 330618 -2934 330854
rect -2698 330618 -2614 330854
rect -2378 330618 5546 330854
rect 5782 330618 5866 330854
rect 6102 330618 41546 330854
rect 41782 330618 41866 330854
rect 42102 330618 77546 330854
rect 77782 330618 77866 330854
rect 78102 330618 113546 330854
rect 113782 330618 113866 330854
rect 114102 330618 149546 330854
rect 149782 330618 149866 330854
rect 150102 330618 177610 330854
rect 177846 330618 208330 330854
rect 208566 330618 221546 330854
rect 221782 330618 221866 330854
rect 222102 330618 257546 330854
rect 257782 330618 257866 330854
rect 258102 330618 293546 330854
rect 293782 330618 293866 330854
rect 294102 330618 329546 330854
rect 329782 330618 329866 330854
rect 330102 330618 365546 330854
rect 365782 330618 365866 330854
rect 366102 330618 401546 330854
rect 401782 330618 401866 330854
rect 402102 330618 437546 330854
rect 437782 330618 437866 330854
rect 438102 330618 473546 330854
rect 473782 330618 473866 330854
rect 474102 330618 509546 330854
rect 509782 330618 509866 330854
rect 510102 330618 545546 330854
rect 545782 330618 545866 330854
rect 546102 330618 581546 330854
rect 581782 330618 581866 330854
rect 582102 330618 586302 330854
rect 586538 330618 586622 330854
rect 586858 330618 592650 330854
rect -8726 330586 592650 330618
rect -8726 327454 592650 327486
rect -8726 327218 -1974 327454
rect -1738 327218 -1654 327454
rect -1418 327218 1826 327454
rect 2062 327218 2146 327454
rect 2382 327218 37826 327454
rect 38062 327218 38146 327454
rect 38382 327218 73826 327454
rect 74062 327218 74146 327454
rect 74382 327218 109826 327454
rect 110062 327218 110146 327454
rect 110382 327218 145826 327454
rect 146062 327218 146146 327454
rect 146382 327218 162250 327454
rect 162486 327218 192970 327454
rect 193206 327218 217826 327454
rect 218062 327218 218146 327454
rect 218382 327218 253826 327454
rect 254062 327218 254146 327454
rect 254382 327218 289826 327454
rect 290062 327218 290146 327454
rect 290382 327218 325826 327454
rect 326062 327218 326146 327454
rect 326382 327218 361826 327454
rect 362062 327218 362146 327454
rect 362382 327218 397826 327454
rect 398062 327218 398146 327454
rect 398382 327218 433826 327454
rect 434062 327218 434146 327454
rect 434382 327218 469826 327454
rect 470062 327218 470146 327454
rect 470382 327218 505826 327454
rect 506062 327218 506146 327454
rect 506382 327218 541826 327454
rect 542062 327218 542146 327454
rect 542382 327218 577826 327454
rect 578062 327218 578146 327454
rect 578382 327218 585342 327454
rect 585578 327218 585662 327454
rect 585898 327218 592650 327454
rect -8726 327134 592650 327218
rect -8726 326898 -1974 327134
rect -1738 326898 -1654 327134
rect -1418 326898 1826 327134
rect 2062 326898 2146 327134
rect 2382 326898 37826 327134
rect 38062 326898 38146 327134
rect 38382 326898 73826 327134
rect 74062 326898 74146 327134
rect 74382 326898 109826 327134
rect 110062 326898 110146 327134
rect 110382 326898 145826 327134
rect 146062 326898 146146 327134
rect 146382 326898 162250 327134
rect 162486 326898 192970 327134
rect 193206 326898 217826 327134
rect 218062 326898 218146 327134
rect 218382 326898 253826 327134
rect 254062 326898 254146 327134
rect 254382 326898 289826 327134
rect 290062 326898 290146 327134
rect 290382 326898 325826 327134
rect 326062 326898 326146 327134
rect 326382 326898 361826 327134
rect 362062 326898 362146 327134
rect 362382 326898 397826 327134
rect 398062 326898 398146 327134
rect 398382 326898 433826 327134
rect 434062 326898 434146 327134
rect 434382 326898 469826 327134
rect 470062 326898 470146 327134
rect 470382 326898 505826 327134
rect 506062 326898 506146 327134
rect 506382 326898 541826 327134
rect 542062 326898 542146 327134
rect 542382 326898 577826 327134
rect 578062 326898 578146 327134
rect 578382 326898 585342 327134
rect 585578 326898 585662 327134
rect 585898 326898 592650 327134
rect -8726 326866 592650 326898
rect -8726 317494 592650 317526
rect -8726 317258 -8694 317494
rect -8458 317258 -8374 317494
rect -8138 317258 27866 317494
rect 28102 317258 28186 317494
rect 28422 317258 135866 317494
rect 136102 317258 136186 317494
rect 136422 317258 243866 317494
rect 244102 317258 244186 317494
rect 244422 317258 567866 317494
rect 568102 317258 568186 317494
rect 568422 317258 592062 317494
rect 592298 317258 592382 317494
rect 592618 317258 592650 317494
rect -8726 317174 592650 317258
rect -8726 316938 -8694 317174
rect -8458 316938 -8374 317174
rect -8138 316938 27866 317174
rect 28102 316938 28186 317174
rect 28422 316938 135866 317174
rect 136102 316938 136186 317174
rect 136422 316938 243866 317174
rect 244102 316938 244186 317174
rect 244422 316938 567866 317174
rect 568102 316938 568186 317174
rect 568422 316938 592062 317174
rect 592298 316938 592382 317174
rect 592618 316938 592650 317174
rect -8726 316906 592650 316938
rect -8726 313774 592650 313806
rect -8726 313538 -7734 313774
rect -7498 313538 -7414 313774
rect -7178 313538 24146 313774
rect 24382 313538 24466 313774
rect 24702 313538 60146 313774
rect 60382 313538 60466 313774
rect 60702 313538 132146 313774
rect 132382 313538 132466 313774
rect 132702 313538 240146 313774
rect 240382 313538 240466 313774
rect 240702 313538 564146 313774
rect 564382 313538 564466 313774
rect 564702 313538 591102 313774
rect 591338 313538 591422 313774
rect 591658 313538 592650 313774
rect -8726 313454 592650 313538
rect -8726 313218 -7734 313454
rect -7498 313218 -7414 313454
rect -7178 313218 24146 313454
rect 24382 313218 24466 313454
rect 24702 313218 60146 313454
rect 60382 313218 60466 313454
rect 60702 313218 132146 313454
rect 132382 313218 132466 313454
rect 132702 313218 240146 313454
rect 240382 313218 240466 313454
rect 240702 313218 564146 313454
rect 564382 313218 564466 313454
rect 564702 313218 591102 313454
rect 591338 313218 591422 313454
rect 591658 313218 592650 313454
rect -8726 313186 592650 313218
rect -8726 310054 592650 310086
rect -8726 309818 -6774 310054
rect -6538 309818 -6454 310054
rect -6218 309818 20426 310054
rect 20662 309818 20746 310054
rect 20982 309818 56426 310054
rect 56662 309818 56746 310054
rect 56982 309818 128426 310054
rect 128662 309818 128746 310054
rect 128982 309818 236426 310054
rect 236662 309818 236746 310054
rect 236982 309818 560426 310054
rect 560662 309818 560746 310054
rect 560982 309818 590142 310054
rect 590378 309818 590462 310054
rect 590698 309818 592650 310054
rect -8726 309734 592650 309818
rect -8726 309498 -6774 309734
rect -6538 309498 -6454 309734
rect -6218 309498 20426 309734
rect 20662 309498 20746 309734
rect 20982 309498 56426 309734
rect 56662 309498 56746 309734
rect 56982 309498 128426 309734
rect 128662 309498 128746 309734
rect 128982 309498 236426 309734
rect 236662 309498 236746 309734
rect 236982 309498 560426 309734
rect 560662 309498 560746 309734
rect 560982 309498 590142 309734
rect 590378 309498 590462 309734
rect 590698 309498 592650 309734
rect -8726 309466 592650 309498
rect -8726 306334 592650 306366
rect -8726 306098 -5814 306334
rect -5578 306098 -5494 306334
rect -5258 306098 16706 306334
rect 16942 306098 17026 306334
rect 17262 306098 52706 306334
rect 52942 306098 53026 306334
rect 53262 306098 124706 306334
rect 124942 306098 125026 306334
rect 125262 306098 232706 306334
rect 232942 306098 233026 306334
rect 233262 306098 556706 306334
rect 556942 306098 557026 306334
rect 557262 306098 589182 306334
rect 589418 306098 589502 306334
rect 589738 306098 592650 306334
rect -8726 306014 592650 306098
rect -8726 305778 -5814 306014
rect -5578 305778 -5494 306014
rect -5258 305778 16706 306014
rect 16942 305778 17026 306014
rect 17262 305778 52706 306014
rect 52942 305778 53026 306014
rect 53262 305778 124706 306014
rect 124942 305778 125026 306014
rect 125262 305778 232706 306014
rect 232942 305778 233026 306014
rect 233262 305778 556706 306014
rect 556942 305778 557026 306014
rect 557262 305778 589182 306014
rect 589418 305778 589502 306014
rect 589738 305778 592650 306014
rect -8726 305746 592650 305778
rect -8726 302614 592650 302646
rect -8726 302378 -4854 302614
rect -4618 302378 -4534 302614
rect -4298 302378 12986 302614
rect 13222 302378 13306 302614
rect 13542 302378 120986 302614
rect 121222 302378 121306 302614
rect 121542 302378 228986 302614
rect 229222 302378 229306 302614
rect 229542 302378 552986 302614
rect 553222 302378 553306 302614
rect 553542 302378 588222 302614
rect 588458 302378 588542 302614
rect 588778 302378 592650 302614
rect -8726 302294 592650 302378
rect -8726 302058 -4854 302294
rect -4618 302058 -4534 302294
rect -4298 302058 12986 302294
rect 13222 302058 13306 302294
rect 13542 302058 120986 302294
rect 121222 302058 121306 302294
rect 121542 302058 228986 302294
rect 229222 302058 229306 302294
rect 229542 302058 552986 302294
rect 553222 302058 553306 302294
rect 553542 302058 588222 302294
rect 588458 302058 588542 302294
rect 588778 302058 592650 302294
rect -8726 302026 592650 302058
rect -8726 298894 592650 298926
rect -8726 298658 -3894 298894
rect -3658 298658 -3574 298894
rect -3338 298658 9266 298894
rect 9502 298658 9586 298894
rect 9822 298658 45266 298894
rect 45502 298658 45586 298894
rect 45822 298658 117266 298894
rect 117502 298658 117586 298894
rect 117822 298658 153266 298894
rect 153502 298658 153586 298894
rect 153822 298658 225266 298894
rect 225502 298658 225586 298894
rect 225822 298658 587262 298894
rect 587498 298658 587582 298894
rect 587818 298658 592650 298894
rect -8726 298574 592650 298658
rect -8726 298338 -3894 298574
rect -3658 298338 -3574 298574
rect -3338 298338 9266 298574
rect 9502 298338 9586 298574
rect 9822 298338 45266 298574
rect 45502 298338 45586 298574
rect 45822 298338 117266 298574
rect 117502 298338 117586 298574
rect 117822 298338 153266 298574
rect 153502 298338 153586 298574
rect 153822 298338 225266 298574
rect 225502 298338 225586 298574
rect 225822 298338 587262 298574
rect 587498 298338 587582 298574
rect 587818 298338 592650 298574
rect -8726 298306 592650 298338
rect -8726 295174 592650 295206
rect -8726 294938 -2934 295174
rect -2698 294938 -2614 295174
rect -2378 294938 5546 295174
rect 5782 294938 5866 295174
rect 6102 294938 41546 295174
rect 41782 294938 41866 295174
rect 42102 294938 49610 295174
rect 49846 294938 80330 295174
rect 80566 294938 113546 295174
rect 113782 294938 113866 295174
rect 114102 294938 149546 295174
rect 149782 294938 149866 295174
rect 150102 294938 177610 295174
rect 177846 294938 208330 295174
rect 208566 294938 221546 295174
rect 221782 294938 221866 295174
rect 222102 294938 257546 295174
rect 257782 294938 257866 295174
rect 258102 294938 279610 295174
rect 279846 294938 310330 295174
rect 310566 294938 341050 295174
rect 341286 294938 371770 295174
rect 372006 294938 402490 295174
rect 402726 294938 433210 295174
rect 433446 294938 463930 295174
rect 464166 294938 494650 295174
rect 494886 294938 525370 295174
rect 525606 294938 581546 295174
rect 581782 294938 581866 295174
rect 582102 294938 586302 295174
rect 586538 294938 586622 295174
rect 586858 294938 592650 295174
rect -8726 294854 592650 294938
rect -8726 294618 -2934 294854
rect -2698 294618 -2614 294854
rect -2378 294618 5546 294854
rect 5782 294618 5866 294854
rect 6102 294618 41546 294854
rect 41782 294618 41866 294854
rect 42102 294618 49610 294854
rect 49846 294618 80330 294854
rect 80566 294618 113546 294854
rect 113782 294618 113866 294854
rect 114102 294618 149546 294854
rect 149782 294618 149866 294854
rect 150102 294618 177610 294854
rect 177846 294618 208330 294854
rect 208566 294618 221546 294854
rect 221782 294618 221866 294854
rect 222102 294618 257546 294854
rect 257782 294618 257866 294854
rect 258102 294618 279610 294854
rect 279846 294618 310330 294854
rect 310566 294618 341050 294854
rect 341286 294618 371770 294854
rect 372006 294618 402490 294854
rect 402726 294618 433210 294854
rect 433446 294618 463930 294854
rect 464166 294618 494650 294854
rect 494886 294618 525370 294854
rect 525606 294618 581546 294854
rect 581782 294618 581866 294854
rect 582102 294618 586302 294854
rect 586538 294618 586622 294854
rect 586858 294618 592650 294854
rect -8726 294586 592650 294618
rect -8726 291454 592650 291486
rect -8726 291218 -1974 291454
rect -1738 291218 -1654 291454
rect -1418 291218 1826 291454
rect 2062 291218 2146 291454
rect 2382 291218 34250 291454
rect 34486 291218 37826 291454
rect 38062 291218 38146 291454
rect 38382 291218 64970 291454
rect 65206 291218 95690 291454
rect 95926 291218 109826 291454
rect 110062 291218 110146 291454
rect 110382 291218 145826 291454
rect 146062 291218 146146 291454
rect 146382 291218 162250 291454
rect 162486 291218 192970 291454
rect 193206 291218 217826 291454
rect 218062 291218 218146 291454
rect 218382 291218 253826 291454
rect 254062 291218 254146 291454
rect 254382 291218 264250 291454
rect 264486 291218 294970 291454
rect 295206 291218 325690 291454
rect 325926 291218 356410 291454
rect 356646 291218 387130 291454
rect 387366 291218 417850 291454
rect 418086 291218 448570 291454
rect 448806 291218 479290 291454
rect 479526 291218 510010 291454
rect 510246 291218 540730 291454
rect 540966 291218 577826 291454
rect 578062 291218 578146 291454
rect 578382 291218 585342 291454
rect 585578 291218 585662 291454
rect 585898 291218 592650 291454
rect -8726 291134 592650 291218
rect -8726 290898 -1974 291134
rect -1738 290898 -1654 291134
rect -1418 290898 1826 291134
rect 2062 290898 2146 291134
rect 2382 290898 34250 291134
rect 34486 290898 37826 291134
rect 38062 290898 38146 291134
rect 38382 290898 64970 291134
rect 65206 290898 95690 291134
rect 95926 290898 109826 291134
rect 110062 290898 110146 291134
rect 110382 290898 145826 291134
rect 146062 290898 146146 291134
rect 146382 290898 162250 291134
rect 162486 290898 192970 291134
rect 193206 290898 217826 291134
rect 218062 290898 218146 291134
rect 218382 290898 253826 291134
rect 254062 290898 254146 291134
rect 254382 290898 264250 291134
rect 264486 290898 294970 291134
rect 295206 290898 325690 291134
rect 325926 290898 356410 291134
rect 356646 290898 387130 291134
rect 387366 290898 417850 291134
rect 418086 290898 448570 291134
rect 448806 290898 479290 291134
rect 479526 290898 510010 291134
rect 510246 290898 540730 291134
rect 540966 290898 577826 291134
rect 578062 290898 578146 291134
rect 578382 290898 585342 291134
rect 585578 290898 585662 291134
rect 585898 290898 592650 291134
rect -8726 290866 592650 290898
rect -8726 281494 592650 281526
rect -8726 281258 -8694 281494
rect -8458 281258 -8374 281494
rect -8138 281258 27866 281494
rect 28102 281258 28186 281494
rect 28422 281258 135866 281494
rect 136102 281258 136186 281494
rect 136422 281258 243866 281494
rect 244102 281258 244186 281494
rect 244422 281258 567866 281494
rect 568102 281258 568186 281494
rect 568422 281258 592062 281494
rect 592298 281258 592382 281494
rect 592618 281258 592650 281494
rect -8726 281174 592650 281258
rect -8726 280938 -8694 281174
rect -8458 280938 -8374 281174
rect -8138 280938 27866 281174
rect 28102 280938 28186 281174
rect 28422 280938 135866 281174
rect 136102 280938 136186 281174
rect 136422 280938 243866 281174
rect 244102 280938 244186 281174
rect 244422 280938 567866 281174
rect 568102 280938 568186 281174
rect 568422 280938 592062 281174
rect 592298 280938 592382 281174
rect 592618 280938 592650 281174
rect -8726 280906 592650 280938
rect -8726 277774 592650 277806
rect -8726 277538 -7734 277774
rect -7498 277538 -7414 277774
rect -7178 277538 24146 277774
rect 24382 277538 24466 277774
rect 24702 277538 60146 277774
rect 60382 277538 60466 277774
rect 60702 277538 132146 277774
rect 132382 277538 132466 277774
rect 132702 277538 240146 277774
rect 240382 277538 240466 277774
rect 240702 277538 564146 277774
rect 564382 277538 564466 277774
rect 564702 277538 591102 277774
rect 591338 277538 591422 277774
rect 591658 277538 592650 277774
rect -8726 277454 592650 277538
rect -8726 277218 -7734 277454
rect -7498 277218 -7414 277454
rect -7178 277218 24146 277454
rect 24382 277218 24466 277454
rect 24702 277218 60146 277454
rect 60382 277218 60466 277454
rect 60702 277218 132146 277454
rect 132382 277218 132466 277454
rect 132702 277218 240146 277454
rect 240382 277218 240466 277454
rect 240702 277218 564146 277454
rect 564382 277218 564466 277454
rect 564702 277218 591102 277454
rect 591338 277218 591422 277454
rect 591658 277218 592650 277454
rect -8726 277186 592650 277218
rect -8726 274054 592650 274086
rect -8726 273818 -6774 274054
rect -6538 273818 -6454 274054
rect -6218 273818 20426 274054
rect 20662 273818 20746 274054
rect 20982 273818 56426 274054
rect 56662 273818 56746 274054
rect 56982 273818 128426 274054
rect 128662 273818 128746 274054
rect 128982 273818 236426 274054
rect 236662 273818 236746 274054
rect 236982 273818 560426 274054
rect 560662 273818 560746 274054
rect 560982 273818 590142 274054
rect 590378 273818 590462 274054
rect 590698 273818 592650 274054
rect -8726 273734 592650 273818
rect -8726 273498 -6774 273734
rect -6538 273498 -6454 273734
rect -6218 273498 20426 273734
rect 20662 273498 20746 273734
rect 20982 273498 56426 273734
rect 56662 273498 56746 273734
rect 56982 273498 128426 273734
rect 128662 273498 128746 273734
rect 128982 273498 236426 273734
rect 236662 273498 236746 273734
rect 236982 273498 560426 273734
rect 560662 273498 560746 273734
rect 560982 273498 590142 273734
rect 590378 273498 590462 273734
rect 590698 273498 592650 273734
rect -8726 273466 592650 273498
rect -8726 270334 592650 270366
rect -8726 270098 -5814 270334
rect -5578 270098 -5494 270334
rect -5258 270098 16706 270334
rect 16942 270098 17026 270334
rect 17262 270098 52706 270334
rect 52942 270098 53026 270334
rect 53262 270098 124706 270334
rect 124942 270098 125026 270334
rect 125262 270098 232706 270334
rect 232942 270098 233026 270334
rect 233262 270098 556706 270334
rect 556942 270098 557026 270334
rect 557262 270098 589182 270334
rect 589418 270098 589502 270334
rect 589738 270098 592650 270334
rect -8726 270014 592650 270098
rect -8726 269778 -5814 270014
rect -5578 269778 -5494 270014
rect -5258 269778 16706 270014
rect 16942 269778 17026 270014
rect 17262 269778 52706 270014
rect 52942 269778 53026 270014
rect 53262 269778 124706 270014
rect 124942 269778 125026 270014
rect 125262 269778 232706 270014
rect 232942 269778 233026 270014
rect 233262 269778 556706 270014
rect 556942 269778 557026 270014
rect 557262 269778 589182 270014
rect 589418 269778 589502 270014
rect 589738 269778 592650 270014
rect -8726 269746 592650 269778
rect -8726 266614 592650 266646
rect -8726 266378 -4854 266614
rect -4618 266378 -4534 266614
rect -4298 266378 12986 266614
rect 13222 266378 13306 266614
rect 13542 266378 120986 266614
rect 121222 266378 121306 266614
rect 121542 266378 156986 266614
rect 157222 266378 157306 266614
rect 157542 266378 192986 266614
rect 193222 266378 193306 266614
rect 193542 266378 228986 266614
rect 229222 266378 229306 266614
rect 229542 266378 552986 266614
rect 553222 266378 553306 266614
rect 553542 266378 588222 266614
rect 588458 266378 588542 266614
rect 588778 266378 592650 266614
rect -8726 266294 592650 266378
rect -8726 266058 -4854 266294
rect -4618 266058 -4534 266294
rect -4298 266058 12986 266294
rect 13222 266058 13306 266294
rect 13542 266058 120986 266294
rect 121222 266058 121306 266294
rect 121542 266058 156986 266294
rect 157222 266058 157306 266294
rect 157542 266058 192986 266294
rect 193222 266058 193306 266294
rect 193542 266058 228986 266294
rect 229222 266058 229306 266294
rect 229542 266058 552986 266294
rect 553222 266058 553306 266294
rect 553542 266058 588222 266294
rect 588458 266058 588542 266294
rect 588778 266058 592650 266294
rect -8726 266026 592650 266058
rect -8726 262894 592650 262926
rect -8726 262658 -3894 262894
rect -3658 262658 -3574 262894
rect -3338 262658 9266 262894
rect 9502 262658 9586 262894
rect 9822 262658 45266 262894
rect 45502 262658 45586 262894
rect 45822 262658 117266 262894
rect 117502 262658 117586 262894
rect 117822 262658 153266 262894
rect 153502 262658 153586 262894
rect 153822 262658 189266 262894
rect 189502 262658 189586 262894
rect 189822 262658 225266 262894
rect 225502 262658 225586 262894
rect 225822 262658 587262 262894
rect 587498 262658 587582 262894
rect 587818 262658 592650 262894
rect -8726 262574 592650 262658
rect -8726 262338 -3894 262574
rect -3658 262338 -3574 262574
rect -3338 262338 9266 262574
rect 9502 262338 9586 262574
rect 9822 262338 45266 262574
rect 45502 262338 45586 262574
rect 45822 262338 117266 262574
rect 117502 262338 117586 262574
rect 117822 262338 153266 262574
rect 153502 262338 153586 262574
rect 153822 262338 189266 262574
rect 189502 262338 189586 262574
rect 189822 262338 225266 262574
rect 225502 262338 225586 262574
rect 225822 262338 587262 262574
rect 587498 262338 587582 262574
rect 587818 262338 592650 262574
rect -8726 262306 592650 262338
rect -8726 259174 592650 259206
rect -8726 258938 -2934 259174
rect -2698 258938 -2614 259174
rect -2378 258938 5546 259174
rect 5782 258938 5866 259174
rect 6102 258938 41546 259174
rect 41782 258938 41866 259174
rect 42102 258938 49610 259174
rect 49846 258938 80330 259174
rect 80566 258938 113546 259174
rect 113782 258938 113866 259174
rect 114102 258938 149546 259174
rect 149782 258938 149866 259174
rect 150102 258938 185546 259174
rect 185782 258938 185866 259174
rect 186102 258938 221546 259174
rect 221782 258938 221866 259174
rect 222102 258938 257546 259174
rect 257782 258938 257866 259174
rect 258102 258938 279610 259174
rect 279846 258938 310330 259174
rect 310566 258938 341050 259174
rect 341286 258938 371770 259174
rect 372006 258938 402490 259174
rect 402726 258938 433210 259174
rect 433446 258938 463930 259174
rect 464166 258938 494650 259174
rect 494886 258938 525370 259174
rect 525606 258938 581546 259174
rect 581782 258938 581866 259174
rect 582102 258938 586302 259174
rect 586538 258938 586622 259174
rect 586858 258938 592650 259174
rect -8726 258854 592650 258938
rect -8726 258618 -2934 258854
rect -2698 258618 -2614 258854
rect -2378 258618 5546 258854
rect 5782 258618 5866 258854
rect 6102 258618 41546 258854
rect 41782 258618 41866 258854
rect 42102 258618 49610 258854
rect 49846 258618 80330 258854
rect 80566 258618 113546 258854
rect 113782 258618 113866 258854
rect 114102 258618 149546 258854
rect 149782 258618 149866 258854
rect 150102 258618 185546 258854
rect 185782 258618 185866 258854
rect 186102 258618 221546 258854
rect 221782 258618 221866 258854
rect 222102 258618 257546 258854
rect 257782 258618 257866 258854
rect 258102 258618 279610 258854
rect 279846 258618 310330 258854
rect 310566 258618 341050 258854
rect 341286 258618 371770 258854
rect 372006 258618 402490 258854
rect 402726 258618 433210 258854
rect 433446 258618 463930 258854
rect 464166 258618 494650 258854
rect 494886 258618 525370 258854
rect 525606 258618 581546 258854
rect 581782 258618 581866 258854
rect 582102 258618 586302 258854
rect 586538 258618 586622 258854
rect 586858 258618 592650 258854
rect -8726 258586 592650 258618
rect -8726 255454 592650 255486
rect -8726 255218 -1974 255454
rect -1738 255218 -1654 255454
rect -1418 255218 1826 255454
rect 2062 255218 2146 255454
rect 2382 255218 34250 255454
rect 34486 255218 37826 255454
rect 38062 255218 38146 255454
rect 38382 255218 64970 255454
rect 65206 255218 95690 255454
rect 95926 255218 109826 255454
rect 110062 255218 110146 255454
rect 110382 255218 145826 255454
rect 146062 255218 146146 255454
rect 146382 255218 181826 255454
rect 182062 255218 182146 255454
rect 182382 255218 217826 255454
rect 218062 255218 218146 255454
rect 218382 255218 253826 255454
rect 254062 255218 254146 255454
rect 254382 255218 264250 255454
rect 264486 255218 294970 255454
rect 295206 255218 325690 255454
rect 325926 255218 356410 255454
rect 356646 255218 387130 255454
rect 387366 255218 417850 255454
rect 418086 255218 448570 255454
rect 448806 255218 479290 255454
rect 479526 255218 510010 255454
rect 510246 255218 540730 255454
rect 540966 255218 577826 255454
rect 578062 255218 578146 255454
rect 578382 255218 585342 255454
rect 585578 255218 585662 255454
rect 585898 255218 592650 255454
rect -8726 255134 592650 255218
rect -8726 254898 -1974 255134
rect -1738 254898 -1654 255134
rect -1418 254898 1826 255134
rect 2062 254898 2146 255134
rect 2382 254898 34250 255134
rect 34486 254898 37826 255134
rect 38062 254898 38146 255134
rect 38382 254898 64970 255134
rect 65206 254898 95690 255134
rect 95926 254898 109826 255134
rect 110062 254898 110146 255134
rect 110382 254898 145826 255134
rect 146062 254898 146146 255134
rect 146382 254898 181826 255134
rect 182062 254898 182146 255134
rect 182382 254898 217826 255134
rect 218062 254898 218146 255134
rect 218382 254898 253826 255134
rect 254062 254898 254146 255134
rect 254382 254898 264250 255134
rect 264486 254898 294970 255134
rect 295206 254898 325690 255134
rect 325926 254898 356410 255134
rect 356646 254898 387130 255134
rect 387366 254898 417850 255134
rect 418086 254898 448570 255134
rect 448806 254898 479290 255134
rect 479526 254898 510010 255134
rect 510246 254898 540730 255134
rect 540966 254898 577826 255134
rect 578062 254898 578146 255134
rect 578382 254898 585342 255134
rect 585578 254898 585662 255134
rect 585898 254898 592650 255134
rect -8726 254866 592650 254898
rect -8726 245494 592650 245526
rect -8726 245258 -8694 245494
rect -8458 245258 -8374 245494
rect -8138 245258 27866 245494
rect 28102 245258 28186 245494
rect 28422 245258 135866 245494
rect 136102 245258 136186 245494
rect 136422 245258 171866 245494
rect 172102 245258 172186 245494
rect 172422 245258 207866 245494
rect 208102 245258 208186 245494
rect 208422 245258 243866 245494
rect 244102 245258 244186 245494
rect 244422 245258 567866 245494
rect 568102 245258 568186 245494
rect 568422 245258 592062 245494
rect 592298 245258 592382 245494
rect 592618 245258 592650 245494
rect -8726 245174 592650 245258
rect -8726 244938 -8694 245174
rect -8458 244938 -8374 245174
rect -8138 244938 27866 245174
rect 28102 244938 28186 245174
rect 28422 244938 135866 245174
rect 136102 244938 136186 245174
rect 136422 244938 171866 245174
rect 172102 244938 172186 245174
rect 172422 244938 207866 245174
rect 208102 244938 208186 245174
rect 208422 244938 243866 245174
rect 244102 244938 244186 245174
rect 244422 244938 567866 245174
rect 568102 244938 568186 245174
rect 568422 244938 592062 245174
rect 592298 244938 592382 245174
rect 592618 244938 592650 245174
rect -8726 244906 592650 244938
rect -8726 241774 592650 241806
rect -8726 241538 -7734 241774
rect -7498 241538 -7414 241774
rect -7178 241538 24146 241774
rect 24382 241538 24466 241774
rect 24702 241538 60146 241774
rect 60382 241538 60466 241774
rect 60702 241538 132146 241774
rect 132382 241538 132466 241774
rect 132702 241538 168146 241774
rect 168382 241538 168466 241774
rect 168702 241538 204146 241774
rect 204382 241538 204466 241774
rect 204702 241538 240146 241774
rect 240382 241538 240466 241774
rect 240702 241538 564146 241774
rect 564382 241538 564466 241774
rect 564702 241538 591102 241774
rect 591338 241538 591422 241774
rect 591658 241538 592650 241774
rect -8726 241454 592650 241538
rect -8726 241218 -7734 241454
rect -7498 241218 -7414 241454
rect -7178 241218 24146 241454
rect 24382 241218 24466 241454
rect 24702 241218 60146 241454
rect 60382 241218 60466 241454
rect 60702 241218 132146 241454
rect 132382 241218 132466 241454
rect 132702 241218 168146 241454
rect 168382 241218 168466 241454
rect 168702 241218 204146 241454
rect 204382 241218 204466 241454
rect 204702 241218 240146 241454
rect 240382 241218 240466 241454
rect 240702 241218 564146 241454
rect 564382 241218 564466 241454
rect 564702 241218 591102 241454
rect 591338 241218 591422 241454
rect 591658 241218 592650 241454
rect -8726 241186 592650 241218
rect -8726 238054 592650 238086
rect -8726 237818 -6774 238054
rect -6538 237818 -6454 238054
rect -6218 237818 20426 238054
rect 20662 237818 20746 238054
rect 20982 237818 56426 238054
rect 56662 237818 56746 238054
rect 56982 237818 128426 238054
rect 128662 237818 128746 238054
rect 128982 237818 164426 238054
rect 164662 237818 164746 238054
rect 164982 237818 200426 238054
rect 200662 237818 200746 238054
rect 200982 237818 236426 238054
rect 236662 237818 236746 238054
rect 236982 237818 560426 238054
rect 560662 237818 560746 238054
rect 560982 237818 590142 238054
rect 590378 237818 590462 238054
rect 590698 237818 592650 238054
rect -8726 237734 592650 237818
rect -8726 237498 -6774 237734
rect -6538 237498 -6454 237734
rect -6218 237498 20426 237734
rect 20662 237498 20746 237734
rect 20982 237498 56426 237734
rect 56662 237498 56746 237734
rect 56982 237498 128426 237734
rect 128662 237498 128746 237734
rect 128982 237498 164426 237734
rect 164662 237498 164746 237734
rect 164982 237498 200426 237734
rect 200662 237498 200746 237734
rect 200982 237498 236426 237734
rect 236662 237498 236746 237734
rect 236982 237498 560426 237734
rect 560662 237498 560746 237734
rect 560982 237498 590142 237734
rect 590378 237498 590462 237734
rect 590698 237498 592650 237734
rect -8726 237466 592650 237498
rect -8726 234334 592650 234366
rect -8726 234098 -5814 234334
rect -5578 234098 -5494 234334
rect -5258 234098 16706 234334
rect 16942 234098 17026 234334
rect 17262 234098 52706 234334
rect 52942 234098 53026 234334
rect 53262 234098 124706 234334
rect 124942 234098 125026 234334
rect 125262 234098 160706 234334
rect 160942 234098 161026 234334
rect 161262 234098 196706 234334
rect 196942 234098 197026 234334
rect 197262 234098 232706 234334
rect 232942 234098 233026 234334
rect 233262 234098 556706 234334
rect 556942 234098 557026 234334
rect 557262 234098 589182 234334
rect 589418 234098 589502 234334
rect 589738 234098 592650 234334
rect -8726 234014 592650 234098
rect -8726 233778 -5814 234014
rect -5578 233778 -5494 234014
rect -5258 233778 16706 234014
rect 16942 233778 17026 234014
rect 17262 233778 52706 234014
rect 52942 233778 53026 234014
rect 53262 233778 124706 234014
rect 124942 233778 125026 234014
rect 125262 233778 160706 234014
rect 160942 233778 161026 234014
rect 161262 233778 196706 234014
rect 196942 233778 197026 234014
rect 197262 233778 232706 234014
rect 232942 233778 233026 234014
rect 233262 233778 556706 234014
rect 556942 233778 557026 234014
rect 557262 233778 589182 234014
rect 589418 233778 589502 234014
rect 589738 233778 592650 234014
rect -8726 233746 592650 233778
rect -8726 230614 592650 230646
rect -8726 230378 -4854 230614
rect -4618 230378 -4534 230614
rect -4298 230378 12986 230614
rect 13222 230378 13306 230614
rect 13542 230378 120986 230614
rect 121222 230378 121306 230614
rect 121542 230378 156986 230614
rect 157222 230378 157306 230614
rect 157542 230378 192986 230614
rect 193222 230378 193306 230614
rect 193542 230378 228986 230614
rect 229222 230378 229306 230614
rect 229542 230378 552986 230614
rect 553222 230378 553306 230614
rect 553542 230378 588222 230614
rect 588458 230378 588542 230614
rect 588778 230378 592650 230614
rect -8726 230294 592650 230378
rect -8726 230058 -4854 230294
rect -4618 230058 -4534 230294
rect -4298 230058 12986 230294
rect 13222 230058 13306 230294
rect 13542 230058 120986 230294
rect 121222 230058 121306 230294
rect 121542 230058 156986 230294
rect 157222 230058 157306 230294
rect 157542 230058 192986 230294
rect 193222 230058 193306 230294
rect 193542 230058 228986 230294
rect 229222 230058 229306 230294
rect 229542 230058 552986 230294
rect 553222 230058 553306 230294
rect 553542 230058 588222 230294
rect 588458 230058 588542 230294
rect 588778 230058 592650 230294
rect -8726 230026 592650 230058
rect -8726 226894 592650 226926
rect -8726 226658 -3894 226894
rect -3658 226658 -3574 226894
rect -3338 226658 9266 226894
rect 9502 226658 9586 226894
rect 9822 226658 45266 226894
rect 45502 226658 45586 226894
rect 45822 226658 117266 226894
rect 117502 226658 117586 226894
rect 117822 226658 153266 226894
rect 153502 226658 153586 226894
rect 153822 226658 189266 226894
rect 189502 226658 189586 226894
rect 189822 226658 225266 226894
rect 225502 226658 225586 226894
rect 225822 226658 587262 226894
rect 587498 226658 587582 226894
rect 587818 226658 592650 226894
rect -8726 226574 592650 226658
rect -8726 226338 -3894 226574
rect -3658 226338 -3574 226574
rect -3338 226338 9266 226574
rect 9502 226338 9586 226574
rect 9822 226338 45266 226574
rect 45502 226338 45586 226574
rect 45822 226338 117266 226574
rect 117502 226338 117586 226574
rect 117822 226338 153266 226574
rect 153502 226338 153586 226574
rect 153822 226338 189266 226574
rect 189502 226338 189586 226574
rect 189822 226338 225266 226574
rect 225502 226338 225586 226574
rect 225822 226338 587262 226574
rect 587498 226338 587582 226574
rect 587818 226338 592650 226574
rect -8726 226306 592650 226338
rect -8726 223174 592650 223206
rect -8726 222938 -2934 223174
rect -2698 222938 -2614 223174
rect -2378 222938 5546 223174
rect 5782 222938 5866 223174
rect 6102 222938 41546 223174
rect 41782 222938 41866 223174
rect 42102 222938 49610 223174
rect 49846 222938 80330 223174
rect 80566 222938 113546 223174
rect 113782 222938 113866 223174
rect 114102 222938 149546 223174
rect 149782 222938 149866 223174
rect 150102 222938 185546 223174
rect 185782 222938 185866 223174
rect 186102 222938 221546 223174
rect 221782 222938 221866 223174
rect 222102 222938 257546 223174
rect 257782 222938 257866 223174
rect 258102 222938 279610 223174
rect 279846 222938 310330 223174
rect 310566 222938 341050 223174
rect 341286 222938 371770 223174
rect 372006 222938 402490 223174
rect 402726 222938 433210 223174
rect 433446 222938 463930 223174
rect 464166 222938 494650 223174
rect 494886 222938 525370 223174
rect 525606 222938 581546 223174
rect 581782 222938 581866 223174
rect 582102 222938 586302 223174
rect 586538 222938 586622 223174
rect 586858 222938 592650 223174
rect -8726 222854 592650 222938
rect -8726 222618 -2934 222854
rect -2698 222618 -2614 222854
rect -2378 222618 5546 222854
rect 5782 222618 5866 222854
rect 6102 222618 41546 222854
rect 41782 222618 41866 222854
rect 42102 222618 49610 222854
rect 49846 222618 80330 222854
rect 80566 222618 113546 222854
rect 113782 222618 113866 222854
rect 114102 222618 149546 222854
rect 149782 222618 149866 222854
rect 150102 222618 185546 222854
rect 185782 222618 185866 222854
rect 186102 222618 221546 222854
rect 221782 222618 221866 222854
rect 222102 222618 257546 222854
rect 257782 222618 257866 222854
rect 258102 222618 279610 222854
rect 279846 222618 310330 222854
rect 310566 222618 341050 222854
rect 341286 222618 371770 222854
rect 372006 222618 402490 222854
rect 402726 222618 433210 222854
rect 433446 222618 463930 222854
rect 464166 222618 494650 222854
rect 494886 222618 525370 222854
rect 525606 222618 581546 222854
rect 581782 222618 581866 222854
rect 582102 222618 586302 222854
rect 586538 222618 586622 222854
rect 586858 222618 592650 222854
rect -8726 222586 592650 222618
rect -8726 219454 592650 219486
rect -8726 219218 -1974 219454
rect -1738 219218 -1654 219454
rect -1418 219218 1826 219454
rect 2062 219218 2146 219454
rect 2382 219218 34250 219454
rect 34486 219218 37826 219454
rect 38062 219218 38146 219454
rect 38382 219218 64970 219454
rect 65206 219218 95690 219454
rect 95926 219218 109826 219454
rect 110062 219218 110146 219454
rect 110382 219218 145826 219454
rect 146062 219218 146146 219454
rect 146382 219218 181826 219454
rect 182062 219218 182146 219454
rect 182382 219218 217826 219454
rect 218062 219218 218146 219454
rect 218382 219218 253826 219454
rect 254062 219218 254146 219454
rect 254382 219218 264250 219454
rect 264486 219218 294970 219454
rect 295206 219218 325690 219454
rect 325926 219218 356410 219454
rect 356646 219218 387130 219454
rect 387366 219218 417850 219454
rect 418086 219218 448570 219454
rect 448806 219218 479290 219454
rect 479526 219218 510010 219454
rect 510246 219218 540730 219454
rect 540966 219218 577826 219454
rect 578062 219218 578146 219454
rect 578382 219218 585342 219454
rect 585578 219218 585662 219454
rect 585898 219218 592650 219454
rect -8726 219134 592650 219218
rect -8726 218898 -1974 219134
rect -1738 218898 -1654 219134
rect -1418 218898 1826 219134
rect 2062 218898 2146 219134
rect 2382 218898 34250 219134
rect 34486 218898 37826 219134
rect 38062 218898 38146 219134
rect 38382 218898 64970 219134
rect 65206 218898 95690 219134
rect 95926 218898 109826 219134
rect 110062 218898 110146 219134
rect 110382 218898 145826 219134
rect 146062 218898 146146 219134
rect 146382 218898 181826 219134
rect 182062 218898 182146 219134
rect 182382 218898 217826 219134
rect 218062 218898 218146 219134
rect 218382 218898 253826 219134
rect 254062 218898 254146 219134
rect 254382 218898 264250 219134
rect 264486 218898 294970 219134
rect 295206 218898 325690 219134
rect 325926 218898 356410 219134
rect 356646 218898 387130 219134
rect 387366 218898 417850 219134
rect 418086 218898 448570 219134
rect 448806 218898 479290 219134
rect 479526 218898 510010 219134
rect 510246 218898 540730 219134
rect 540966 218898 577826 219134
rect 578062 218898 578146 219134
rect 578382 218898 585342 219134
rect 585578 218898 585662 219134
rect 585898 218898 592650 219134
rect -8726 218866 592650 218898
rect -8726 209494 592650 209526
rect -8726 209258 -8694 209494
rect -8458 209258 -8374 209494
rect -8138 209258 27866 209494
rect 28102 209258 28186 209494
rect 28422 209258 135866 209494
rect 136102 209258 136186 209494
rect 136422 209258 171866 209494
rect 172102 209258 172186 209494
rect 172422 209258 207866 209494
rect 208102 209258 208186 209494
rect 208422 209258 243866 209494
rect 244102 209258 244186 209494
rect 244422 209258 567866 209494
rect 568102 209258 568186 209494
rect 568422 209258 592062 209494
rect 592298 209258 592382 209494
rect 592618 209258 592650 209494
rect -8726 209174 592650 209258
rect -8726 208938 -8694 209174
rect -8458 208938 -8374 209174
rect -8138 208938 27866 209174
rect 28102 208938 28186 209174
rect 28422 208938 135866 209174
rect 136102 208938 136186 209174
rect 136422 208938 171866 209174
rect 172102 208938 172186 209174
rect 172422 208938 207866 209174
rect 208102 208938 208186 209174
rect 208422 208938 243866 209174
rect 244102 208938 244186 209174
rect 244422 208938 567866 209174
rect 568102 208938 568186 209174
rect 568422 208938 592062 209174
rect 592298 208938 592382 209174
rect 592618 208938 592650 209174
rect -8726 208906 592650 208938
rect -8726 205774 592650 205806
rect -8726 205538 -7734 205774
rect -7498 205538 -7414 205774
rect -7178 205538 24146 205774
rect 24382 205538 24466 205774
rect 24702 205538 60146 205774
rect 60382 205538 60466 205774
rect 60702 205538 132146 205774
rect 132382 205538 132466 205774
rect 132702 205538 168146 205774
rect 168382 205538 168466 205774
rect 168702 205538 204146 205774
rect 204382 205538 204466 205774
rect 204702 205538 240146 205774
rect 240382 205538 240466 205774
rect 240702 205538 564146 205774
rect 564382 205538 564466 205774
rect 564702 205538 591102 205774
rect 591338 205538 591422 205774
rect 591658 205538 592650 205774
rect -8726 205454 592650 205538
rect -8726 205218 -7734 205454
rect -7498 205218 -7414 205454
rect -7178 205218 24146 205454
rect 24382 205218 24466 205454
rect 24702 205218 60146 205454
rect 60382 205218 60466 205454
rect 60702 205218 132146 205454
rect 132382 205218 132466 205454
rect 132702 205218 168146 205454
rect 168382 205218 168466 205454
rect 168702 205218 204146 205454
rect 204382 205218 204466 205454
rect 204702 205218 240146 205454
rect 240382 205218 240466 205454
rect 240702 205218 564146 205454
rect 564382 205218 564466 205454
rect 564702 205218 591102 205454
rect 591338 205218 591422 205454
rect 591658 205218 592650 205454
rect -8726 205186 592650 205218
rect -8726 202054 592650 202086
rect -8726 201818 -6774 202054
rect -6538 201818 -6454 202054
rect -6218 201818 20426 202054
rect 20662 201818 20746 202054
rect 20982 201818 56426 202054
rect 56662 201818 56746 202054
rect 56982 201818 128426 202054
rect 128662 201818 128746 202054
rect 128982 201818 164426 202054
rect 164662 201818 164746 202054
rect 164982 201818 200426 202054
rect 200662 201818 200746 202054
rect 200982 201818 236426 202054
rect 236662 201818 236746 202054
rect 236982 201818 560426 202054
rect 560662 201818 560746 202054
rect 560982 201818 590142 202054
rect 590378 201818 590462 202054
rect 590698 201818 592650 202054
rect -8726 201734 592650 201818
rect -8726 201498 -6774 201734
rect -6538 201498 -6454 201734
rect -6218 201498 20426 201734
rect 20662 201498 20746 201734
rect 20982 201498 56426 201734
rect 56662 201498 56746 201734
rect 56982 201498 128426 201734
rect 128662 201498 128746 201734
rect 128982 201498 164426 201734
rect 164662 201498 164746 201734
rect 164982 201498 200426 201734
rect 200662 201498 200746 201734
rect 200982 201498 236426 201734
rect 236662 201498 236746 201734
rect 236982 201498 560426 201734
rect 560662 201498 560746 201734
rect 560982 201498 590142 201734
rect 590378 201498 590462 201734
rect 590698 201498 592650 201734
rect -8726 201466 592650 201498
rect -8726 198334 592650 198366
rect -8726 198098 -5814 198334
rect -5578 198098 -5494 198334
rect -5258 198098 16706 198334
rect 16942 198098 17026 198334
rect 17262 198098 52706 198334
rect 52942 198098 53026 198334
rect 53262 198098 124706 198334
rect 124942 198098 125026 198334
rect 125262 198098 160706 198334
rect 160942 198098 161026 198334
rect 161262 198098 196706 198334
rect 196942 198098 197026 198334
rect 197262 198098 232706 198334
rect 232942 198098 233026 198334
rect 233262 198098 556706 198334
rect 556942 198098 557026 198334
rect 557262 198098 589182 198334
rect 589418 198098 589502 198334
rect 589738 198098 592650 198334
rect -8726 198014 592650 198098
rect -8726 197778 -5814 198014
rect -5578 197778 -5494 198014
rect -5258 197778 16706 198014
rect 16942 197778 17026 198014
rect 17262 197778 52706 198014
rect 52942 197778 53026 198014
rect 53262 197778 124706 198014
rect 124942 197778 125026 198014
rect 125262 197778 160706 198014
rect 160942 197778 161026 198014
rect 161262 197778 196706 198014
rect 196942 197778 197026 198014
rect 197262 197778 232706 198014
rect 232942 197778 233026 198014
rect 233262 197778 556706 198014
rect 556942 197778 557026 198014
rect 557262 197778 589182 198014
rect 589418 197778 589502 198014
rect 589738 197778 592650 198014
rect -8726 197746 592650 197778
rect -8726 194614 592650 194646
rect -8726 194378 -4854 194614
rect -4618 194378 -4534 194614
rect -4298 194378 12986 194614
rect 13222 194378 13306 194614
rect 13542 194378 120986 194614
rect 121222 194378 121306 194614
rect 121542 194378 156986 194614
rect 157222 194378 157306 194614
rect 157542 194378 192986 194614
rect 193222 194378 193306 194614
rect 193542 194378 228986 194614
rect 229222 194378 229306 194614
rect 229542 194378 552986 194614
rect 553222 194378 553306 194614
rect 553542 194378 588222 194614
rect 588458 194378 588542 194614
rect 588778 194378 592650 194614
rect -8726 194294 592650 194378
rect -8726 194058 -4854 194294
rect -4618 194058 -4534 194294
rect -4298 194058 12986 194294
rect 13222 194058 13306 194294
rect 13542 194058 120986 194294
rect 121222 194058 121306 194294
rect 121542 194058 156986 194294
rect 157222 194058 157306 194294
rect 157542 194058 192986 194294
rect 193222 194058 193306 194294
rect 193542 194058 228986 194294
rect 229222 194058 229306 194294
rect 229542 194058 552986 194294
rect 553222 194058 553306 194294
rect 553542 194058 588222 194294
rect 588458 194058 588542 194294
rect 588778 194058 592650 194294
rect -8726 194026 592650 194058
rect -8726 190894 592650 190926
rect -8726 190658 -3894 190894
rect -3658 190658 -3574 190894
rect -3338 190658 9266 190894
rect 9502 190658 9586 190894
rect 9822 190658 45266 190894
rect 45502 190658 45586 190894
rect 45822 190658 117266 190894
rect 117502 190658 117586 190894
rect 117822 190658 153266 190894
rect 153502 190658 153586 190894
rect 153822 190658 189266 190894
rect 189502 190658 189586 190894
rect 189822 190658 225266 190894
rect 225502 190658 225586 190894
rect 225822 190658 587262 190894
rect 587498 190658 587582 190894
rect 587818 190658 592650 190894
rect -8726 190574 592650 190658
rect -8726 190338 -3894 190574
rect -3658 190338 -3574 190574
rect -3338 190338 9266 190574
rect 9502 190338 9586 190574
rect 9822 190338 45266 190574
rect 45502 190338 45586 190574
rect 45822 190338 117266 190574
rect 117502 190338 117586 190574
rect 117822 190338 153266 190574
rect 153502 190338 153586 190574
rect 153822 190338 189266 190574
rect 189502 190338 189586 190574
rect 189822 190338 225266 190574
rect 225502 190338 225586 190574
rect 225822 190338 587262 190574
rect 587498 190338 587582 190574
rect 587818 190338 592650 190574
rect -8726 190306 592650 190338
rect -8726 187174 592650 187206
rect -8726 186938 -2934 187174
rect -2698 186938 -2614 187174
rect -2378 186938 5546 187174
rect 5782 186938 5866 187174
rect 6102 186938 41546 187174
rect 41782 186938 41866 187174
rect 42102 186938 49610 187174
rect 49846 186938 80330 187174
rect 80566 186938 113546 187174
rect 113782 186938 113866 187174
rect 114102 186938 149546 187174
rect 149782 186938 149866 187174
rect 150102 186938 185546 187174
rect 185782 186938 185866 187174
rect 186102 186938 221546 187174
rect 221782 186938 221866 187174
rect 222102 186938 257546 187174
rect 257782 186938 257866 187174
rect 258102 186938 279610 187174
rect 279846 186938 310330 187174
rect 310566 186938 341050 187174
rect 341286 186938 371770 187174
rect 372006 186938 402490 187174
rect 402726 186938 433210 187174
rect 433446 186938 463930 187174
rect 464166 186938 494650 187174
rect 494886 186938 525370 187174
rect 525606 186938 581546 187174
rect 581782 186938 581866 187174
rect 582102 186938 586302 187174
rect 586538 186938 586622 187174
rect 586858 186938 592650 187174
rect -8726 186854 592650 186938
rect -8726 186618 -2934 186854
rect -2698 186618 -2614 186854
rect -2378 186618 5546 186854
rect 5782 186618 5866 186854
rect 6102 186618 41546 186854
rect 41782 186618 41866 186854
rect 42102 186618 49610 186854
rect 49846 186618 80330 186854
rect 80566 186618 113546 186854
rect 113782 186618 113866 186854
rect 114102 186618 149546 186854
rect 149782 186618 149866 186854
rect 150102 186618 185546 186854
rect 185782 186618 185866 186854
rect 186102 186618 221546 186854
rect 221782 186618 221866 186854
rect 222102 186618 257546 186854
rect 257782 186618 257866 186854
rect 258102 186618 279610 186854
rect 279846 186618 310330 186854
rect 310566 186618 341050 186854
rect 341286 186618 371770 186854
rect 372006 186618 402490 186854
rect 402726 186618 433210 186854
rect 433446 186618 463930 186854
rect 464166 186618 494650 186854
rect 494886 186618 525370 186854
rect 525606 186618 581546 186854
rect 581782 186618 581866 186854
rect 582102 186618 586302 186854
rect 586538 186618 586622 186854
rect 586858 186618 592650 186854
rect -8726 186586 592650 186618
rect -8726 183454 592650 183486
rect -8726 183218 -1974 183454
rect -1738 183218 -1654 183454
rect -1418 183218 1826 183454
rect 2062 183218 2146 183454
rect 2382 183218 34250 183454
rect 34486 183218 37826 183454
rect 38062 183218 38146 183454
rect 38382 183218 64970 183454
rect 65206 183218 95690 183454
rect 95926 183218 109826 183454
rect 110062 183218 110146 183454
rect 110382 183218 145826 183454
rect 146062 183218 146146 183454
rect 146382 183218 181826 183454
rect 182062 183218 182146 183454
rect 182382 183218 217826 183454
rect 218062 183218 218146 183454
rect 218382 183218 253826 183454
rect 254062 183218 254146 183454
rect 254382 183218 264250 183454
rect 264486 183218 294970 183454
rect 295206 183218 325690 183454
rect 325926 183218 356410 183454
rect 356646 183218 387130 183454
rect 387366 183218 417850 183454
rect 418086 183218 448570 183454
rect 448806 183218 479290 183454
rect 479526 183218 510010 183454
rect 510246 183218 540730 183454
rect 540966 183218 577826 183454
rect 578062 183218 578146 183454
rect 578382 183218 585342 183454
rect 585578 183218 585662 183454
rect 585898 183218 592650 183454
rect -8726 183134 592650 183218
rect -8726 182898 -1974 183134
rect -1738 182898 -1654 183134
rect -1418 182898 1826 183134
rect 2062 182898 2146 183134
rect 2382 182898 34250 183134
rect 34486 182898 37826 183134
rect 38062 182898 38146 183134
rect 38382 182898 64970 183134
rect 65206 182898 95690 183134
rect 95926 182898 109826 183134
rect 110062 182898 110146 183134
rect 110382 182898 145826 183134
rect 146062 182898 146146 183134
rect 146382 182898 181826 183134
rect 182062 182898 182146 183134
rect 182382 182898 217826 183134
rect 218062 182898 218146 183134
rect 218382 182898 253826 183134
rect 254062 182898 254146 183134
rect 254382 182898 264250 183134
rect 264486 182898 294970 183134
rect 295206 182898 325690 183134
rect 325926 182898 356410 183134
rect 356646 182898 387130 183134
rect 387366 182898 417850 183134
rect 418086 182898 448570 183134
rect 448806 182898 479290 183134
rect 479526 182898 510010 183134
rect 510246 182898 540730 183134
rect 540966 182898 577826 183134
rect 578062 182898 578146 183134
rect 578382 182898 585342 183134
rect 585578 182898 585662 183134
rect 585898 182898 592650 183134
rect -8726 182866 592650 182898
rect -8726 173494 592650 173526
rect -8726 173258 -8694 173494
rect -8458 173258 -8374 173494
rect -8138 173258 27866 173494
rect 28102 173258 28186 173494
rect 28422 173258 135866 173494
rect 136102 173258 136186 173494
rect 136422 173258 171866 173494
rect 172102 173258 172186 173494
rect 172422 173258 207866 173494
rect 208102 173258 208186 173494
rect 208422 173258 243866 173494
rect 244102 173258 244186 173494
rect 244422 173258 567866 173494
rect 568102 173258 568186 173494
rect 568422 173258 592062 173494
rect 592298 173258 592382 173494
rect 592618 173258 592650 173494
rect -8726 173174 592650 173258
rect -8726 172938 -8694 173174
rect -8458 172938 -8374 173174
rect -8138 172938 27866 173174
rect 28102 172938 28186 173174
rect 28422 172938 135866 173174
rect 136102 172938 136186 173174
rect 136422 172938 171866 173174
rect 172102 172938 172186 173174
rect 172422 172938 207866 173174
rect 208102 172938 208186 173174
rect 208422 172938 243866 173174
rect 244102 172938 244186 173174
rect 244422 172938 567866 173174
rect 568102 172938 568186 173174
rect 568422 172938 592062 173174
rect 592298 172938 592382 173174
rect 592618 172938 592650 173174
rect -8726 172906 592650 172938
rect -8726 169774 592650 169806
rect -8726 169538 -7734 169774
rect -7498 169538 -7414 169774
rect -7178 169538 24146 169774
rect 24382 169538 24466 169774
rect 24702 169538 60146 169774
rect 60382 169538 60466 169774
rect 60702 169538 132146 169774
rect 132382 169538 132466 169774
rect 132702 169538 168146 169774
rect 168382 169538 168466 169774
rect 168702 169538 204146 169774
rect 204382 169538 204466 169774
rect 204702 169538 240146 169774
rect 240382 169538 240466 169774
rect 240702 169538 564146 169774
rect 564382 169538 564466 169774
rect 564702 169538 591102 169774
rect 591338 169538 591422 169774
rect 591658 169538 592650 169774
rect -8726 169454 592650 169538
rect -8726 169218 -7734 169454
rect -7498 169218 -7414 169454
rect -7178 169218 24146 169454
rect 24382 169218 24466 169454
rect 24702 169218 60146 169454
rect 60382 169218 60466 169454
rect 60702 169218 132146 169454
rect 132382 169218 132466 169454
rect 132702 169218 168146 169454
rect 168382 169218 168466 169454
rect 168702 169218 204146 169454
rect 204382 169218 204466 169454
rect 204702 169218 240146 169454
rect 240382 169218 240466 169454
rect 240702 169218 564146 169454
rect 564382 169218 564466 169454
rect 564702 169218 591102 169454
rect 591338 169218 591422 169454
rect 591658 169218 592650 169454
rect -8726 169186 592650 169218
rect -8726 166054 592650 166086
rect -8726 165818 -6774 166054
rect -6538 165818 -6454 166054
rect -6218 165818 20426 166054
rect 20662 165818 20746 166054
rect 20982 165818 56426 166054
rect 56662 165818 56746 166054
rect 56982 165818 92426 166054
rect 92662 165818 92746 166054
rect 92982 165818 128426 166054
rect 128662 165818 128746 166054
rect 128982 165818 164426 166054
rect 164662 165818 164746 166054
rect 164982 165818 200426 166054
rect 200662 165818 200746 166054
rect 200982 165818 236426 166054
rect 236662 165818 236746 166054
rect 236982 165818 560426 166054
rect 560662 165818 560746 166054
rect 560982 165818 590142 166054
rect 590378 165818 590462 166054
rect 590698 165818 592650 166054
rect -8726 165734 592650 165818
rect -8726 165498 -6774 165734
rect -6538 165498 -6454 165734
rect -6218 165498 20426 165734
rect 20662 165498 20746 165734
rect 20982 165498 56426 165734
rect 56662 165498 56746 165734
rect 56982 165498 92426 165734
rect 92662 165498 92746 165734
rect 92982 165498 128426 165734
rect 128662 165498 128746 165734
rect 128982 165498 164426 165734
rect 164662 165498 164746 165734
rect 164982 165498 200426 165734
rect 200662 165498 200746 165734
rect 200982 165498 236426 165734
rect 236662 165498 236746 165734
rect 236982 165498 560426 165734
rect 560662 165498 560746 165734
rect 560982 165498 590142 165734
rect 590378 165498 590462 165734
rect 590698 165498 592650 165734
rect -8726 165466 592650 165498
rect -8726 162334 592650 162366
rect -8726 162098 -5814 162334
rect -5578 162098 -5494 162334
rect -5258 162098 16706 162334
rect 16942 162098 17026 162334
rect 17262 162098 52706 162334
rect 52942 162098 53026 162334
rect 53262 162098 88706 162334
rect 88942 162098 89026 162334
rect 89262 162098 124706 162334
rect 124942 162098 125026 162334
rect 125262 162098 160706 162334
rect 160942 162098 161026 162334
rect 161262 162098 196706 162334
rect 196942 162098 197026 162334
rect 197262 162098 232706 162334
rect 232942 162098 233026 162334
rect 233262 162098 556706 162334
rect 556942 162098 557026 162334
rect 557262 162098 589182 162334
rect 589418 162098 589502 162334
rect 589738 162098 592650 162334
rect -8726 162014 592650 162098
rect -8726 161778 -5814 162014
rect -5578 161778 -5494 162014
rect -5258 161778 16706 162014
rect 16942 161778 17026 162014
rect 17262 161778 52706 162014
rect 52942 161778 53026 162014
rect 53262 161778 88706 162014
rect 88942 161778 89026 162014
rect 89262 161778 124706 162014
rect 124942 161778 125026 162014
rect 125262 161778 160706 162014
rect 160942 161778 161026 162014
rect 161262 161778 196706 162014
rect 196942 161778 197026 162014
rect 197262 161778 232706 162014
rect 232942 161778 233026 162014
rect 233262 161778 556706 162014
rect 556942 161778 557026 162014
rect 557262 161778 589182 162014
rect 589418 161778 589502 162014
rect 589738 161778 592650 162014
rect -8726 161746 592650 161778
rect -8726 158614 592650 158646
rect -8726 158378 -4854 158614
rect -4618 158378 -4534 158614
rect -4298 158378 12986 158614
rect 13222 158378 13306 158614
rect 13542 158378 120986 158614
rect 121222 158378 121306 158614
rect 121542 158378 156986 158614
rect 157222 158378 157306 158614
rect 157542 158378 192986 158614
rect 193222 158378 193306 158614
rect 193542 158378 228986 158614
rect 229222 158378 229306 158614
rect 229542 158378 552986 158614
rect 553222 158378 553306 158614
rect 553542 158378 588222 158614
rect 588458 158378 588542 158614
rect 588778 158378 592650 158614
rect -8726 158294 592650 158378
rect -8726 158058 -4854 158294
rect -4618 158058 -4534 158294
rect -4298 158058 12986 158294
rect 13222 158058 13306 158294
rect 13542 158058 120986 158294
rect 121222 158058 121306 158294
rect 121542 158058 156986 158294
rect 157222 158058 157306 158294
rect 157542 158058 192986 158294
rect 193222 158058 193306 158294
rect 193542 158058 228986 158294
rect 229222 158058 229306 158294
rect 229542 158058 552986 158294
rect 553222 158058 553306 158294
rect 553542 158058 588222 158294
rect 588458 158058 588542 158294
rect 588778 158058 592650 158294
rect -8726 158026 592650 158058
rect -8726 154894 592650 154926
rect -8726 154658 -3894 154894
rect -3658 154658 -3574 154894
rect -3338 154658 9266 154894
rect 9502 154658 9586 154894
rect 9822 154658 45266 154894
rect 45502 154658 45586 154894
rect 45822 154658 117266 154894
rect 117502 154658 117586 154894
rect 117822 154658 153266 154894
rect 153502 154658 153586 154894
rect 153822 154658 189266 154894
rect 189502 154658 189586 154894
rect 189822 154658 225266 154894
rect 225502 154658 225586 154894
rect 225822 154658 587262 154894
rect 587498 154658 587582 154894
rect 587818 154658 592650 154894
rect -8726 154574 592650 154658
rect -8726 154338 -3894 154574
rect -3658 154338 -3574 154574
rect -3338 154338 9266 154574
rect 9502 154338 9586 154574
rect 9822 154338 45266 154574
rect 45502 154338 45586 154574
rect 45822 154338 117266 154574
rect 117502 154338 117586 154574
rect 117822 154338 153266 154574
rect 153502 154338 153586 154574
rect 153822 154338 189266 154574
rect 189502 154338 189586 154574
rect 189822 154338 225266 154574
rect 225502 154338 225586 154574
rect 225822 154338 587262 154574
rect 587498 154338 587582 154574
rect 587818 154338 592650 154574
rect -8726 154306 592650 154338
rect -8726 151174 592650 151206
rect -8726 150938 -2934 151174
rect -2698 150938 -2614 151174
rect -2378 150938 5546 151174
rect 5782 150938 5866 151174
rect 6102 150938 41546 151174
rect 41782 150938 41866 151174
rect 42102 150938 113546 151174
rect 113782 150938 113866 151174
rect 114102 150938 149546 151174
rect 149782 150938 149866 151174
rect 150102 150938 185546 151174
rect 185782 150938 185866 151174
rect 186102 150938 221546 151174
rect 221782 150938 221866 151174
rect 222102 150938 257546 151174
rect 257782 150938 257866 151174
rect 258102 150938 279610 151174
rect 279846 150938 310330 151174
rect 310566 150938 341050 151174
rect 341286 150938 371770 151174
rect 372006 150938 402490 151174
rect 402726 150938 433210 151174
rect 433446 150938 463930 151174
rect 464166 150938 494650 151174
rect 494886 150938 525370 151174
rect 525606 150938 581546 151174
rect 581782 150938 581866 151174
rect 582102 150938 586302 151174
rect 586538 150938 586622 151174
rect 586858 150938 592650 151174
rect -8726 150854 592650 150938
rect -8726 150618 -2934 150854
rect -2698 150618 -2614 150854
rect -2378 150618 5546 150854
rect 5782 150618 5866 150854
rect 6102 150618 41546 150854
rect 41782 150618 41866 150854
rect 42102 150618 113546 150854
rect 113782 150618 113866 150854
rect 114102 150618 149546 150854
rect 149782 150618 149866 150854
rect 150102 150618 185546 150854
rect 185782 150618 185866 150854
rect 186102 150618 221546 150854
rect 221782 150618 221866 150854
rect 222102 150618 257546 150854
rect 257782 150618 257866 150854
rect 258102 150618 279610 150854
rect 279846 150618 310330 150854
rect 310566 150618 341050 150854
rect 341286 150618 371770 150854
rect 372006 150618 402490 150854
rect 402726 150618 433210 150854
rect 433446 150618 463930 150854
rect 464166 150618 494650 150854
rect 494886 150618 525370 150854
rect 525606 150618 581546 150854
rect 581782 150618 581866 150854
rect 582102 150618 586302 150854
rect 586538 150618 586622 150854
rect 586858 150618 592650 150854
rect -8726 150586 592650 150618
rect -8726 147454 592650 147486
rect -8726 147218 -1974 147454
rect -1738 147218 -1654 147454
rect -1418 147218 1826 147454
rect 2062 147218 2146 147454
rect 2382 147218 37826 147454
rect 38062 147218 38146 147454
rect 38382 147218 109826 147454
rect 110062 147218 110146 147454
rect 110382 147218 145826 147454
rect 146062 147218 146146 147454
rect 146382 147218 181826 147454
rect 182062 147218 182146 147454
rect 182382 147218 217826 147454
rect 218062 147218 218146 147454
rect 218382 147218 253826 147454
rect 254062 147218 254146 147454
rect 254382 147218 264250 147454
rect 264486 147218 294970 147454
rect 295206 147218 325690 147454
rect 325926 147218 356410 147454
rect 356646 147218 387130 147454
rect 387366 147218 417850 147454
rect 418086 147218 448570 147454
rect 448806 147218 479290 147454
rect 479526 147218 510010 147454
rect 510246 147218 540730 147454
rect 540966 147218 577826 147454
rect 578062 147218 578146 147454
rect 578382 147218 585342 147454
rect 585578 147218 585662 147454
rect 585898 147218 592650 147454
rect -8726 147134 592650 147218
rect -8726 146898 -1974 147134
rect -1738 146898 -1654 147134
rect -1418 146898 1826 147134
rect 2062 146898 2146 147134
rect 2382 146898 37826 147134
rect 38062 146898 38146 147134
rect 38382 146898 109826 147134
rect 110062 146898 110146 147134
rect 110382 146898 145826 147134
rect 146062 146898 146146 147134
rect 146382 146898 181826 147134
rect 182062 146898 182146 147134
rect 182382 146898 217826 147134
rect 218062 146898 218146 147134
rect 218382 146898 253826 147134
rect 254062 146898 254146 147134
rect 254382 146898 264250 147134
rect 264486 146898 294970 147134
rect 295206 146898 325690 147134
rect 325926 146898 356410 147134
rect 356646 146898 387130 147134
rect 387366 146898 417850 147134
rect 418086 146898 448570 147134
rect 448806 146898 479290 147134
rect 479526 146898 510010 147134
rect 510246 146898 540730 147134
rect 540966 146898 577826 147134
rect 578062 146898 578146 147134
rect 578382 146898 585342 147134
rect 585578 146898 585662 147134
rect 585898 146898 592650 147134
rect -8726 146866 592650 146898
rect -8726 137494 592650 137526
rect -8726 137258 -8694 137494
rect -8458 137258 -8374 137494
rect -8138 137258 27866 137494
rect 28102 137258 28186 137494
rect 28422 137258 135866 137494
rect 136102 137258 136186 137494
rect 136422 137258 171866 137494
rect 172102 137258 172186 137494
rect 172422 137258 207866 137494
rect 208102 137258 208186 137494
rect 208422 137258 243866 137494
rect 244102 137258 244186 137494
rect 244422 137258 567866 137494
rect 568102 137258 568186 137494
rect 568422 137258 592062 137494
rect 592298 137258 592382 137494
rect 592618 137258 592650 137494
rect -8726 137174 592650 137258
rect -8726 136938 -8694 137174
rect -8458 136938 -8374 137174
rect -8138 136938 27866 137174
rect 28102 136938 28186 137174
rect 28422 136938 135866 137174
rect 136102 136938 136186 137174
rect 136422 136938 171866 137174
rect 172102 136938 172186 137174
rect 172422 136938 207866 137174
rect 208102 136938 208186 137174
rect 208422 136938 243866 137174
rect 244102 136938 244186 137174
rect 244422 136938 567866 137174
rect 568102 136938 568186 137174
rect 568422 136938 592062 137174
rect 592298 136938 592382 137174
rect 592618 136938 592650 137174
rect -8726 136906 592650 136938
rect -8726 133774 592650 133806
rect -8726 133538 -7734 133774
rect -7498 133538 -7414 133774
rect -7178 133538 24146 133774
rect 24382 133538 24466 133774
rect 24702 133538 60146 133774
rect 60382 133538 60466 133774
rect 60702 133538 96146 133774
rect 96382 133538 96466 133774
rect 96702 133538 132146 133774
rect 132382 133538 132466 133774
rect 132702 133538 168146 133774
rect 168382 133538 168466 133774
rect 168702 133538 204146 133774
rect 204382 133538 204466 133774
rect 204702 133538 240146 133774
rect 240382 133538 240466 133774
rect 240702 133538 564146 133774
rect 564382 133538 564466 133774
rect 564702 133538 591102 133774
rect 591338 133538 591422 133774
rect 591658 133538 592650 133774
rect -8726 133454 592650 133538
rect -8726 133218 -7734 133454
rect -7498 133218 -7414 133454
rect -7178 133218 24146 133454
rect 24382 133218 24466 133454
rect 24702 133218 60146 133454
rect 60382 133218 60466 133454
rect 60702 133218 96146 133454
rect 96382 133218 96466 133454
rect 96702 133218 132146 133454
rect 132382 133218 132466 133454
rect 132702 133218 168146 133454
rect 168382 133218 168466 133454
rect 168702 133218 204146 133454
rect 204382 133218 204466 133454
rect 204702 133218 240146 133454
rect 240382 133218 240466 133454
rect 240702 133218 564146 133454
rect 564382 133218 564466 133454
rect 564702 133218 591102 133454
rect 591338 133218 591422 133454
rect 591658 133218 592650 133454
rect -8726 133186 592650 133218
rect -8726 130054 592650 130086
rect -8726 129818 -6774 130054
rect -6538 129818 -6454 130054
rect -6218 129818 20426 130054
rect 20662 129818 20746 130054
rect 20982 129818 200426 130054
rect 200662 129818 200746 130054
rect 200982 129818 236426 130054
rect 236662 129818 236746 130054
rect 236982 129818 560426 130054
rect 560662 129818 560746 130054
rect 560982 129818 590142 130054
rect 590378 129818 590462 130054
rect 590698 129818 592650 130054
rect -8726 129734 592650 129818
rect -8726 129498 -6774 129734
rect -6538 129498 -6454 129734
rect -6218 129498 20426 129734
rect 20662 129498 20746 129734
rect 20982 129498 200426 129734
rect 200662 129498 200746 129734
rect 200982 129498 236426 129734
rect 236662 129498 236746 129734
rect 236982 129498 560426 129734
rect 560662 129498 560746 129734
rect 560982 129498 590142 129734
rect 590378 129498 590462 129734
rect 590698 129498 592650 129734
rect -8726 129466 592650 129498
rect -8726 126334 592650 126366
rect -8726 126098 -5814 126334
rect -5578 126098 -5494 126334
rect -5258 126098 16706 126334
rect 16942 126098 17026 126334
rect 17262 126098 196706 126334
rect 196942 126098 197026 126334
rect 197262 126098 232706 126334
rect 232942 126098 233026 126334
rect 233262 126098 556706 126334
rect 556942 126098 557026 126334
rect 557262 126098 589182 126334
rect 589418 126098 589502 126334
rect 589738 126098 592650 126334
rect -8726 126014 592650 126098
rect -8726 125778 -5814 126014
rect -5578 125778 -5494 126014
rect -5258 125778 16706 126014
rect 16942 125778 17026 126014
rect 17262 125778 196706 126014
rect 196942 125778 197026 126014
rect 197262 125778 232706 126014
rect 232942 125778 233026 126014
rect 233262 125778 556706 126014
rect 556942 125778 557026 126014
rect 557262 125778 589182 126014
rect 589418 125778 589502 126014
rect 589738 125778 592650 126014
rect -8726 125746 592650 125778
rect -8726 122614 592650 122646
rect -8726 122378 -4854 122614
rect -4618 122378 -4534 122614
rect -4298 122378 12986 122614
rect 13222 122378 13306 122614
rect 13542 122378 156986 122614
rect 157222 122378 157306 122614
rect 157542 122378 228986 122614
rect 229222 122378 229306 122614
rect 229542 122378 552986 122614
rect 553222 122378 553306 122614
rect 553542 122378 588222 122614
rect 588458 122378 588542 122614
rect 588778 122378 592650 122614
rect -8726 122294 592650 122378
rect -8726 122058 -4854 122294
rect -4618 122058 -4534 122294
rect -4298 122058 12986 122294
rect 13222 122058 13306 122294
rect 13542 122058 156986 122294
rect 157222 122058 157306 122294
rect 157542 122058 228986 122294
rect 229222 122058 229306 122294
rect 229542 122058 552986 122294
rect 553222 122058 553306 122294
rect 553542 122058 588222 122294
rect 588458 122058 588542 122294
rect 588778 122058 592650 122294
rect -8726 122026 592650 122058
rect -8726 118894 592650 118926
rect -8726 118658 -3894 118894
rect -3658 118658 -3574 118894
rect -3338 118658 9266 118894
rect 9502 118658 9586 118894
rect 9822 118658 153266 118894
rect 153502 118658 153586 118894
rect 153822 118658 225266 118894
rect 225502 118658 225586 118894
rect 225822 118658 587262 118894
rect 587498 118658 587582 118894
rect 587818 118658 592650 118894
rect -8726 118574 592650 118658
rect -8726 118338 -3894 118574
rect -3658 118338 -3574 118574
rect -3338 118338 9266 118574
rect 9502 118338 9586 118574
rect 9822 118338 153266 118574
rect 153502 118338 153586 118574
rect 153822 118338 225266 118574
rect 225502 118338 225586 118574
rect 225822 118338 587262 118574
rect 587498 118338 587582 118574
rect 587818 118338 592650 118574
rect -8726 118306 592650 118338
rect -8726 115174 592650 115206
rect -8726 114938 -2934 115174
rect -2698 114938 -2614 115174
rect -2378 114938 5546 115174
rect 5782 114938 5866 115174
rect 6102 114938 43610 115174
rect 43846 114938 74330 115174
rect 74566 114938 105050 115174
rect 105286 114938 149546 115174
rect 149782 114938 149866 115174
rect 150102 114938 177610 115174
rect 177846 114938 208330 115174
rect 208566 114938 221546 115174
rect 221782 114938 221866 115174
rect 222102 114938 257546 115174
rect 257782 114938 257866 115174
rect 258102 114938 279610 115174
rect 279846 114938 310330 115174
rect 310566 114938 341050 115174
rect 341286 114938 371770 115174
rect 372006 114938 402490 115174
rect 402726 114938 433210 115174
rect 433446 114938 463930 115174
rect 464166 114938 494650 115174
rect 494886 114938 525370 115174
rect 525606 114938 581546 115174
rect 581782 114938 581866 115174
rect 582102 114938 586302 115174
rect 586538 114938 586622 115174
rect 586858 114938 592650 115174
rect -8726 114854 592650 114938
rect -8726 114618 -2934 114854
rect -2698 114618 -2614 114854
rect -2378 114618 5546 114854
rect 5782 114618 5866 114854
rect 6102 114618 43610 114854
rect 43846 114618 74330 114854
rect 74566 114618 105050 114854
rect 105286 114618 149546 114854
rect 149782 114618 149866 114854
rect 150102 114618 177610 114854
rect 177846 114618 208330 114854
rect 208566 114618 221546 114854
rect 221782 114618 221866 114854
rect 222102 114618 257546 114854
rect 257782 114618 257866 114854
rect 258102 114618 279610 114854
rect 279846 114618 310330 114854
rect 310566 114618 341050 114854
rect 341286 114618 371770 114854
rect 372006 114618 402490 114854
rect 402726 114618 433210 114854
rect 433446 114618 463930 114854
rect 464166 114618 494650 114854
rect 494886 114618 525370 114854
rect 525606 114618 581546 114854
rect 581782 114618 581866 114854
rect 582102 114618 586302 114854
rect 586538 114618 586622 114854
rect 586858 114618 592650 114854
rect -8726 114586 592650 114618
rect -8726 111454 592650 111486
rect -8726 111218 -1974 111454
rect -1738 111218 -1654 111454
rect -1418 111218 1826 111454
rect 2062 111218 2146 111454
rect 2382 111218 28250 111454
rect 28486 111218 58970 111454
rect 59206 111218 89690 111454
rect 89926 111218 120410 111454
rect 120646 111218 145826 111454
rect 146062 111218 146146 111454
rect 146382 111218 162250 111454
rect 162486 111218 192970 111454
rect 193206 111218 217826 111454
rect 218062 111218 218146 111454
rect 218382 111218 253826 111454
rect 254062 111218 254146 111454
rect 254382 111218 264250 111454
rect 264486 111218 294970 111454
rect 295206 111218 325690 111454
rect 325926 111218 356410 111454
rect 356646 111218 387130 111454
rect 387366 111218 417850 111454
rect 418086 111218 448570 111454
rect 448806 111218 479290 111454
rect 479526 111218 510010 111454
rect 510246 111218 540730 111454
rect 540966 111218 577826 111454
rect 578062 111218 578146 111454
rect 578382 111218 585342 111454
rect 585578 111218 585662 111454
rect 585898 111218 592650 111454
rect -8726 111134 592650 111218
rect -8726 110898 -1974 111134
rect -1738 110898 -1654 111134
rect -1418 110898 1826 111134
rect 2062 110898 2146 111134
rect 2382 110898 28250 111134
rect 28486 110898 58970 111134
rect 59206 110898 89690 111134
rect 89926 110898 120410 111134
rect 120646 110898 145826 111134
rect 146062 110898 146146 111134
rect 146382 110898 162250 111134
rect 162486 110898 192970 111134
rect 193206 110898 217826 111134
rect 218062 110898 218146 111134
rect 218382 110898 253826 111134
rect 254062 110898 254146 111134
rect 254382 110898 264250 111134
rect 264486 110898 294970 111134
rect 295206 110898 325690 111134
rect 325926 110898 356410 111134
rect 356646 110898 387130 111134
rect 387366 110898 417850 111134
rect 418086 110898 448570 111134
rect 448806 110898 479290 111134
rect 479526 110898 510010 111134
rect 510246 110898 540730 111134
rect 540966 110898 577826 111134
rect 578062 110898 578146 111134
rect 578382 110898 585342 111134
rect 585578 110898 585662 111134
rect 585898 110898 592650 111134
rect -8726 110866 592650 110898
rect -8726 101494 592650 101526
rect -8726 101258 -8694 101494
rect -8458 101258 -8374 101494
rect -8138 101258 135866 101494
rect 136102 101258 136186 101494
rect 136422 101258 243866 101494
rect 244102 101258 244186 101494
rect 244422 101258 567866 101494
rect 568102 101258 568186 101494
rect 568422 101258 592062 101494
rect 592298 101258 592382 101494
rect 592618 101258 592650 101494
rect -8726 101174 592650 101258
rect -8726 100938 -8694 101174
rect -8458 100938 -8374 101174
rect -8138 100938 135866 101174
rect 136102 100938 136186 101174
rect 136422 100938 243866 101174
rect 244102 100938 244186 101174
rect 244422 100938 567866 101174
rect 568102 100938 568186 101174
rect 568422 100938 592062 101174
rect 592298 100938 592382 101174
rect 592618 100938 592650 101174
rect -8726 100906 592650 100938
rect -8726 97774 592650 97806
rect -8726 97538 -7734 97774
rect -7498 97538 -7414 97774
rect -7178 97538 24146 97774
rect 24382 97538 24466 97774
rect 24702 97538 204146 97774
rect 204382 97538 204466 97774
rect 204702 97538 240146 97774
rect 240382 97538 240466 97774
rect 240702 97538 564146 97774
rect 564382 97538 564466 97774
rect 564702 97538 591102 97774
rect 591338 97538 591422 97774
rect 591658 97538 592650 97774
rect -8726 97454 592650 97538
rect -8726 97218 -7734 97454
rect -7498 97218 -7414 97454
rect -7178 97218 24146 97454
rect 24382 97218 24466 97454
rect 24702 97218 204146 97454
rect 204382 97218 204466 97454
rect 204702 97218 240146 97454
rect 240382 97218 240466 97454
rect 240702 97218 564146 97454
rect 564382 97218 564466 97454
rect 564702 97218 591102 97454
rect 591338 97218 591422 97454
rect 591658 97218 592650 97454
rect -8726 97186 592650 97218
rect -8726 94054 592650 94086
rect -8726 93818 -6774 94054
rect -6538 93818 -6454 94054
rect -6218 93818 20426 94054
rect 20662 93818 20746 94054
rect 20982 93818 200426 94054
rect 200662 93818 200746 94054
rect 200982 93818 236426 94054
rect 236662 93818 236746 94054
rect 236982 93818 560426 94054
rect 560662 93818 560746 94054
rect 560982 93818 590142 94054
rect 590378 93818 590462 94054
rect 590698 93818 592650 94054
rect -8726 93734 592650 93818
rect -8726 93498 -6774 93734
rect -6538 93498 -6454 93734
rect -6218 93498 20426 93734
rect 20662 93498 20746 93734
rect 20982 93498 200426 93734
rect 200662 93498 200746 93734
rect 200982 93498 236426 93734
rect 236662 93498 236746 93734
rect 236982 93498 560426 93734
rect 560662 93498 560746 93734
rect 560982 93498 590142 93734
rect 590378 93498 590462 93734
rect 590698 93498 592650 93734
rect -8726 93466 592650 93498
rect -8726 90334 592650 90366
rect -8726 90098 -5814 90334
rect -5578 90098 -5494 90334
rect -5258 90098 16706 90334
rect 16942 90098 17026 90334
rect 17262 90098 196706 90334
rect 196942 90098 197026 90334
rect 197262 90098 232706 90334
rect 232942 90098 233026 90334
rect 233262 90098 556706 90334
rect 556942 90098 557026 90334
rect 557262 90098 589182 90334
rect 589418 90098 589502 90334
rect 589738 90098 592650 90334
rect -8726 90014 592650 90098
rect -8726 89778 -5814 90014
rect -5578 89778 -5494 90014
rect -5258 89778 16706 90014
rect 16942 89778 17026 90014
rect 17262 89778 196706 90014
rect 196942 89778 197026 90014
rect 197262 89778 232706 90014
rect 232942 89778 233026 90014
rect 233262 89778 556706 90014
rect 556942 89778 557026 90014
rect 557262 89778 589182 90014
rect 589418 89778 589502 90014
rect 589738 89778 592650 90014
rect -8726 89746 592650 89778
rect -8726 86614 592650 86646
rect -8726 86378 -4854 86614
rect -4618 86378 -4534 86614
rect -4298 86378 12986 86614
rect 13222 86378 13306 86614
rect 13542 86378 156986 86614
rect 157222 86378 157306 86614
rect 157542 86378 228986 86614
rect 229222 86378 229306 86614
rect 229542 86378 552986 86614
rect 553222 86378 553306 86614
rect 553542 86378 588222 86614
rect 588458 86378 588542 86614
rect 588778 86378 592650 86614
rect -8726 86294 592650 86378
rect -8726 86058 -4854 86294
rect -4618 86058 -4534 86294
rect -4298 86058 12986 86294
rect 13222 86058 13306 86294
rect 13542 86058 156986 86294
rect 157222 86058 157306 86294
rect 157542 86058 228986 86294
rect 229222 86058 229306 86294
rect 229542 86058 552986 86294
rect 553222 86058 553306 86294
rect 553542 86058 588222 86294
rect 588458 86058 588542 86294
rect 588778 86058 592650 86294
rect -8726 86026 592650 86058
rect -8726 82894 592650 82926
rect -8726 82658 -3894 82894
rect -3658 82658 -3574 82894
rect -3338 82658 9266 82894
rect 9502 82658 9586 82894
rect 9822 82658 153266 82894
rect 153502 82658 153586 82894
rect 153822 82658 225266 82894
rect 225502 82658 225586 82894
rect 225822 82658 587262 82894
rect 587498 82658 587582 82894
rect 587818 82658 592650 82894
rect -8726 82574 592650 82658
rect -8726 82338 -3894 82574
rect -3658 82338 -3574 82574
rect -3338 82338 9266 82574
rect 9502 82338 9586 82574
rect 9822 82338 153266 82574
rect 153502 82338 153586 82574
rect 153822 82338 225266 82574
rect 225502 82338 225586 82574
rect 225822 82338 587262 82574
rect 587498 82338 587582 82574
rect 587818 82338 592650 82574
rect -8726 82306 592650 82338
rect -8726 79174 592650 79206
rect -8726 78938 -2934 79174
rect -2698 78938 -2614 79174
rect -2378 78938 5546 79174
rect 5782 78938 5866 79174
rect 6102 78938 43610 79174
rect 43846 78938 74330 79174
rect 74566 78938 105050 79174
rect 105286 78938 149546 79174
rect 149782 78938 149866 79174
rect 150102 78938 177610 79174
rect 177846 78938 208330 79174
rect 208566 78938 221546 79174
rect 221782 78938 221866 79174
rect 222102 78938 257546 79174
rect 257782 78938 257866 79174
rect 258102 78938 279610 79174
rect 279846 78938 310330 79174
rect 310566 78938 341050 79174
rect 341286 78938 371770 79174
rect 372006 78938 402490 79174
rect 402726 78938 433210 79174
rect 433446 78938 463930 79174
rect 464166 78938 494650 79174
rect 494886 78938 525370 79174
rect 525606 78938 581546 79174
rect 581782 78938 581866 79174
rect 582102 78938 586302 79174
rect 586538 78938 586622 79174
rect 586858 78938 592650 79174
rect -8726 78854 592650 78938
rect -8726 78618 -2934 78854
rect -2698 78618 -2614 78854
rect -2378 78618 5546 78854
rect 5782 78618 5866 78854
rect 6102 78618 43610 78854
rect 43846 78618 74330 78854
rect 74566 78618 105050 78854
rect 105286 78618 149546 78854
rect 149782 78618 149866 78854
rect 150102 78618 177610 78854
rect 177846 78618 208330 78854
rect 208566 78618 221546 78854
rect 221782 78618 221866 78854
rect 222102 78618 257546 78854
rect 257782 78618 257866 78854
rect 258102 78618 279610 78854
rect 279846 78618 310330 78854
rect 310566 78618 341050 78854
rect 341286 78618 371770 78854
rect 372006 78618 402490 78854
rect 402726 78618 433210 78854
rect 433446 78618 463930 78854
rect 464166 78618 494650 78854
rect 494886 78618 525370 78854
rect 525606 78618 581546 78854
rect 581782 78618 581866 78854
rect 582102 78618 586302 78854
rect 586538 78618 586622 78854
rect 586858 78618 592650 78854
rect -8726 78586 592650 78618
rect -8726 75454 592650 75486
rect -8726 75218 -1974 75454
rect -1738 75218 -1654 75454
rect -1418 75218 1826 75454
rect 2062 75218 2146 75454
rect 2382 75218 28250 75454
rect 28486 75218 58970 75454
rect 59206 75218 89690 75454
rect 89926 75218 120410 75454
rect 120646 75218 145826 75454
rect 146062 75218 146146 75454
rect 146382 75218 162250 75454
rect 162486 75218 192970 75454
rect 193206 75218 217826 75454
rect 218062 75218 218146 75454
rect 218382 75218 253826 75454
rect 254062 75218 254146 75454
rect 254382 75218 264250 75454
rect 264486 75218 294970 75454
rect 295206 75218 325690 75454
rect 325926 75218 356410 75454
rect 356646 75218 387130 75454
rect 387366 75218 417850 75454
rect 418086 75218 448570 75454
rect 448806 75218 479290 75454
rect 479526 75218 510010 75454
rect 510246 75218 540730 75454
rect 540966 75218 577826 75454
rect 578062 75218 578146 75454
rect 578382 75218 585342 75454
rect 585578 75218 585662 75454
rect 585898 75218 592650 75454
rect -8726 75134 592650 75218
rect -8726 74898 -1974 75134
rect -1738 74898 -1654 75134
rect -1418 74898 1826 75134
rect 2062 74898 2146 75134
rect 2382 74898 28250 75134
rect 28486 74898 58970 75134
rect 59206 74898 89690 75134
rect 89926 74898 120410 75134
rect 120646 74898 145826 75134
rect 146062 74898 146146 75134
rect 146382 74898 162250 75134
rect 162486 74898 192970 75134
rect 193206 74898 217826 75134
rect 218062 74898 218146 75134
rect 218382 74898 253826 75134
rect 254062 74898 254146 75134
rect 254382 74898 264250 75134
rect 264486 74898 294970 75134
rect 295206 74898 325690 75134
rect 325926 74898 356410 75134
rect 356646 74898 387130 75134
rect 387366 74898 417850 75134
rect 418086 74898 448570 75134
rect 448806 74898 479290 75134
rect 479526 74898 510010 75134
rect 510246 74898 540730 75134
rect 540966 74898 577826 75134
rect 578062 74898 578146 75134
rect 578382 74898 585342 75134
rect 585578 74898 585662 75134
rect 585898 74898 592650 75134
rect -8726 74866 592650 74898
rect -8726 65494 592650 65526
rect -8726 65258 -8694 65494
rect -8458 65258 -8374 65494
rect -8138 65258 135866 65494
rect 136102 65258 136186 65494
rect 136422 65258 243866 65494
rect 244102 65258 244186 65494
rect 244422 65258 567866 65494
rect 568102 65258 568186 65494
rect 568422 65258 592062 65494
rect 592298 65258 592382 65494
rect 592618 65258 592650 65494
rect -8726 65174 592650 65258
rect -8726 64938 -8694 65174
rect -8458 64938 -8374 65174
rect -8138 64938 135866 65174
rect 136102 64938 136186 65174
rect 136422 64938 243866 65174
rect 244102 64938 244186 65174
rect 244422 64938 567866 65174
rect 568102 64938 568186 65174
rect 568422 64938 592062 65174
rect 592298 64938 592382 65174
rect 592618 64938 592650 65174
rect -8726 64906 592650 64938
rect -8726 61774 592650 61806
rect -8726 61538 -7734 61774
rect -7498 61538 -7414 61774
rect -7178 61538 24146 61774
rect 24382 61538 24466 61774
rect 24702 61538 204146 61774
rect 204382 61538 204466 61774
rect 204702 61538 240146 61774
rect 240382 61538 240466 61774
rect 240702 61538 564146 61774
rect 564382 61538 564466 61774
rect 564702 61538 591102 61774
rect 591338 61538 591422 61774
rect 591658 61538 592650 61774
rect -8726 61454 592650 61538
rect -8726 61218 -7734 61454
rect -7498 61218 -7414 61454
rect -7178 61218 24146 61454
rect 24382 61218 24466 61454
rect 24702 61218 204146 61454
rect 204382 61218 204466 61454
rect 204702 61218 240146 61454
rect 240382 61218 240466 61454
rect 240702 61218 564146 61454
rect 564382 61218 564466 61454
rect 564702 61218 591102 61454
rect 591338 61218 591422 61454
rect 591658 61218 592650 61454
rect -8726 61186 592650 61218
rect -8726 58054 592650 58086
rect -8726 57818 -6774 58054
rect -6538 57818 -6454 58054
rect -6218 57818 20426 58054
rect 20662 57818 20746 58054
rect 20982 57818 200426 58054
rect 200662 57818 200746 58054
rect 200982 57818 236426 58054
rect 236662 57818 236746 58054
rect 236982 57818 560426 58054
rect 560662 57818 560746 58054
rect 560982 57818 590142 58054
rect 590378 57818 590462 58054
rect 590698 57818 592650 58054
rect -8726 57734 592650 57818
rect -8726 57498 -6774 57734
rect -6538 57498 -6454 57734
rect -6218 57498 20426 57734
rect 20662 57498 20746 57734
rect 20982 57498 200426 57734
rect 200662 57498 200746 57734
rect 200982 57498 236426 57734
rect 236662 57498 236746 57734
rect 236982 57498 560426 57734
rect 560662 57498 560746 57734
rect 560982 57498 590142 57734
rect 590378 57498 590462 57734
rect 590698 57498 592650 57734
rect -8726 57466 592650 57498
rect -8726 54334 592650 54366
rect -8726 54098 -5814 54334
rect -5578 54098 -5494 54334
rect -5258 54098 16706 54334
rect 16942 54098 17026 54334
rect 17262 54098 196706 54334
rect 196942 54098 197026 54334
rect 197262 54098 232706 54334
rect 232942 54098 233026 54334
rect 233262 54098 556706 54334
rect 556942 54098 557026 54334
rect 557262 54098 589182 54334
rect 589418 54098 589502 54334
rect 589738 54098 592650 54334
rect -8726 54014 592650 54098
rect -8726 53778 -5814 54014
rect -5578 53778 -5494 54014
rect -5258 53778 16706 54014
rect 16942 53778 17026 54014
rect 17262 53778 196706 54014
rect 196942 53778 197026 54014
rect 197262 53778 232706 54014
rect 232942 53778 233026 54014
rect 233262 53778 556706 54014
rect 556942 53778 557026 54014
rect 557262 53778 589182 54014
rect 589418 53778 589502 54014
rect 589738 53778 592650 54014
rect -8726 53746 592650 53778
rect -8726 50614 592650 50646
rect -8726 50378 -4854 50614
rect -4618 50378 -4534 50614
rect -4298 50378 12986 50614
rect 13222 50378 13306 50614
rect 13542 50378 156986 50614
rect 157222 50378 157306 50614
rect 157542 50378 192986 50614
rect 193222 50378 193306 50614
rect 193542 50378 228986 50614
rect 229222 50378 229306 50614
rect 229542 50378 552986 50614
rect 553222 50378 553306 50614
rect 553542 50378 588222 50614
rect 588458 50378 588542 50614
rect 588778 50378 592650 50614
rect -8726 50294 592650 50378
rect -8726 50058 -4854 50294
rect -4618 50058 -4534 50294
rect -4298 50058 12986 50294
rect 13222 50058 13306 50294
rect 13542 50058 156986 50294
rect 157222 50058 157306 50294
rect 157542 50058 192986 50294
rect 193222 50058 193306 50294
rect 193542 50058 228986 50294
rect 229222 50058 229306 50294
rect 229542 50058 552986 50294
rect 553222 50058 553306 50294
rect 553542 50058 588222 50294
rect 588458 50058 588542 50294
rect 588778 50058 592650 50294
rect -8726 50026 592650 50058
rect -8726 46894 592650 46926
rect -8726 46658 -3894 46894
rect -3658 46658 -3574 46894
rect -3338 46658 9266 46894
rect 9502 46658 9586 46894
rect 9822 46658 153266 46894
rect 153502 46658 153586 46894
rect 153822 46658 189266 46894
rect 189502 46658 189586 46894
rect 189822 46658 225266 46894
rect 225502 46658 225586 46894
rect 225822 46658 587262 46894
rect 587498 46658 587582 46894
rect 587818 46658 592650 46894
rect -8726 46574 592650 46658
rect -8726 46338 -3894 46574
rect -3658 46338 -3574 46574
rect -3338 46338 9266 46574
rect 9502 46338 9586 46574
rect 9822 46338 153266 46574
rect 153502 46338 153586 46574
rect 153822 46338 189266 46574
rect 189502 46338 189586 46574
rect 189822 46338 225266 46574
rect 225502 46338 225586 46574
rect 225822 46338 587262 46574
rect 587498 46338 587582 46574
rect 587818 46338 592650 46574
rect -8726 46306 592650 46338
rect -8726 43174 592650 43206
rect -8726 42938 -2934 43174
rect -2698 42938 -2614 43174
rect -2378 42938 5546 43174
rect 5782 42938 5866 43174
rect 6102 42938 43610 43174
rect 43846 42938 74330 43174
rect 74566 42938 105050 43174
rect 105286 42938 149546 43174
rect 149782 42938 149866 43174
rect 150102 42938 185546 43174
rect 185782 42938 185866 43174
rect 186102 42938 221546 43174
rect 221782 42938 221866 43174
rect 222102 42938 257546 43174
rect 257782 42938 257866 43174
rect 258102 42938 279610 43174
rect 279846 42938 310330 43174
rect 310566 42938 341050 43174
rect 341286 42938 371770 43174
rect 372006 42938 402490 43174
rect 402726 42938 433210 43174
rect 433446 42938 463930 43174
rect 464166 42938 494650 43174
rect 494886 42938 525370 43174
rect 525606 42938 581546 43174
rect 581782 42938 581866 43174
rect 582102 42938 586302 43174
rect 586538 42938 586622 43174
rect 586858 42938 592650 43174
rect -8726 42854 592650 42938
rect -8726 42618 -2934 42854
rect -2698 42618 -2614 42854
rect -2378 42618 5546 42854
rect 5782 42618 5866 42854
rect 6102 42618 43610 42854
rect 43846 42618 74330 42854
rect 74566 42618 105050 42854
rect 105286 42618 149546 42854
rect 149782 42618 149866 42854
rect 150102 42618 185546 42854
rect 185782 42618 185866 42854
rect 186102 42618 221546 42854
rect 221782 42618 221866 42854
rect 222102 42618 257546 42854
rect 257782 42618 257866 42854
rect 258102 42618 279610 42854
rect 279846 42618 310330 42854
rect 310566 42618 341050 42854
rect 341286 42618 371770 42854
rect 372006 42618 402490 42854
rect 402726 42618 433210 42854
rect 433446 42618 463930 42854
rect 464166 42618 494650 42854
rect 494886 42618 525370 42854
rect 525606 42618 581546 42854
rect 581782 42618 581866 42854
rect 582102 42618 586302 42854
rect 586538 42618 586622 42854
rect 586858 42618 592650 42854
rect -8726 42586 592650 42618
rect -8726 39454 592650 39486
rect -8726 39218 -1974 39454
rect -1738 39218 -1654 39454
rect -1418 39218 1826 39454
rect 2062 39218 2146 39454
rect 2382 39218 28250 39454
rect 28486 39218 58970 39454
rect 59206 39218 89690 39454
rect 89926 39218 120410 39454
rect 120646 39218 145826 39454
rect 146062 39218 146146 39454
rect 146382 39218 181826 39454
rect 182062 39218 182146 39454
rect 182382 39218 217826 39454
rect 218062 39218 218146 39454
rect 218382 39218 253826 39454
rect 254062 39218 254146 39454
rect 254382 39218 289826 39454
rect 290062 39218 290146 39454
rect 290382 39218 325826 39454
rect 326062 39218 326146 39454
rect 326382 39218 361826 39454
rect 362062 39218 362146 39454
rect 362382 39218 397826 39454
rect 398062 39218 398146 39454
rect 398382 39218 433826 39454
rect 434062 39218 434146 39454
rect 434382 39218 469826 39454
rect 470062 39218 470146 39454
rect 470382 39218 505826 39454
rect 506062 39218 506146 39454
rect 506382 39218 541826 39454
rect 542062 39218 542146 39454
rect 542382 39218 577826 39454
rect 578062 39218 578146 39454
rect 578382 39218 585342 39454
rect 585578 39218 585662 39454
rect 585898 39218 592650 39454
rect -8726 39134 592650 39218
rect -8726 38898 -1974 39134
rect -1738 38898 -1654 39134
rect -1418 38898 1826 39134
rect 2062 38898 2146 39134
rect 2382 38898 28250 39134
rect 28486 38898 58970 39134
rect 59206 38898 89690 39134
rect 89926 38898 120410 39134
rect 120646 38898 145826 39134
rect 146062 38898 146146 39134
rect 146382 38898 181826 39134
rect 182062 38898 182146 39134
rect 182382 38898 217826 39134
rect 218062 38898 218146 39134
rect 218382 38898 253826 39134
rect 254062 38898 254146 39134
rect 254382 38898 289826 39134
rect 290062 38898 290146 39134
rect 290382 38898 325826 39134
rect 326062 38898 326146 39134
rect 326382 38898 361826 39134
rect 362062 38898 362146 39134
rect 362382 38898 397826 39134
rect 398062 38898 398146 39134
rect 398382 38898 433826 39134
rect 434062 38898 434146 39134
rect 434382 38898 469826 39134
rect 470062 38898 470146 39134
rect 470382 38898 505826 39134
rect 506062 38898 506146 39134
rect 506382 38898 541826 39134
rect 542062 38898 542146 39134
rect 542382 38898 577826 39134
rect 578062 38898 578146 39134
rect 578382 38898 585342 39134
rect 585578 38898 585662 39134
rect 585898 38898 592650 39134
rect -8726 38866 592650 38898
rect -8726 29494 592650 29526
rect -8726 29258 -8694 29494
rect -8458 29258 -8374 29494
rect -8138 29258 135866 29494
rect 136102 29258 136186 29494
rect 136422 29258 171866 29494
rect 172102 29258 172186 29494
rect 172422 29258 207866 29494
rect 208102 29258 208186 29494
rect 208422 29258 243866 29494
rect 244102 29258 244186 29494
rect 244422 29258 279866 29494
rect 280102 29258 280186 29494
rect 280422 29258 315866 29494
rect 316102 29258 316186 29494
rect 316422 29258 351866 29494
rect 352102 29258 352186 29494
rect 352422 29258 387866 29494
rect 388102 29258 388186 29494
rect 388422 29258 423866 29494
rect 424102 29258 424186 29494
rect 424422 29258 459866 29494
rect 460102 29258 460186 29494
rect 460422 29258 495866 29494
rect 496102 29258 496186 29494
rect 496422 29258 531866 29494
rect 532102 29258 532186 29494
rect 532422 29258 567866 29494
rect 568102 29258 568186 29494
rect 568422 29258 592062 29494
rect 592298 29258 592382 29494
rect 592618 29258 592650 29494
rect -8726 29174 592650 29258
rect -8726 28938 -8694 29174
rect -8458 28938 -8374 29174
rect -8138 28938 135866 29174
rect 136102 28938 136186 29174
rect 136422 28938 171866 29174
rect 172102 28938 172186 29174
rect 172422 28938 207866 29174
rect 208102 28938 208186 29174
rect 208422 28938 243866 29174
rect 244102 28938 244186 29174
rect 244422 28938 279866 29174
rect 280102 28938 280186 29174
rect 280422 28938 315866 29174
rect 316102 28938 316186 29174
rect 316422 28938 351866 29174
rect 352102 28938 352186 29174
rect 352422 28938 387866 29174
rect 388102 28938 388186 29174
rect 388422 28938 423866 29174
rect 424102 28938 424186 29174
rect 424422 28938 459866 29174
rect 460102 28938 460186 29174
rect 460422 28938 495866 29174
rect 496102 28938 496186 29174
rect 496422 28938 531866 29174
rect 532102 28938 532186 29174
rect 532422 28938 567866 29174
rect 568102 28938 568186 29174
rect 568422 28938 592062 29174
rect 592298 28938 592382 29174
rect 592618 28938 592650 29174
rect -8726 28906 592650 28938
rect -8726 25774 592650 25806
rect -8726 25538 -7734 25774
rect -7498 25538 -7414 25774
rect -7178 25538 24146 25774
rect 24382 25538 24466 25774
rect 24702 25538 168146 25774
rect 168382 25538 168466 25774
rect 168702 25538 204146 25774
rect 204382 25538 204466 25774
rect 204702 25538 240146 25774
rect 240382 25538 240466 25774
rect 240702 25538 276146 25774
rect 276382 25538 276466 25774
rect 276702 25538 312146 25774
rect 312382 25538 312466 25774
rect 312702 25538 348146 25774
rect 348382 25538 348466 25774
rect 348702 25538 384146 25774
rect 384382 25538 384466 25774
rect 384702 25538 420146 25774
rect 420382 25538 420466 25774
rect 420702 25538 456146 25774
rect 456382 25538 456466 25774
rect 456702 25538 492146 25774
rect 492382 25538 492466 25774
rect 492702 25538 528146 25774
rect 528382 25538 528466 25774
rect 528702 25538 564146 25774
rect 564382 25538 564466 25774
rect 564702 25538 591102 25774
rect 591338 25538 591422 25774
rect 591658 25538 592650 25774
rect -8726 25454 592650 25538
rect -8726 25218 -7734 25454
rect -7498 25218 -7414 25454
rect -7178 25218 24146 25454
rect 24382 25218 24466 25454
rect 24702 25218 168146 25454
rect 168382 25218 168466 25454
rect 168702 25218 204146 25454
rect 204382 25218 204466 25454
rect 204702 25218 240146 25454
rect 240382 25218 240466 25454
rect 240702 25218 276146 25454
rect 276382 25218 276466 25454
rect 276702 25218 312146 25454
rect 312382 25218 312466 25454
rect 312702 25218 348146 25454
rect 348382 25218 348466 25454
rect 348702 25218 384146 25454
rect 384382 25218 384466 25454
rect 384702 25218 420146 25454
rect 420382 25218 420466 25454
rect 420702 25218 456146 25454
rect 456382 25218 456466 25454
rect 456702 25218 492146 25454
rect 492382 25218 492466 25454
rect 492702 25218 528146 25454
rect 528382 25218 528466 25454
rect 528702 25218 564146 25454
rect 564382 25218 564466 25454
rect 564702 25218 591102 25454
rect 591338 25218 591422 25454
rect 591658 25218 592650 25454
rect -8726 25186 592650 25218
rect -8726 22054 592650 22086
rect -8726 21818 -6774 22054
rect -6538 21818 -6454 22054
rect -6218 21818 20426 22054
rect 20662 21818 20746 22054
rect 20982 21818 56426 22054
rect 56662 21818 56746 22054
rect 56982 21818 92426 22054
rect 92662 21818 92746 22054
rect 92982 21818 128426 22054
rect 128662 21818 128746 22054
rect 128982 21818 164426 22054
rect 164662 21818 164746 22054
rect 164982 21818 200426 22054
rect 200662 21818 200746 22054
rect 200982 21818 236426 22054
rect 236662 21818 236746 22054
rect 236982 21818 272426 22054
rect 272662 21818 272746 22054
rect 272982 21818 308426 22054
rect 308662 21818 308746 22054
rect 308982 21818 344426 22054
rect 344662 21818 344746 22054
rect 344982 21818 380426 22054
rect 380662 21818 380746 22054
rect 380982 21818 416426 22054
rect 416662 21818 416746 22054
rect 416982 21818 452426 22054
rect 452662 21818 452746 22054
rect 452982 21818 488426 22054
rect 488662 21818 488746 22054
rect 488982 21818 524426 22054
rect 524662 21818 524746 22054
rect 524982 21818 560426 22054
rect 560662 21818 560746 22054
rect 560982 21818 590142 22054
rect 590378 21818 590462 22054
rect 590698 21818 592650 22054
rect -8726 21734 592650 21818
rect -8726 21498 -6774 21734
rect -6538 21498 -6454 21734
rect -6218 21498 20426 21734
rect 20662 21498 20746 21734
rect 20982 21498 56426 21734
rect 56662 21498 56746 21734
rect 56982 21498 92426 21734
rect 92662 21498 92746 21734
rect 92982 21498 128426 21734
rect 128662 21498 128746 21734
rect 128982 21498 164426 21734
rect 164662 21498 164746 21734
rect 164982 21498 200426 21734
rect 200662 21498 200746 21734
rect 200982 21498 236426 21734
rect 236662 21498 236746 21734
rect 236982 21498 272426 21734
rect 272662 21498 272746 21734
rect 272982 21498 308426 21734
rect 308662 21498 308746 21734
rect 308982 21498 344426 21734
rect 344662 21498 344746 21734
rect 344982 21498 380426 21734
rect 380662 21498 380746 21734
rect 380982 21498 416426 21734
rect 416662 21498 416746 21734
rect 416982 21498 452426 21734
rect 452662 21498 452746 21734
rect 452982 21498 488426 21734
rect 488662 21498 488746 21734
rect 488982 21498 524426 21734
rect 524662 21498 524746 21734
rect 524982 21498 560426 21734
rect 560662 21498 560746 21734
rect 560982 21498 590142 21734
rect 590378 21498 590462 21734
rect 590698 21498 592650 21734
rect -8726 21466 592650 21498
rect -8726 18334 592650 18366
rect -8726 18098 -5814 18334
rect -5578 18098 -5494 18334
rect -5258 18098 16706 18334
rect 16942 18098 17026 18334
rect 17262 18098 52706 18334
rect 52942 18098 53026 18334
rect 53262 18098 88706 18334
rect 88942 18098 89026 18334
rect 89262 18098 124706 18334
rect 124942 18098 125026 18334
rect 125262 18098 160706 18334
rect 160942 18098 161026 18334
rect 161262 18098 196706 18334
rect 196942 18098 197026 18334
rect 197262 18098 232706 18334
rect 232942 18098 233026 18334
rect 233262 18098 268706 18334
rect 268942 18098 269026 18334
rect 269262 18098 304706 18334
rect 304942 18098 305026 18334
rect 305262 18098 340706 18334
rect 340942 18098 341026 18334
rect 341262 18098 376706 18334
rect 376942 18098 377026 18334
rect 377262 18098 412706 18334
rect 412942 18098 413026 18334
rect 413262 18098 448706 18334
rect 448942 18098 449026 18334
rect 449262 18098 484706 18334
rect 484942 18098 485026 18334
rect 485262 18098 520706 18334
rect 520942 18098 521026 18334
rect 521262 18098 556706 18334
rect 556942 18098 557026 18334
rect 557262 18098 589182 18334
rect 589418 18098 589502 18334
rect 589738 18098 592650 18334
rect -8726 18014 592650 18098
rect -8726 17778 -5814 18014
rect -5578 17778 -5494 18014
rect -5258 17778 16706 18014
rect 16942 17778 17026 18014
rect 17262 17778 52706 18014
rect 52942 17778 53026 18014
rect 53262 17778 88706 18014
rect 88942 17778 89026 18014
rect 89262 17778 124706 18014
rect 124942 17778 125026 18014
rect 125262 17778 160706 18014
rect 160942 17778 161026 18014
rect 161262 17778 196706 18014
rect 196942 17778 197026 18014
rect 197262 17778 232706 18014
rect 232942 17778 233026 18014
rect 233262 17778 268706 18014
rect 268942 17778 269026 18014
rect 269262 17778 304706 18014
rect 304942 17778 305026 18014
rect 305262 17778 340706 18014
rect 340942 17778 341026 18014
rect 341262 17778 376706 18014
rect 376942 17778 377026 18014
rect 377262 17778 412706 18014
rect 412942 17778 413026 18014
rect 413262 17778 448706 18014
rect 448942 17778 449026 18014
rect 449262 17778 484706 18014
rect 484942 17778 485026 18014
rect 485262 17778 520706 18014
rect 520942 17778 521026 18014
rect 521262 17778 556706 18014
rect 556942 17778 557026 18014
rect 557262 17778 589182 18014
rect 589418 17778 589502 18014
rect 589738 17778 592650 18014
rect -8726 17746 592650 17778
rect -8726 14614 592650 14646
rect -8726 14378 -4854 14614
rect -4618 14378 -4534 14614
rect -4298 14378 12986 14614
rect 13222 14378 13306 14614
rect 13542 14378 48986 14614
rect 49222 14378 49306 14614
rect 49542 14378 84986 14614
rect 85222 14378 85306 14614
rect 85542 14378 120986 14614
rect 121222 14378 121306 14614
rect 121542 14378 156986 14614
rect 157222 14378 157306 14614
rect 157542 14378 192986 14614
rect 193222 14378 193306 14614
rect 193542 14378 228986 14614
rect 229222 14378 229306 14614
rect 229542 14378 264986 14614
rect 265222 14378 265306 14614
rect 265542 14378 300986 14614
rect 301222 14378 301306 14614
rect 301542 14378 336986 14614
rect 337222 14378 337306 14614
rect 337542 14378 372986 14614
rect 373222 14378 373306 14614
rect 373542 14378 408986 14614
rect 409222 14378 409306 14614
rect 409542 14378 444986 14614
rect 445222 14378 445306 14614
rect 445542 14378 480986 14614
rect 481222 14378 481306 14614
rect 481542 14378 516986 14614
rect 517222 14378 517306 14614
rect 517542 14378 552986 14614
rect 553222 14378 553306 14614
rect 553542 14378 588222 14614
rect 588458 14378 588542 14614
rect 588778 14378 592650 14614
rect -8726 14294 592650 14378
rect -8726 14058 -4854 14294
rect -4618 14058 -4534 14294
rect -4298 14058 12986 14294
rect 13222 14058 13306 14294
rect 13542 14058 48986 14294
rect 49222 14058 49306 14294
rect 49542 14058 84986 14294
rect 85222 14058 85306 14294
rect 85542 14058 120986 14294
rect 121222 14058 121306 14294
rect 121542 14058 156986 14294
rect 157222 14058 157306 14294
rect 157542 14058 192986 14294
rect 193222 14058 193306 14294
rect 193542 14058 228986 14294
rect 229222 14058 229306 14294
rect 229542 14058 264986 14294
rect 265222 14058 265306 14294
rect 265542 14058 300986 14294
rect 301222 14058 301306 14294
rect 301542 14058 336986 14294
rect 337222 14058 337306 14294
rect 337542 14058 372986 14294
rect 373222 14058 373306 14294
rect 373542 14058 408986 14294
rect 409222 14058 409306 14294
rect 409542 14058 444986 14294
rect 445222 14058 445306 14294
rect 445542 14058 480986 14294
rect 481222 14058 481306 14294
rect 481542 14058 516986 14294
rect 517222 14058 517306 14294
rect 517542 14058 552986 14294
rect 553222 14058 553306 14294
rect 553542 14058 588222 14294
rect 588458 14058 588542 14294
rect 588778 14058 592650 14294
rect -8726 14026 592650 14058
rect -8726 10894 592650 10926
rect -8726 10658 -3894 10894
rect -3658 10658 -3574 10894
rect -3338 10658 9266 10894
rect 9502 10658 9586 10894
rect 9822 10658 45266 10894
rect 45502 10658 45586 10894
rect 45822 10658 81266 10894
rect 81502 10658 81586 10894
rect 81822 10658 117266 10894
rect 117502 10658 117586 10894
rect 117822 10658 153266 10894
rect 153502 10658 153586 10894
rect 153822 10658 189266 10894
rect 189502 10658 189586 10894
rect 189822 10658 225266 10894
rect 225502 10658 225586 10894
rect 225822 10658 261266 10894
rect 261502 10658 261586 10894
rect 261822 10658 297266 10894
rect 297502 10658 297586 10894
rect 297822 10658 333266 10894
rect 333502 10658 333586 10894
rect 333822 10658 369266 10894
rect 369502 10658 369586 10894
rect 369822 10658 405266 10894
rect 405502 10658 405586 10894
rect 405822 10658 441266 10894
rect 441502 10658 441586 10894
rect 441822 10658 477266 10894
rect 477502 10658 477586 10894
rect 477822 10658 513266 10894
rect 513502 10658 513586 10894
rect 513822 10658 549266 10894
rect 549502 10658 549586 10894
rect 549822 10658 587262 10894
rect 587498 10658 587582 10894
rect 587818 10658 592650 10894
rect -8726 10574 592650 10658
rect -8726 10338 -3894 10574
rect -3658 10338 -3574 10574
rect -3338 10338 9266 10574
rect 9502 10338 9586 10574
rect 9822 10338 45266 10574
rect 45502 10338 45586 10574
rect 45822 10338 81266 10574
rect 81502 10338 81586 10574
rect 81822 10338 117266 10574
rect 117502 10338 117586 10574
rect 117822 10338 153266 10574
rect 153502 10338 153586 10574
rect 153822 10338 189266 10574
rect 189502 10338 189586 10574
rect 189822 10338 225266 10574
rect 225502 10338 225586 10574
rect 225822 10338 261266 10574
rect 261502 10338 261586 10574
rect 261822 10338 297266 10574
rect 297502 10338 297586 10574
rect 297822 10338 333266 10574
rect 333502 10338 333586 10574
rect 333822 10338 369266 10574
rect 369502 10338 369586 10574
rect 369822 10338 405266 10574
rect 405502 10338 405586 10574
rect 405822 10338 441266 10574
rect 441502 10338 441586 10574
rect 441822 10338 477266 10574
rect 477502 10338 477586 10574
rect 477822 10338 513266 10574
rect 513502 10338 513586 10574
rect 513822 10338 549266 10574
rect 549502 10338 549586 10574
rect 549822 10338 587262 10574
rect 587498 10338 587582 10574
rect 587818 10338 592650 10574
rect -8726 10306 592650 10338
rect -8726 7174 592650 7206
rect -8726 6938 -2934 7174
rect -2698 6938 -2614 7174
rect -2378 6938 5546 7174
rect 5782 6938 5866 7174
rect 6102 6938 41546 7174
rect 41782 6938 41866 7174
rect 42102 6938 77546 7174
rect 77782 6938 77866 7174
rect 78102 6938 113546 7174
rect 113782 6938 113866 7174
rect 114102 6938 149546 7174
rect 149782 6938 149866 7174
rect 150102 6938 185546 7174
rect 185782 6938 185866 7174
rect 186102 6938 221546 7174
rect 221782 6938 221866 7174
rect 222102 6938 257546 7174
rect 257782 6938 257866 7174
rect 258102 6938 293546 7174
rect 293782 6938 293866 7174
rect 294102 6938 329546 7174
rect 329782 6938 329866 7174
rect 330102 6938 365546 7174
rect 365782 6938 365866 7174
rect 366102 6938 401546 7174
rect 401782 6938 401866 7174
rect 402102 6938 437546 7174
rect 437782 6938 437866 7174
rect 438102 6938 473546 7174
rect 473782 6938 473866 7174
rect 474102 6938 509546 7174
rect 509782 6938 509866 7174
rect 510102 6938 545546 7174
rect 545782 6938 545866 7174
rect 546102 6938 581546 7174
rect 581782 6938 581866 7174
rect 582102 6938 586302 7174
rect 586538 6938 586622 7174
rect 586858 6938 592650 7174
rect -8726 6854 592650 6938
rect -8726 6618 -2934 6854
rect -2698 6618 -2614 6854
rect -2378 6618 5546 6854
rect 5782 6618 5866 6854
rect 6102 6618 41546 6854
rect 41782 6618 41866 6854
rect 42102 6618 77546 6854
rect 77782 6618 77866 6854
rect 78102 6618 113546 6854
rect 113782 6618 113866 6854
rect 114102 6618 149546 6854
rect 149782 6618 149866 6854
rect 150102 6618 185546 6854
rect 185782 6618 185866 6854
rect 186102 6618 221546 6854
rect 221782 6618 221866 6854
rect 222102 6618 257546 6854
rect 257782 6618 257866 6854
rect 258102 6618 293546 6854
rect 293782 6618 293866 6854
rect 294102 6618 329546 6854
rect 329782 6618 329866 6854
rect 330102 6618 365546 6854
rect 365782 6618 365866 6854
rect 366102 6618 401546 6854
rect 401782 6618 401866 6854
rect 402102 6618 437546 6854
rect 437782 6618 437866 6854
rect 438102 6618 473546 6854
rect 473782 6618 473866 6854
rect 474102 6618 509546 6854
rect 509782 6618 509866 6854
rect 510102 6618 545546 6854
rect 545782 6618 545866 6854
rect 546102 6618 581546 6854
rect 581782 6618 581866 6854
rect 582102 6618 586302 6854
rect 586538 6618 586622 6854
rect 586858 6618 592650 6854
rect -8726 6586 592650 6618
rect -8726 3454 592650 3486
rect -8726 3218 -1974 3454
rect -1738 3218 -1654 3454
rect -1418 3218 1826 3454
rect 2062 3218 2146 3454
rect 2382 3218 37826 3454
rect 38062 3218 38146 3454
rect 38382 3218 73826 3454
rect 74062 3218 74146 3454
rect 74382 3218 109826 3454
rect 110062 3218 110146 3454
rect 110382 3218 145826 3454
rect 146062 3218 146146 3454
rect 146382 3218 181826 3454
rect 182062 3218 182146 3454
rect 182382 3218 217826 3454
rect 218062 3218 218146 3454
rect 218382 3218 253826 3454
rect 254062 3218 254146 3454
rect 254382 3218 289826 3454
rect 290062 3218 290146 3454
rect 290382 3218 325826 3454
rect 326062 3218 326146 3454
rect 326382 3218 361826 3454
rect 362062 3218 362146 3454
rect 362382 3218 397826 3454
rect 398062 3218 398146 3454
rect 398382 3218 433826 3454
rect 434062 3218 434146 3454
rect 434382 3218 469826 3454
rect 470062 3218 470146 3454
rect 470382 3218 505826 3454
rect 506062 3218 506146 3454
rect 506382 3218 541826 3454
rect 542062 3218 542146 3454
rect 542382 3218 577826 3454
rect 578062 3218 578146 3454
rect 578382 3218 585342 3454
rect 585578 3218 585662 3454
rect 585898 3218 592650 3454
rect -8726 3134 592650 3218
rect -8726 2898 -1974 3134
rect -1738 2898 -1654 3134
rect -1418 2898 1826 3134
rect 2062 2898 2146 3134
rect 2382 2898 37826 3134
rect 38062 2898 38146 3134
rect 38382 2898 73826 3134
rect 74062 2898 74146 3134
rect 74382 2898 109826 3134
rect 110062 2898 110146 3134
rect 110382 2898 145826 3134
rect 146062 2898 146146 3134
rect 146382 2898 181826 3134
rect 182062 2898 182146 3134
rect 182382 2898 217826 3134
rect 218062 2898 218146 3134
rect 218382 2898 253826 3134
rect 254062 2898 254146 3134
rect 254382 2898 289826 3134
rect 290062 2898 290146 3134
rect 290382 2898 325826 3134
rect 326062 2898 326146 3134
rect 326382 2898 361826 3134
rect 362062 2898 362146 3134
rect 362382 2898 397826 3134
rect 398062 2898 398146 3134
rect 398382 2898 433826 3134
rect 434062 2898 434146 3134
rect 434382 2898 469826 3134
rect 470062 2898 470146 3134
rect 470382 2898 505826 3134
rect 506062 2898 506146 3134
rect 506382 2898 541826 3134
rect 542062 2898 542146 3134
rect 542382 2898 577826 3134
rect 578062 2898 578146 3134
rect 578382 2898 585342 3134
rect 585578 2898 585662 3134
rect 585898 2898 592650 3134
rect -8726 2866 592650 2898
rect -2006 -346 585930 -314
rect -2006 -582 -1974 -346
rect -1738 -582 -1654 -346
rect -1418 -582 1826 -346
rect 2062 -582 2146 -346
rect 2382 -582 37826 -346
rect 38062 -582 38146 -346
rect 38382 -582 73826 -346
rect 74062 -582 74146 -346
rect 74382 -582 109826 -346
rect 110062 -582 110146 -346
rect 110382 -582 145826 -346
rect 146062 -582 146146 -346
rect 146382 -582 181826 -346
rect 182062 -582 182146 -346
rect 182382 -582 217826 -346
rect 218062 -582 218146 -346
rect 218382 -582 253826 -346
rect 254062 -582 254146 -346
rect 254382 -582 289826 -346
rect 290062 -582 290146 -346
rect 290382 -582 325826 -346
rect 326062 -582 326146 -346
rect 326382 -582 361826 -346
rect 362062 -582 362146 -346
rect 362382 -582 397826 -346
rect 398062 -582 398146 -346
rect 398382 -582 433826 -346
rect 434062 -582 434146 -346
rect 434382 -582 469826 -346
rect 470062 -582 470146 -346
rect 470382 -582 505826 -346
rect 506062 -582 506146 -346
rect 506382 -582 541826 -346
rect 542062 -582 542146 -346
rect 542382 -582 577826 -346
rect 578062 -582 578146 -346
rect 578382 -582 585342 -346
rect 585578 -582 585662 -346
rect 585898 -582 585930 -346
rect -2006 -666 585930 -582
rect -2006 -902 -1974 -666
rect -1738 -902 -1654 -666
rect -1418 -902 1826 -666
rect 2062 -902 2146 -666
rect 2382 -902 37826 -666
rect 38062 -902 38146 -666
rect 38382 -902 73826 -666
rect 74062 -902 74146 -666
rect 74382 -902 109826 -666
rect 110062 -902 110146 -666
rect 110382 -902 145826 -666
rect 146062 -902 146146 -666
rect 146382 -902 181826 -666
rect 182062 -902 182146 -666
rect 182382 -902 217826 -666
rect 218062 -902 218146 -666
rect 218382 -902 253826 -666
rect 254062 -902 254146 -666
rect 254382 -902 289826 -666
rect 290062 -902 290146 -666
rect 290382 -902 325826 -666
rect 326062 -902 326146 -666
rect 326382 -902 361826 -666
rect 362062 -902 362146 -666
rect 362382 -902 397826 -666
rect 398062 -902 398146 -666
rect 398382 -902 433826 -666
rect 434062 -902 434146 -666
rect 434382 -902 469826 -666
rect 470062 -902 470146 -666
rect 470382 -902 505826 -666
rect 506062 -902 506146 -666
rect 506382 -902 541826 -666
rect 542062 -902 542146 -666
rect 542382 -902 577826 -666
rect 578062 -902 578146 -666
rect 578382 -902 585342 -666
rect 585578 -902 585662 -666
rect 585898 -902 585930 -666
rect -2006 -934 585930 -902
rect -2966 -1306 586890 -1274
rect -2966 -1542 -2934 -1306
rect -2698 -1542 -2614 -1306
rect -2378 -1542 5546 -1306
rect 5782 -1542 5866 -1306
rect 6102 -1542 41546 -1306
rect 41782 -1542 41866 -1306
rect 42102 -1542 77546 -1306
rect 77782 -1542 77866 -1306
rect 78102 -1542 113546 -1306
rect 113782 -1542 113866 -1306
rect 114102 -1542 149546 -1306
rect 149782 -1542 149866 -1306
rect 150102 -1542 185546 -1306
rect 185782 -1542 185866 -1306
rect 186102 -1542 221546 -1306
rect 221782 -1542 221866 -1306
rect 222102 -1542 257546 -1306
rect 257782 -1542 257866 -1306
rect 258102 -1542 293546 -1306
rect 293782 -1542 293866 -1306
rect 294102 -1542 329546 -1306
rect 329782 -1542 329866 -1306
rect 330102 -1542 365546 -1306
rect 365782 -1542 365866 -1306
rect 366102 -1542 401546 -1306
rect 401782 -1542 401866 -1306
rect 402102 -1542 437546 -1306
rect 437782 -1542 437866 -1306
rect 438102 -1542 473546 -1306
rect 473782 -1542 473866 -1306
rect 474102 -1542 509546 -1306
rect 509782 -1542 509866 -1306
rect 510102 -1542 545546 -1306
rect 545782 -1542 545866 -1306
rect 546102 -1542 581546 -1306
rect 581782 -1542 581866 -1306
rect 582102 -1542 586302 -1306
rect 586538 -1542 586622 -1306
rect 586858 -1542 586890 -1306
rect -2966 -1626 586890 -1542
rect -2966 -1862 -2934 -1626
rect -2698 -1862 -2614 -1626
rect -2378 -1862 5546 -1626
rect 5782 -1862 5866 -1626
rect 6102 -1862 41546 -1626
rect 41782 -1862 41866 -1626
rect 42102 -1862 77546 -1626
rect 77782 -1862 77866 -1626
rect 78102 -1862 113546 -1626
rect 113782 -1862 113866 -1626
rect 114102 -1862 149546 -1626
rect 149782 -1862 149866 -1626
rect 150102 -1862 185546 -1626
rect 185782 -1862 185866 -1626
rect 186102 -1862 221546 -1626
rect 221782 -1862 221866 -1626
rect 222102 -1862 257546 -1626
rect 257782 -1862 257866 -1626
rect 258102 -1862 293546 -1626
rect 293782 -1862 293866 -1626
rect 294102 -1862 329546 -1626
rect 329782 -1862 329866 -1626
rect 330102 -1862 365546 -1626
rect 365782 -1862 365866 -1626
rect 366102 -1862 401546 -1626
rect 401782 -1862 401866 -1626
rect 402102 -1862 437546 -1626
rect 437782 -1862 437866 -1626
rect 438102 -1862 473546 -1626
rect 473782 -1862 473866 -1626
rect 474102 -1862 509546 -1626
rect 509782 -1862 509866 -1626
rect 510102 -1862 545546 -1626
rect 545782 -1862 545866 -1626
rect 546102 -1862 581546 -1626
rect 581782 -1862 581866 -1626
rect 582102 -1862 586302 -1626
rect 586538 -1862 586622 -1626
rect 586858 -1862 586890 -1626
rect -2966 -1894 586890 -1862
rect -3926 -2266 587850 -2234
rect -3926 -2502 -3894 -2266
rect -3658 -2502 -3574 -2266
rect -3338 -2502 9266 -2266
rect 9502 -2502 9586 -2266
rect 9822 -2502 45266 -2266
rect 45502 -2502 45586 -2266
rect 45822 -2502 81266 -2266
rect 81502 -2502 81586 -2266
rect 81822 -2502 117266 -2266
rect 117502 -2502 117586 -2266
rect 117822 -2502 153266 -2266
rect 153502 -2502 153586 -2266
rect 153822 -2502 189266 -2266
rect 189502 -2502 189586 -2266
rect 189822 -2502 225266 -2266
rect 225502 -2502 225586 -2266
rect 225822 -2502 261266 -2266
rect 261502 -2502 261586 -2266
rect 261822 -2502 297266 -2266
rect 297502 -2502 297586 -2266
rect 297822 -2502 333266 -2266
rect 333502 -2502 333586 -2266
rect 333822 -2502 369266 -2266
rect 369502 -2502 369586 -2266
rect 369822 -2502 405266 -2266
rect 405502 -2502 405586 -2266
rect 405822 -2502 441266 -2266
rect 441502 -2502 441586 -2266
rect 441822 -2502 477266 -2266
rect 477502 -2502 477586 -2266
rect 477822 -2502 513266 -2266
rect 513502 -2502 513586 -2266
rect 513822 -2502 549266 -2266
rect 549502 -2502 549586 -2266
rect 549822 -2502 587262 -2266
rect 587498 -2502 587582 -2266
rect 587818 -2502 587850 -2266
rect -3926 -2586 587850 -2502
rect -3926 -2822 -3894 -2586
rect -3658 -2822 -3574 -2586
rect -3338 -2822 9266 -2586
rect 9502 -2822 9586 -2586
rect 9822 -2822 45266 -2586
rect 45502 -2822 45586 -2586
rect 45822 -2822 81266 -2586
rect 81502 -2822 81586 -2586
rect 81822 -2822 117266 -2586
rect 117502 -2822 117586 -2586
rect 117822 -2822 153266 -2586
rect 153502 -2822 153586 -2586
rect 153822 -2822 189266 -2586
rect 189502 -2822 189586 -2586
rect 189822 -2822 225266 -2586
rect 225502 -2822 225586 -2586
rect 225822 -2822 261266 -2586
rect 261502 -2822 261586 -2586
rect 261822 -2822 297266 -2586
rect 297502 -2822 297586 -2586
rect 297822 -2822 333266 -2586
rect 333502 -2822 333586 -2586
rect 333822 -2822 369266 -2586
rect 369502 -2822 369586 -2586
rect 369822 -2822 405266 -2586
rect 405502 -2822 405586 -2586
rect 405822 -2822 441266 -2586
rect 441502 -2822 441586 -2586
rect 441822 -2822 477266 -2586
rect 477502 -2822 477586 -2586
rect 477822 -2822 513266 -2586
rect 513502 -2822 513586 -2586
rect 513822 -2822 549266 -2586
rect 549502 -2822 549586 -2586
rect 549822 -2822 587262 -2586
rect 587498 -2822 587582 -2586
rect 587818 -2822 587850 -2586
rect -3926 -2854 587850 -2822
rect -4886 -3226 588810 -3194
rect -4886 -3462 -4854 -3226
rect -4618 -3462 -4534 -3226
rect -4298 -3462 12986 -3226
rect 13222 -3462 13306 -3226
rect 13542 -3462 48986 -3226
rect 49222 -3462 49306 -3226
rect 49542 -3462 84986 -3226
rect 85222 -3462 85306 -3226
rect 85542 -3462 120986 -3226
rect 121222 -3462 121306 -3226
rect 121542 -3462 156986 -3226
rect 157222 -3462 157306 -3226
rect 157542 -3462 192986 -3226
rect 193222 -3462 193306 -3226
rect 193542 -3462 228986 -3226
rect 229222 -3462 229306 -3226
rect 229542 -3462 264986 -3226
rect 265222 -3462 265306 -3226
rect 265542 -3462 300986 -3226
rect 301222 -3462 301306 -3226
rect 301542 -3462 336986 -3226
rect 337222 -3462 337306 -3226
rect 337542 -3462 372986 -3226
rect 373222 -3462 373306 -3226
rect 373542 -3462 408986 -3226
rect 409222 -3462 409306 -3226
rect 409542 -3462 444986 -3226
rect 445222 -3462 445306 -3226
rect 445542 -3462 480986 -3226
rect 481222 -3462 481306 -3226
rect 481542 -3462 516986 -3226
rect 517222 -3462 517306 -3226
rect 517542 -3462 552986 -3226
rect 553222 -3462 553306 -3226
rect 553542 -3462 588222 -3226
rect 588458 -3462 588542 -3226
rect 588778 -3462 588810 -3226
rect -4886 -3546 588810 -3462
rect -4886 -3782 -4854 -3546
rect -4618 -3782 -4534 -3546
rect -4298 -3782 12986 -3546
rect 13222 -3782 13306 -3546
rect 13542 -3782 48986 -3546
rect 49222 -3782 49306 -3546
rect 49542 -3782 84986 -3546
rect 85222 -3782 85306 -3546
rect 85542 -3782 120986 -3546
rect 121222 -3782 121306 -3546
rect 121542 -3782 156986 -3546
rect 157222 -3782 157306 -3546
rect 157542 -3782 192986 -3546
rect 193222 -3782 193306 -3546
rect 193542 -3782 228986 -3546
rect 229222 -3782 229306 -3546
rect 229542 -3782 264986 -3546
rect 265222 -3782 265306 -3546
rect 265542 -3782 300986 -3546
rect 301222 -3782 301306 -3546
rect 301542 -3782 336986 -3546
rect 337222 -3782 337306 -3546
rect 337542 -3782 372986 -3546
rect 373222 -3782 373306 -3546
rect 373542 -3782 408986 -3546
rect 409222 -3782 409306 -3546
rect 409542 -3782 444986 -3546
rect 445222 -3782 445306 -3546
rect 445542 -3782 480986 -3546
rect 481222 -3782 481306 -3546
rect 481542 -3782 516986 -3546
rect 517222 -3782 517306 -3546
rect 517542 -3782 552986 -3546
rect 553222 -3782 553306 -3546
rect 553542 -3782 588222 -3546
rect 588458 -3782 588542 -3546
rect 588778 -3782 588810 -3546
rect -4886 -3814 588810 -3782
rect -5846 -4186 589770 -4154
rect -5846 -4422 -5814 -4186
rect -5578 -4422 -5494 -4186
rect -5258 -4422 16706 -4186
rect 16942 -4422 17026 -4186
rect 17262 -4422 52706 -4186
rect 52942 -4422 53026 -4186
rect 53262 -4422 88706 -4186
rect 88942 -4422 89026 -4186
rect 89262 -4422 124706 -4186
rect 124942 -4422 125026 -4186
rect 125262 -4422 160706 -4186
rect 160942 -4422 161026 -4186
rect 161262 -4422 196706 -4186
rect 196942 -4422 197026 -4186
rect 197262 -4422 232706 -4186
rect 232942 -4422 233026 -4186
rect 233262 -4422 268706 -4186
rect 268942 -4422 269026 -4186
rect 269262 -4422 304706 -4186
rect 304942 -4422 305026 -4186
rect 305262 -4422 340706 -4186
rect 340942 -4422 341026 -4186
rect 341262 -4422 376706 -4186
rect 376942 -4422 377026 -4186
rect 377262 -4422 412706 -4186
rect 412942 -4422 413026 -4186
rect 413262 -4422 448706 -4186
rect 448942 -4422 449026 -4186
rect 449262 -4422 484706 -4186
rect 484942 -4422 485026 -4186
rect 485262 -4422 520706 -4186
rect 520942 -4422 521026 -4186
rect 521262 -4422 556706 -4186
rect 556942 -4422 557026 -4186
rect 557262 -4422 589182 -4186
rect 589418 -4422 589502 -4186
rect 589738 -4422 589770 -4186
rect -5846 -4506 589770 -4422
rect -5846 -4742 -5814 -4506
rect -5578 -4742 -5494 -4506
rect -5258 -4742 16706 -4506
rect 16942 -4742 17026 -4506
rect 17262 -4742 52706 -4506
rect 52942 -4742 53026 -4506
rect 53262 -4742 88706 -4506
rect 88942 -4742 89026 -4506
rect 89262 -4742 124706 -4506
rect 124942 -4742 125026 -4506
rect 125262 -4742 160706 -4506
rect 160942 -4742 161026 -4506
rect 161262 -4742 196706 -4506
rect 196942 -4742 197026 -4506
rect 197262 -4742 232706 -4506
rect 232942 -4742 233026 -4506
rect 233262 -4742 268706 -4506
rect 268942 -4742 269026 -4506
rect 269262 -4742 304706 -4506
rect 304942 -4742 305026 -4506
rect 305262 -4742 340706 -4506
rect 340942 -4742 341026 -4506
rect 341262 -4742 376706 -4506
rect 376942 -4742 377026 -4506
rect 377262 -4742 412706 -4506
rect 412942 -4742 413026 -4506
rect 413262 -4742 448706 -4506
rect 448942 -4742 449026 -4506
rect 449262 -4742 484706 -4506
rect 484942 -4742 485026 -4506
rect 485262 -4742 520706 -4506
rect 520942 -4742 521026 -4506
rect 521262 -4742 556706 -4506
rect 556942 -4742 557026 -4506
rect 557262 -4742 589182 -4506
rect 589418 -4742 589502 -4506
rect 589738 -4742 589770 -4506
rect -5846 -4774 589770 -4742
rect -6806 -5146 590730 -5114
rect -6806 -5382 -6774 -5146
rect -6538 -5382 -6454 -5146
rect -6218 -5382 20426 -5146
rect 20662 -5382 20746 -5146
rect 20982 -5382 56426 -5146
rect 56662 -5382 56746 -5146
rect 56982 -5382 92426 -5146
rect 92662 -5382 92746 -5146
rect 92982 -5382 128426 -5146
rect 128662 -5382 128746 -5146
rect 128982 -5382 164426 -5146
rect 164662 -5382 164746 -5146
rect 164982 -5382 200426 -5146
rect 200662 -5382 200746 -5146
rect 200982 -5382 236426 -5146
rect 236662 -5382 236746 -5146
rect 236982 -5382 272426 -5146
rect 272662 -5382 272746 -5146
rect 272982 -5382 308426 -5146
rect 308662 -5382 308746 -5146
rect 308982 -5382 344426 -5146
rect 344662 -5382 344746 -5146
rect 344982 -5382 380426 -5146
rect 380662 -5382 380746 -5146
rect 380982 -5382 416426 -5146
rect 416662 -5382 416746 -5146
rect 416982 -5382 452426 -5146
rect 452662 -5382 452746 -5146
rect 452982 -5382 488426 -5146
rect 488662 -5382 488746 -5146
rect 488982 -5382 524426 -5146
rect 524662 -5382 524746 -5146
rect 524982 -5382 560426 -5146
rect 560662 -5382 560746 -5146
rect 560982 -5382 590142 -5146
rect 590378 -5382 590462 -5146
rect 590698 -5382 590730 -5146
rect -6806 -5466 590730 -5382
rect -6806 -5702 -6774 -5466
rect -6538 -5702 -6454 -5466
rect -6218 -5702 20426 -5466
rect 20662 -5702 20746 -5466
rect 20982 -5702 56426 -5466
rect 56662 -5702 56746 -5466
rect 56982 -5702 92426 -5466
rect 92662 -5702 92746 -5466
rect 92982 -5702 128426 -5466
rect 128662 -5702 128746 -5466
rect 128982 -5702 164426 -5466
rect 164662 -5702 164746 -5466
rect 164982 -5702 200426 -5466
rect 200662 -5702 200746 -5466
rect 200982 -5702 236426 -5466
rect 236662 -5702 236746 -5466
rect 236982 -5702 272426 -5466
rect 272662 -5702 272746 -5466
rect 272982 -5702 308426 -5466
rect 308662 -5702 308746 -5466
rect 308982 -5702 344426 -5466
rect 344662 -5702 344746 -5466
rect 344982 -5702 380426 -5466
rect 380662 -5702 380746 -5466
rect 380982 -5702 416426 -5466
rect 416662 -5702 416746 -5466
rect 416982 -5702 452426 -5466
rect 452662 -5702 452746 -5466
rect 452982 -5702 488426 -5466
rect 488662 -5702 488746 -5466
rect 488982 -5702 524426 -5466
rect 524662 -5702 524746 -5466
rect 524982 -5702 560426 -5466
rect 560662 -5702 560746 -5466
rect 560982 -5702 590142 -5466
rect 590378 -5702 590462 -5466
rect 590698 -5702 590730 -5466
rect -6806 -5734 590730 -5702
rect -7766 -6106 591690 -6074
rect -7766 -6342 -7734 -6106
rect -7498 -6342 -7414 -6106
rect -7178 -6342 24146 -6106
rect 24382 -6342 24466 -6106
rect 24702 -6342 168146 -6106
rect 168382 -6342 168466 -6106
rect 168702 -6342 204146 -6106
rect 204382 -6342 204466 -6106
rect 204702 -6342 240146 -6106
rect 240382 -6342 240466 -6106
rect 240702 -6342 276146 -6106
rect 276382 -6342 276466 -6106
rect 276702 -6342 312146 -6106
rect 312382 -6342 312466 -6106
rect 312702 -6342 348146 -6106
rect 348382 -6342 348466 -6106
rect 348702 -6342 384146 -6106
rect 384382 -6342 384466 -6106
rect 384702 -6342 420146 -6106
rect 420382 -6342 420466 -6106
rect 420702 -6342 456146 -6106
rect 456382 -6342 456466 -6106
rect 456702 -6342 492146 -6106
rect 492382 -6342 492466 -6106
rect 492702 -6342 528146 -6106
rect 528382 -6342 528466 -6106
rect 528702 -6342 564146 -6106
rect 564382 -6342 564466 -6106
rect 564702 -6342 591102 -6106
rect 591338 -6342 591422 -6106
rect 591658 -6342 591690 -6106
rect -7766 -6426 591690 -6342
rect -7766 -6662 -7734 -6426
rect -7498 -6662 -7414 -6426
rect -7178 -6662 24146 -6426
rect 24382 -6662 24466 -6426
rect 24702 -6662 168146 -6426
rect 168382 -6662 168466 -6426
rect 168702 -6662 204146 -6426
rect 204382 -6662 204466 -6426
rect 204702 -6662 240146 -6426
rect 240382 -6662 240466 -6426
rect 240702 -6662 276146 -6426
rect 276382 -6662 276466 -6426
rect 276702 -6662 312146 -6426
rect 312382 -6662 312466 -6426
rect 312702 -6662 348146 -6426
rect 348382 -6662 348466 -6426
rect 348702 -6662 384146 -6426
rect 384382 -6662 384466 -6426
rect 384702 -6662 420146 -6426
rect 420382 -6662 420466 -6426
rect 420702 -6662 456146 -6426
rect 456382 -6662 456466 -6426
rect 456702 -6662 492146 -6426
rect 492382 -6662 492466 -6426
rect 492702 -6662 528146 -6426
rect 528382 -6662 528466 -6426
rect 528702 -6662 564146 -6426
rect 564382 -6662 564466 -6426
rect 564702 -6662 591102 -6426
rect 591338 -6662 591422 -6426
rect 591658 -6662 591690 -6426
rect -7766 -6694 591690 -6662
rect -8726 -7066 592650 -7034
rect -8726 -7302 -8694 -7066
rect -8458 -7302 -8374 -7066
rect -8138 -7302 135866 -7066
rect 136102 -7302 136186 -7066
rect 136422 -7302 171866 -7066
rect 172102 -7302 172186 -7066
rect 172422 -7302 207866 -7066
rect 208102 -7302 208186 -7066
rect 208422 -7302 243866 -7066
rect 244102 -7302 244186 -7066
rect 244422 -7302 279866 -7066
rect 280102 -7302 280186 -7066
rect 280422 -7302 315866 -7066
rect 316102 -7302 316186 -7066
rect 316422 -7302 351866 -7066
rect 352102 -7302 352186 -7066
rect 352422 -7302 387866 -7066
rect 388102 -7302 388186 -7066
rect 388422 -7302 423866 -7066
rect 424102 -7302 424186 -7066
rect 424422 -7302 459866 -7066
rect 460102 -7302 460186 -7066
rect 460422 -7302 495866 -7066
rect 496102 -7302 496186 -7066
rect 496422 -7302 531866 -7066
rect 532102 -7302 532186 -7066
rect 532422 -7302 567866 -7066
rect 568102 -7302 568186 -7066
rect 568422 -7302 592062 -7066
rect 592298 -7302 592382 -7066
rect 592618 -7302 592650 -7066
rect -8726 -7386 592650 -7302
rect -8726 -7622 -8694 -7386
rect -8458 -7622 -8374 -7386
rect -8138 -7622 135866 -7386
rect 136102 -7622 136186 -7386
rect 136422 -7622 171866 -7386
rect 172102 -7622 172186 -7386
rect 172422 -7622 207866 -7386
rect 208102 -7622 208186 -7386
rect 208422 -7622 243866 -7386
rect 244102 -7622 244186 -7386
rect 244422 -7622 279866 -7386
rect 280102 -7622 280186 -7386
rect 280422 -7622 315866 -7386
rect 316102 -7622 316186 -7386
rect 316422 -7622 351866 -7386
rect 352102 -7622 352186 -7386
rect 352422 -7622 387866 -7386
rect 388102 -7622 388186 -7386
rect 388422 -7622 423866 -7386
rect 424102 -7622 424186 -7386
rect 424422 -7622 459866 -7386
rect 460102 -7622 460186 -7386
rect 460422 -7622 495866 -7386
rect 496102 -7622 496186 -7386
rect 496422 -7622 531866 -7386
rect 532102 -7622 532186 -7386
rect 532422 -7622 567866 -7386
rect 568102 -7622 568186 -7386
rect 568422 -7622 592062 -7386
rect 592298 -7622 592382 -7386
rect 592618 -7622 592650 -7386
rect -8726 -7654 592650 -7622
use core0  mprj_core0
timestamp 0
transform 1 0 30000 0 1 160000
box 1066 2128 80000 161616
use core1  mprj_core1
timestamp 0
transform 1 0 30000 0 1 440000
box 1066 2128 80000 157808
use dcache  mprj_dcache
timestamp 0
transform 1 0 260000 0 1 40000
box 0 2128 289971 278361
use icache  mprj_icache_0
timestamp 0
transform 1 0 253600 0 1 380000
box 0 2128 318872 117552
use icache  mprj_icache_1
timestamp 0
transform 1 0 253600 0 1 529600
box 0 2128 318872 117552
use int_ram  mprj_int_ram
timestamp 0
transform 1 0 24000 0 1 24000
box 1066 1838 110000 107760
use interconnect_inner  mprj_interconnect_inner
timestamp 0
transform 1 0 158000 0 1 270000
box 0 0 60000 157808
use interconnect_outer  mprj_interconnect_outer
timestamp 0
transform 1 0 158000 0 1 52000
box 0 0 58880 80000
<< labels >>
flabel metal3 s 583520 285276 584960 285516 0 FreeSans 960 0 0 0 analog_io[0]
port 0 nsew signal bidirectional
flabel metal2 s 446098 703520 446210 704960 0 FreeSans 448 90 0 0 analog_io[10]
port 1 nsew signal bidirectional
flabel metal2 s 381146 703520 381258 704960 0 FreeSans 448 90 0 0 analog_io[11]
port 2 nsew signal bidirectional
flabel metal2 s 316286 703520 316398 704960 0 FreeSans 448 90 0 0 analog_io[12]
port 3 nsew signal bidirectional
flabel metal2 s 251426 703520 251538 704960 0 FreeSans 448 90 0 0 analog_io[13]
port 4 nsew signal bidirectional
flabel metal2 s 186474 703520 186586 704960 0 FreeSans 448 90 0 0 analog_io[14]
port 5 nsew signal bidirectional
flabel metal2 s 121614 703520 121726 704960 0 FreeSans 448 90 0 0 analog_io[15]
port 6 nsew signal bidirectional
flabel metal2 s 56754 703520 56866 704960 0 FreeSans 448 90 0 0 analog_io[16]
port 7 nsew signal bidirectional
flabel metal3 s -960 697220 480 697460 0 FreeSans 960 0 0 0 analog_io[17]
port 8 nsew signal bidirectional
flabel metal3 s -960 644996 480 645236 0 FreeSans 960 0 0 0 analog_io[18]
port 9 nsew signal bidirectional
flabel metal3 s -960 592908 480 593148 0 FreeSans 960 0 0 0 analog_io[19]
port 10 nsew signal bidirectional
flabel metal3 s 583520 338452 584960 338692 0 FreeSans 960 0 0 0 analog_io[1]
port 11 nsew signal bidirectional
flabel metal3 s -960 540684 480 540924 0 FreeSans 960 0 0 0 analog_io[20]
port 12 nsew signal bidirectional
flabel metal3 s -960 488596 480 488836 0 FreeSans 960 0 0 0 analog_io[21]
port 13 nsew signal bidirectional
flabel metal3 s -960 436508 480 436748 0 FreeSans 960 0 0 0 analog_io[22]
port 14 nsew signal bidirectional
flabel metal3 s -960 384284 480 384524 0 FreeSans 960 0 0 0 analog_io[23]
port 15 nsew signal bidirectional
flabel metal3 s -960 332196 480 332436 0 FreeSans 960 0 0 0 analog_io[24]
port 16 nsew signal bidirectional
flabel metal3 s -960 279972 480 280212 0 FreeSans 960 0 0 0 analog_io[25]
port 17 nsew signal bidirectional
flabel metal3 s -960 227884 480 228124 0 FreeSans 960 0 0 0 analog_io[26]
port 18 nsew signal bidirectional
flabel metal3 s -960 175796 480 176036 0 FreeSans 960 0 0 0 analog_io[27]
port 19 nsew signal bidirectional
flabel metal3 s -960 123572 480 123812 0 FreeSans 960 0 0 0 analog_io[28]
port 20 nsew signal bidirectional
flabel metal3 s 583520 391628 584960 391868 0 FreeSans 960 0 0 0 analog_io[2]
port 21 nsew signal bidirectional
flabel metal3 s 583520 444668 584960 444908 0 FreeSans 960 0 0 0 analog_io[3]
port 22 nsew signal bidirectional
flabel metal3 s 583520 497844 584960 498084 0 FreeSans 960 0 0 0 analog_io[4]
port 23 nsew signal bidirectional
flabel metal3 s 583520 551020 584960 551260 0 FreeSans 960 0 0 0 analog_io[5]
port 24 nsew signal bidirectional
flabel metal3 s 583520 604060 584960 604300 0 FreeSans 960 0 0 0 analog_io[6]
port 25 nsew signal bidirectional
flabel metal3 s 583520 657236 584960 657476 0 FreeSans 960 0 0 0 analog_io[7]
port 26 nsew signal bidirectional
flabel metal2 s 575818 703520 575930 704960 0 FreeSans 448 90 0 0 analog_io[8]
port 27 nsew signal bidirectional
flabel metal2 s 510958 703520 511070 704960 0 FreeSans 448 90 0 0 analog_io[9]
port 28 nsew signal bidirectional
flabel metal3 s 583520 6476 584960 6716 0 FreeSans 960 0 0 0 io_in[0]
port 29 nsew signal input
flabel metal3 s 583520 457996 584960 458236 0 FreeSans 960 0 0 0 io_in[10]
port 30 nsew signal input
flabel metal3 s 583520 511172 584960 511412 0 FreeSans 960 0 0 0 io_in[11]
port 31 nsew signal input
flabel metal3 s 583520 564212 584960 564452 0 FreeSans 960 0 0 0 io_in[12]
port 32 nsew signal input
flabel metal3 s 583520 617388 584960 617628 0 FreeSans 960 0 0 0 io_in[13]
port 33 nsew signal input
flabel metal3 s 583520 670564 584960 670804 0 FreeSans 960 0 0 0 io_in[14]
port 34 nsew signal input
flabel metal2 s 559626 703520 559738 704960 0 FreeSans 448 90 0 0 io_in[15]
port 35 nsew signal input
flabel metal2 s 494766 703520 494878 704960 0 FreeSans 448 90 0 0 io_in[16]
port 36 nsew signal input
flabel metal2 s 429814 703520 429926 704960 0 FreeSans 448 90 0 0 io_in[17]
port 37 nsew signal input
flabel metal2 s 364954 703520 365066 704960 0 FreeSans 448 90 0 0 io_in[18]
port 38 nsew signal input
flabel metal2 s 300094 703520 300206 704960 0 FreeSans 448 90 0 0 io_in[19]
port 39 nsew signal input
flabel metal3 s 583520 46188 584960 46428 0 FreeSans 960 0 0 0 io_in[1]
port 40 nsew signal input
flabel metal2 s 235142 703520 235254 704960 0 FreeSans 448 90 0 0 io_in[20]
port 41 nsew signal input
flabel metal2 s 170282 703520 170394 704960 0 FreeSans 448 90 0 0 io_in[21]
port 42 nsew signal input
flabel metal2 s 105422 703520 105534 704960 0 FreeSans 448 90 0 0 io_in[22]
port 43 nsew signal input
flabel metal2 s 40470 703520 40582 704960 0 FreeSans 448 90 0 0 io_in[23]
port 44 nsew signal input
flabel metal3 s -960 684164 480 684404 0 FreeSans 960 0 0 0 io_in[24]
port 45 nsew signal input
flabel metal3 s -960 631940 480 632180 0 FreeSans 960 0 0 0 io_in[25]
port 46 nsew signal input
flabel metal3 s -960 579852 480 580092 0 FreeSans 960 0 0 0 io_in[26]
port 47 nsew signal input
flabel metal3 s -960 527764 480 528004 0 FreeSans 960 0 0 0 io_in[27]
port 48 nsew signal input
flabel metal3 s -960 475540 480 475780 0 FreeSans 960 0 0 0 io_in[28]
port 49 nsew signal input
flabel metal3 s -960 423452 480 423692 0 FreeSans 960 0 0 0 io_in[29]
port 50 nsew signal input
flabel metal3 s 583520 86036 584960 86276 0 FreeSans 960 0 0 0 io_in[2]
port 51 nsew signal input
flabel metal3 s -960 371228 480 371468 0 FreeSans 960 0 0 0 io_in[30]
port 52 nsew signal input
flabel metal3 s -960 319140 480 319380 0 FreeSans 960 0 0 0 io_in[31]
port 53 nsew signal input
flabel metal3 s -960 267052 480 267292 0 FreeSans 960 0 0 0 io_in[32]
port 54 nsew signal input
flabel metal3 s -960 214828 480 215068 0 FreeSans 960 0 0 0 io_in[33]
port 55 nsew signal input
flabel metal3 s -960 162740 480 162980 0 FreeSans 960 0 0 0 io_in[34]
port 56 nsew signal input
flabel metal3 s -960 110516 480 110756 0 FreeSans 960 0 0 0 io_in[35]
port 57 nsew signal input
flabel metal3 s -960 71484 480 71724 0 FreeSans 960 0 0 0 io_in[36]
port 58 nsew signal input
flabel metal3 s -960 32316 480 32556 0 FreeSans 960 0 0 0 io_in[37]
port 59 nsew signal input
flabel metal3 s 583520 125884 584960 126124 0 FreeSans 960 0 0 0 io_in[3]
port 60 nsew signal input
flabel metal3 s 583520 165732 584960 165972 0 FreeSans 960 0 0 0 io_in[4]
port 61 nsew signal input
flabel metal3 s 583520 205580 584960 205820 0 FreeSans 960 0 0 0 io_in[5]
port 62 nsew signal input
flabel metal3 s 583520 245428 584960 245668 0 FreeSans 960 0 0 0 io_in[6]
port 63 nsew signal input
flabel metal3 s 583520 298604 584960 298844 0 FreeSans 960 0 0 0 io_in[7]
port 64 nsew signal input
flabel metal3 s 583520 351780 584960 352020 0 FreeSans 960 0 0 0 io_in[8]
port 65 nsew signal input
flabel metal3 s 583520 404820 584960 405060 0 FreeSans 960 0 0 0 io_in[9]
port 66 nsew signal input
flabel metal3 s 583520 32996 584960 33236 0 FreeSans 960 0 0 0 io_oeb[0]
port 67 nsew signal tristate
flabel metal3 s 583520 484516 584960 484756 0 FreeSans 960 0 0 0 io_oeb[10]
port 68 nsew signal tristate
flabel metal3 s 583520 537692 584960 537932 0 FreeSans 960 0 0 0 io_oeb[11]
port 69 nsew signal tristate
flabel metal3 s 583520 590868 584960 591108 0 FreeSans 960 0 0 0 io_oeb[12]
port 70 nsew signal tristate
flabel metal3 s 583520 643908 584960 644148 0 FreeSans 960 0 0 0 io_oeb[13]
port 71 nsew signal tristate
flabel metal3 s 583520 697084 584960 697324 0 FreeSans 960 0 0 0 io_oeb[14]
port 72 nsew signal tristate
flabel metal2 s 527150 703520 527262 704960 0 FreeSans 448 90 0 0 io_oeb[15]
port 73 nsew signal tristate
flabel metal2 s 462290 703520 462402 704960 0 FreeSans 448 90 0 0 io_oeb[16]
port 74 nsew signal tristate
flabel metal2 s 397430 703520 397542 704960 0 FreeSans 448 90 0 0 io_oeb[17]
port 75 nsew signal tristate
flabel metal2 s 332478 703520 332590 704960 0 FreeSans 448 90 0 0 io_oeb[18]
port 76 nsew signal tristate
flabel metal2 s 267618 703520 267730 704960 0 FreeSans 448 90 0 0 io_oeb[19]
port 77 nsew signal tristate
flabel metal3 s 583520 72844 584960 73084 0 FreeSans 960 0 0 0 io_oeb[1]
port 78 nsew signal tristate
flabel metal2 s 202758 703520 202870 704960 0 FreeSans 448 90 0 0 io_oeb[20]
port 79 nsew signal tristate
flabel metal2 s 137806 703520 137918 704960 0 FreeSans 448 90 0 0 io_oeb[21]
port 80 nsew signal tristate
flabel metal2 s 72946 703520 73058 704960 0 FreeSans 448 90 0 0 io_oeb[22]
port 81 nsew signal tristate
flabel metal2 s 8086 703520 8198 704960 0 FreeSans 448 90 0 0 io_oeb[23]
port 82 nsew signal tristate
flabel metal3 s -960 658052 480 658292 0 FreeSans 960 0 0 0 io_oeb[24]
port 83 nsew signal tristate
flabel metal3 s -960 605964 480 606204 0 FreeSans 960 0 0 0 io_oeb[25]
port 84 nsew signal tristate
flabel metal3 s -960 553740 480 553980 0 FreeSans 960 0 0 0 io_oeb[26]
port 85 nsew signal tristate
flabel metal3 s -960 501652 480 501892 0 FreeSans 960 0 0 0 io_oeb[27]
port 86 nsew signal tristate
flabel metal3 s -960 449428 480 449668 0 FreeSans 960 0 0 0 io_oeb[28]
port 87 nsew signal tristate
flabel metal3 s -960 397340 480 397580 0 FreeSans 960 0 0 0 io_oeb[29]
port 88 nsew signal tristate
flabel metal3 s 583520 112692 584960 112932 0 FreeSans 960 0 0 0 io_oeb[2]
port 89 nsew signal tristate
flabel metal3 s -960 345252 480 345492 0 FreeSans 960 0 0 0 io_oeb[30]
port 90 nsew signal tristate
flabel metal3 s -960 293028 480 293268 0 FreeSans 960 0 0 0 io_oeb[31]
port 91 nsew signal tristate
flabel metal3 s -960 240940 480 241180 0 FreeSans 960 0 0 0 io_oeb[32]
port 92 nsew signal tristate
flabel metal3 s -960 188716 480 188956 0 FreeSans 960 0 0 0 io_oeb[33]
port 93 nsew signal tristate
flabel metal3 s -960 136628 480 136868 0 FreeSans 960 0 0 0 io_oeb[34]
port 94 nsew signal tristate
flabel metal3 s -960 84540 480 84780 0 FreeSans 960 0 0 0 io_oeb[35]
port 95 nsew signal tristate
flabel metal3 s -960 45372 480 45612 0 FreeSans 960 0 0 0 io_oeb[36]
port 96 nsew signal tristate
flabel metal3 s -960 6340 480 6580 0 FreeSans 960 0 0 0 io_oeb[37]
port 97 nsew signal tristate
flabel metal3 s 583520 152540 584960 152780 0 FreeSans 960 0 0 0 io_oeb[3]
port 98 nsew signal tristate
flabel metal3 s 583520 192388 584960 192628 0 FreeSans 960 0 0 0 io_oeb[4]
port 99 nsew signal tristate
flabel metal3 s 583520 232236 584960 232476 0 FreeSans 960 0 0 0 io_oeb[5]
port 100 nsew signal tristate
flabel metal3 s 583520 272084 584960 272324 0 FreeSans 960 0 0 0 io_oeb[6]
port 101 nsew signal tristate
flabel metal3 s 583520 325124 584960 325364 0 FreeSans 960 0 0 0 io_oeb[7]
port 102 nsew signal tristate
flabel metal3 s 583520 378300 584960 378540 0 FreeSans 960 0 0 0 io_oeb[8]
port 103 nsew signal tristate
flabel metal3 s 583520 431476 584960 431716 0 FreeSans 960 0 0 0 io_oeb[9]
port 104 nsew signal tristate
flabel metal3 s 583520 19668 584960 19908 0 FreeSans 960 0 0 0 io_out[0]
port 105 nsew signal tristate
flabel metal3 s 583520 471324 584960 471564 0 FreeSans 960 0 0 0 io_out[10]
port 106 nsew signal tristate
flabel metal3 s 583520 524364 584960 524604 0 FreeSans 960 0 0 0 io_out[11]
port 107 nsew signal tristate
flabel metal3 s 583520 577540 584960 577780 0 FreeSans 960 0 0 0 io_out[12]
port 108 nsew signal tristate
flabel metal3 s 583520 630716 584960 630956 0 FreeSans 960 0 0 0 io_out[13]
port 109 nsew signal tristate
flabel metal3 s 583520 683756 584960 683996 0 FreeSans 960 0 0 0 io_out[14]
port 110 nsew signal tristate
flabel metal2 s 543434 703520 543546 704960 0 FreeSans 448 90 0 0 io_out[15]
port 111 nsew signal tristate
flabel metal2 s 478482 703520 478594 704960 0 FreeSans 448 90 0 0 io_out[16]
port 112 nsew signal tristate
flabel metal2 s 413622 703520 413734 704960 0 FreeSans 448 90 0 0 io_out[17]
port 113 nsew signal tristate
flabel metal2 s 348762 703520 348874 704960 0 FreeSans 448 90 0 0 io_out[18]
port 114 nsew signal tristate
flabel metal2 s 283810 703520 283922 704960 0 FreeSans 448 90 0 0 io_out[19]
port 115 nsew signal tristate
flabel metal3 s 583520 59516 584960 59756 0 FreeSans 960 0 0 0 io_out[1]
port 116 nsew signal tristate
flabel metal2 s 218950 703520 219062 704960 0 FreeSans 448 90 0 0 io_out[20]
port 117 nsew signal tristate
flabel metal2 s 154090 703520 154202 704960 0 FreeSans 448 90 0 0 io_out[21]
port 118 nsew signal tristate
flabel metal2 s 89138 703520 89250 704960 0 FreeSans 448 90 0 0 io_out[22]
port 119 nsew signal tristate
flabel metal2 s 24278 703520 24390 704960 0 FreeSans 448 90 0 0 io_out[23]
port 120 nsew signal tristate
flabel metal3 s -960 671108 480 671348 0 FreeSans 960 0 0 0 io_out[24]
port 121 nsew signal tristate
flabel metal3 s -960 619020 480 619260 0 FreeSans 960 0 0 0 io_out[25]
port 122 nsew signal tristate
flabel metal3 s -960 566796 480 567036 0 FreeSans 960 0 0 0 io_out[26]
port 123 nsew signal tristate
flabel metal3 s -960 514708 480 514948 0 FreeSans 960 0 0 0 io_out[27]
port 124 nsew signal tristate
flabel metal3 s -960 462484 480 462724 0 FreeSans 960 0 0 0 io_out[28]
port 125 nsew signal tristate
flabel metal3 s -960 410396 480 410636 0 FreeSans 960 0 0 0 io_out[29]
port 126 nsew signal tristate
flabel metal3 s 583520 99364 584960 99604 0 FreeSans 960 0 0 0 io_out[2]
port 127 nsew signal tristate
flabel metal3 s -960 358308 480 358548 0 FreeSans 960 0 0 0 io_out[30]
port 128 nsew signal tristate
flabel metal3 s -960 306084 480 306324 0 FreeSans 960 0 0 0 io_out[31]
port 129 nsew signal tristate
flabel metal3 s -960 253996 480 254236 0 FreeSans 960 0 0 0 io_out[32]
port 130 nsew signal tristate
flabel metal3 s -960 201772 480 202012 0 FreeSans 960 0 0 0 io_out[33]
port 131 nsew signal tristate
flabel metal3 s -960 149684 480 149924 0 FreeSans 960 0 0 0 io_out[34]
port 132 nsew signal tristate
flabel metal3 s -960 97460 480 97700 0 FreeSans 960 0 0 0 io_out[35]
port 133 nsew signal tristate
flabel metal3 s -960 58428 480 58668 0 FreeSans 960 0 0 0 io_out[36]
port 134 nsew signal tristate
flabel metal3 s -960 19260 480 19500 0 FreeSans 960 0 0 0 io_out[37]
port 135 nsew signal tristate
flabel metal3 s 583520 139212 584960 139452 0 FreeSans 960 0 0 0 io_out[3]
port 136 nsew signal tristate
flabel metal3 s 583520 179060 584960 179300 0 FreeSans 960 0 0 0 io_out[4]
port 137 nsew signal tristate
flabel metal3 s 583520 218908 584960 219148 0 FreeSans 960 0 0 0 io_out[5]
port 138 nsew signal tristate
flabel metal3 s 583520 258756 584960 258996 0 FreeSans 960 0 0 0 io_out[6]
port 139 nsew signal tristate
flabel metal3 s 583520 311932 584960 312172 0 FreeSans 960 0 0 0 io_out[7]
port 140 nsew signal tristate
flabel metal3 s 583520 364972 584960 365212 0 FreeSans 960 0 0 0 io_out[8]
port 141 nsew signal tristate
flabel metal3 s 583520 418148 584960 418388 0 FreeSans 960 0 0 0 io_out[9]
port 142 nsew signal tristate
flabel metal2 s 125846 -960 125958 480 0 FreeSans 448 90 0 0 la_data_in[0]
port 143 nsew signal input
flabel metal2 s 480506 -960 480618 480 0 FreeSans 448 90 0 0 la_data_in[100]
port 144 nsew signal input
flabel metal2 s 484002 -960 484114 480 0 FreeSans 448 90 0 0 la_data_in[101]
port 145 nsew signal input
flabel metal2 s 487590 -960 487702 480 0 FreeSans 448 90 0 0 la_data_in[102]
port 146 nsew signal input
flabel metal2 s 491086 -960 491198 480 0 FreeSans 448 90 0 0 la_data_in[103]
port 147 nsew signal input
flabel metal2 s 494674 -960 494786 480 0 FreeSans 448 90 0 0 la_data_in[104]
port 148 nsew signal input
flabel metal2 s 498170 -960 498282 480 0 FreeSans 448 90 0 0 la_data_in[105]
port 149 nsew signal input
flabel metal2 s 501758 -960 501870 480 0 FreeSans 448 90 0 0 la_data_in[106]
port 150 nsew signal input
flabel metal2 s 505346 -960 505458 480 0 FreeSans 448 90 0 0 la_data_in[107]
port 151 nsew signal input
flabel metal2 s 508842 -960 508954 480 0 FreeSans 448 90 0 0 la_data_in[108]
port 152 nsew signal input
flabel metal2 s 512430 -960 512542 480 0 FreeSans 448 90 0 0 la_data_in[109]
port 153 nsew signal input
flabel metal2 s 161266 -960 161378 480 0 FreeSans 448 90 0 0 la_data_in[10]
port 154 nsew signal input
flabel metal2 s 515926 -960 516038 480 0 FreeSans 448 90 0 0 la_data_in[110]
port 155 nsew signal input
flabel metal2 s 519514 -960 519626 480 0 FreeSans 448 90 0 0 la_data_in[111]
port 156 nsew signal input
flabel metal2 s 523010 -960 523122 480 0 FreeSans 448 90 0 0 la_data_in[112]
port 157 nsew signal input
flabel metal2 s 526598 -960 526710 480 0 FreeSans 448 90 0 0 la_data_in[113]
port 158 nsew signal input
flabel metal2 s 530094 -960 530206 480 0 FreeSans 448 90 0 0 la_data_in[114]
port 159 nsew signal input
flabel metal2 s 533682 -960 533794 480 0 FreeSans 448 90 0 0 la_data_in[115]
port 160 nsew signal input
flabel metal2 s 537178 -960 537290 480 0 FreeSans 448 90 0 0 la_data_in[116]
port 161 nsew signal input
flabel metal2 s 540766 -960 540878 480 0 FreeSans 448 90 0 0 la_data_in[117]
port 162 nsew signal input
flabel metal2 s 544354 -960 544466 480 0 FreeSans 448 90 0 0 la_data_in[118]
port 163 nsew signal input
flabel metal2 s 547850 -960 547962 480 0 FreeSans 448 90 0 0 la_data_in[119]
port 164 nsew signal input
flabel metal2 s 164854 -960 164966 480 0 FreeSans 448 90 0 0 la_data_in[11]
port 165 nsew signal input
flabel metal2 s 551438 -960 551550 480 0 FreeSans 448 90 0 0 la_data_in[120]
port 166 nsew signal input
flabel metal2 s 554934 -960 555046 480 0 FreeSans 448 90 0 0 la_data_in[121]
port 167 nsew signal input
flabel metal2 s 558522 -960 558634 480 0 FreeSans 448 90 0 0 la_data_in[122]
port 168 nsew signal input
flabel metal2 s 562018 -960 562130 480 0 FreeSans 448 90 0 0 la_data_in[123]
port 169 nsew signal input
flabel metal2 s 565606 -960 565718 480 0 FreeSans 448 90 0 0 la_data_in[124]
port 170 nsew signal input
flabel metal2 s 569102 -960 569214 480 0 FreeSans 448 90 0 0 la_data_in[125]
port 171 nsew signal input
flabel metal2 s 572690 -960 572802 480 0 FreeSans 448 90 0 0 la_data_in[126]
port 172 nsew signal input
flabel metal2 s 576278 -960 576390 480 0 FreeSans 448 90 0 0 la_data_in[127]
port 173 nsew signal input
flabel metal2 s 168350 -960 168462 480 0 FreeSans 448 90 0 0 la_data_in[12]
port 174 nsew signal input
flabel metal2 s 171938 -960 172050 480 0 FreeSans 448 90 0 0 la_data_in[13]
port 175 nsew signal input
flabel metal2 s 175434 -960 175546 480 0 FreeSans 448 90 0 0 la_data_in[14]
port 176 nsew signal input
flabel metal2 s 179022 -960 179134 480 0 FreeSans 448 90 0 0 la_data_in[15]
port 177 nsew signal input
flabel metal2 s 182518 -960 182630 480 0 FreeSans 448 90 0 0 la_data_in[16]
port 178 nsew signal input
flabel metal2 s 186106 -960 186218 480 0 FreeSans 448 90 0 0 la_data_in[17]
port 179 nsew signal input
flabel metal2 s 189694 -960 189806 480 0 FreeSans 448 90 0 0 la_data_in[18]
port 180 nsew signal input
flabel metal2 s 193190 -960 193302 480 0 FreeSans 448 90 0 0 la_data_in[19]
port 181 nsew signal input
flabel metal2 s 129342 -960 129454 480 0 FreeSans 448 90 0 0 la_data_in[1]
port 182 nsew signal input
flabel metal2 s 196778 -960 196890 480 0 FreeSans 448 90 0 0 la_data_in[20]
port 183 nsew signal input
flabel metal2 s 200274 -960 200386 480 0 FreeSans 448 90 0 0 la_data_in[21]
port 184 nsew signal input
flabel metal2 s 203862 -960 203974 480 0 FreeSans 448 90 0 0 la_data_in[22]
port 185 nsew signal input
flabel metal2 s 207358 -960 207470 480 0 FreeSans 448 90 0 0 la_data_in[23]
port 186 nsew signal input
flabel metal2 s 210946 -960 211058 480 0 FreeSans 448 90 0 0 la_data_in[24]
port 187 nsew signal input
flabel metal2 s 214442 -960 214554 480 0 FreeSans 448 90 0 0 la_data_in[25]
port 188 nsew signal input
flabel metal2 s 218030 -960 218142 480 0 FreeSans 448 90 0 0 la_data_in[26]
port 189 nsew signal input
flabel metal2 s 221526 -960 221638 480 0 FreeSans 448 90 0 0 la_data_in[27]
port 190 nsew signal input
flabel metal2 s 225114 -960 225226 480 0 FreeSans 448 90 0 0 la_data_in[28]
port 191 nsew signal input
flabel metal2 s 228702 -960 228814 480 0 FreeSans 448 90 0 0 la_data_in[29]
port 192 nsew signal input
flabel metal2 s 132930 -960 133042 480 0 FreeSans 448 90 0 0 la_data_in[2]
port 193 nsew signal input
flabel metal2 s 232198 -960 232310 480 0 FreeSans 448 90 0 0 la_data_in[30]
port 194 nsew signal input
flabel metal2 s 235786 -960 235898 480 0 FreeSans 448 90 0 0 la_data_in[31]
port 195 nsew signal input
flabel metal2 s 239282 -960 239394 480 0 FreeSans 448 90 0 0 la_data_in[32]
port 196 nsew signal input
flabel metal2 s 242870 -960 242982 480 0 FreeSans 448 90 0 0 la_data_in[33]
port 197 nsew signal input
flabel metal2 s 246366 -960 246478 480 0 FreeSans 448 90 0 0 la_data_in[34]
port 198 nsew signal input
flabel metal2 s 249954 -960 250066 480 0 FreeSans 448 90 0 0 la_data_in[35]
port 199 nsew signal input
flabel metal2 s 253450 -960 253562 480 0 FreeSans 448 90 0 0 la_data_in[36]
port 200 nsew signal input
flabel metal2 s 257038 -960 257150 480 0 FreeSans 448 90 0 0 la_data_in[37]
port 201 nsew signal input
flabel metal2 s 260626 -960 260738 480 0 FreeSans 448 90 0 0 la_data_in[38]
port 202 nsew signal input
flabel metal2 s 264122 -960 264234 480 0 FreeSans 448 90 0 0 la_data_in[39]
port 203 nsew signal input
flabel metal2 s 136426 -960 136538 480 0 FreeSans 448 90 0 0 la_data_in[3]
port 204 nsew signal input
flabel metal2 s 267710 -960 267822 480 0 FreeSans 448 90 0 0 la_data_in[40]
port 205 nsew signal input
flabel metal2 s 271206 -960 271318 480 0 FreeSans 448 90 0 0 la_data_in[41]
port 206 nsew signal input
flabel metal2 s 274794 -960 274906 480 0 FreeSans 448 90 0 0 la_data_in[42]
port 207 nsew signal input
flabel metal2 s 278290 -960 278402 480 0 FreeSans 448 90 0 0 la_data_in[43]
port 208 nsew signal input
flabel metal2 s 281878 -960 281990 480 0 FreeSans 448 90 0 0 la_data_in[44]
port 209 nsew signal input
flabel metal2 s 285374 -960 285486 480 0 FreeSans 448 90 0 0 la_data_in[45]
port 210 nsew signal input
flabel metal2 s 288962 -960 289074 480 0 FreeSans 448 90 0 0 la_data_in[46]
port 211 nsew signal input
flabel metal2 s 292550 -960 292662 480 0 FreeSans 448 90 0 0 la_data_in[47]
port 212 nsew signal input
flabel metal2 s 296046 -960 296158 480 0 FreeSans 448 90 0 0 la_data_in[48]
port 213 nsew signal input
flabel metal2 s 299634 -960 299746 480 0 FreeSans 448 90 0 0 la_data_in[49]
port 214 nsew signal input
flabel metal2 s 140014 -960 140126 480 0 FreeSans 448 90 0 0 la_data_in[4]
port 215 nsew signal input
flabel metal2 s 303130 -960 303242 480 0 FreeSans 448 90 0 0 la_data_in[50]
port 216 nsew signal input
flabel metal2 s 306718 -960 306830 480 0 FreeSans 448 90 0 0 la_data_in[51]
port 217 nsew signal input
flabel metal2 s 310214 -960 310326 480 0 FreeSans 448 90 0 0 la_data_in[52]
port 218 nsew signal input
flabel metal2 s 313802 -960 313914 480 0 FreeSans 448 90 0 0 la_data_in[53]
port 219 nsew signal input
flabel metal2 s 317298 -960 317410 480 0 FreeSans 448 90 0 0 la_data_in[54]
port 220 nsew signal input
flabel metal2 s 320886 -960 320998 480 0 FreeSans 448 90 0 0 la_data_in[55]
port 221 nsew signal input
flabel metal2 s 324382 -960 324494 480 0 FreeSans 448 90 0 0 la_data_in[56]
port 222 nsew signal input
flabel metal2 s 327970 -960 328082 480 0 FreeSans 448 90 0 0 la_data_in[57]
port 223 nsew signal input
flabel metal2 s 331558 -960 331670 480 0 FreeSans 448 90 0 0 la_data_in[58]
port 224 nsew signal input
flabel metal2 s 335054 -960 335166 480 0 FreeSans 448 90 0 0 la_data_in[59]
port 225 nsew signal input
flabel metal2 s 143510 -960 143622 480 0 FreeSans 448 90 0 0 la_data_in[5]
port 226 nsew signal input
flabel metal2 s 338642 -960 338754 480 0 FreeSans 448 90 0 0 la_data_in[60]
port 227 nsew signal input
flabel metal2 s 342138 -960 342250 480 0 FreeSans 448 90 0 0 la_data_in[61]
port 228 nsew signal input
flabel metal2 s 345726 -960 345838 480 0 FreeSans 448 90 0 0 la_data_in[62]
port 229 nsew signal input
flabel metal2 s 349222 -960 349334 480 0 FreeSans 448 90 0 0 la_data_in[63]
port 230 nsew signal input
flabel metal2 s 352810 -960 352922 480 0 FreeSans 448 90 0 0 la_data_in[64]
port 231 nsew signal input
flabel metal2 s 356306 -960 356418 480 0 FreeSans 448 90 0 0 la_data_in[65]
port 232 nsew signal input
flabel metal2 s 359894 -960 360006 480 0 FreeSans 448 90 0 0 la_data_in[66]
port 233 nsew signal input
flabel metal2 s 363482 -960 363594 480 0 FreeSans 448 90 0 0 la_data_in[67]
port 234 nsew signal input
flabel metal2 s 366978 -960 367090 480 0 FreeSans 448 90 0 0 la_data_in[68]
port 235 nsew signal input
flabel metal2 s 370566 -960 370678 480 0 FreeSans 448 90 0 0 la_data_in[69]
port 236 nsew signal input
flabel metal2 s 147098 -960 147210 480 0 FreeSans 448 90 0 0 la_data_in[6]
port 237 nsew signal input
flabel metal2 s 374062 -960 374174 480 0 FreeSans 448 90 0 0 la_data_in[70]
port 238 nsew signal input
flabel metal2 s 377650 -960 377762 480 0 FreeSans 448 90 0 0 la_data_in[71]
port 239 nsew signal input
flabel metal2 s 381146 -960 381258 480 0 FreeSans 448 90 0 0 la_data_in[72]
port 240 nsew signal input
flabel metal2 s 384734 -960 384846 480 0 FreeSans 448 90 0 0 la_data_in[73]
port 241 nsew signal input
flabel metal2 s 388230 -960 388342 480 0 FreeSans 448 90 0 0 la_data_in[74]
port 242 nsew signal input
flabel metal2 s 391818 -960 391930 480 0 FreeSans 448 90 0 0 la_data_in[75]
port 243 nsew signal input
flabel metal2 s 395314 -960 395426 480 0 FreeSans 448 90 0 0 la_data_in[76]
port 244 nsew signal input
flabel metal2 s 398902 -960 399014 480 0 FreeSans 448 90 0 0 la_data_in[77]
port 245 nsew signal input
flabel metal2 s 402490 -960 402602 480 0 FreeSans 448 90 0 0 la_data_in[78]
port 246 nsew signal input
flabel metal2 s 405986 -960 406098 480 0 FreeSans 448 90 0 0 la_data_in[79]
port 247 nsew signal input
flabel metal2 s 150594 -960 150706 480 0 FreeSans 448 90 0 0 la_data_in[7]
port 248 nsew signal input
flabel metal2 s 409574 -960 409686 480 0 FreeSans 448 90 0 0 la_data_in[80]
port 249 nsew signal input
flabel metal2 s 413070 -960 413182 480 0 FreeSans 448 90 0 0 la_data_in[81]
port 250 nsew signal input
flabel metal2 s 416658 -960 416770 480 0 FreeSans 448 90 0 0 la_data_in[82]
port 251 nsew signal input
flabel metal2 s 420154 -960 420266 480 0 FreeSans 448 90 0 0 la_data_in[83]
port 252 nsew signal input
flabel metal2 s 423742 -960 423854 480 0 FreeSans 448 90 0 0 la_data_in[84]
port 253 nsew signal input
flabel metal2 s 427238 -960 427350 480 0 FreeSans 448 90 0 0 la_data_in[85]
port 254 nsew signal input
flabel metal2 s 430826 -960 430938 480 0 FreeSans 448 90 0 0 la_data_in[86]
port 255 nsew signal input
flabel metal2 s 434414 -960 434526 480 0 FreeSans 448 90 0 0 la_data_in[87]
port 256 nsew signal input
flabel metal2 s 437910 -960 438022 480 0 FreeSans 448 90 0 0 la_data_in[88]
port 257 nsew signal input
flabel metal2 s 441498 -960 441610 480 0 FreeSans 448 90 0 0 la_data_in[89]
port 258 nsew signal input
flabel metal2 s 154182 -960 154294 480 0 FreeSans 448 90 0 0 la_data_in[8]
port 259 nsew signal input
flabel metal2 s 444994 -960 445106 480 0 FreeSans 448 90 0 0 la_data_in[90]
port 260 nsew signal input
flabel metal2 s 448582 -960 448694 480 0 FreeSans 448 90 0 0 la_data_in[91]
port 261 nsew signal input
flabel metal2 s 452078 -960 452190 480 0 FreeSans 448 90 0 0 la_data_in[92]
port 262 nsew signal input
flabel metal2 s 455666 -960 455778 480 0 FreeSans 448 90 0 0 la_data_in[93]
port 263 nsew signal input
flabel metal2 s 459162 -960 459274 480 0 FreeSans 448 90 0 0 la_data_in[94]
port 264 nsew signal input
flabel metal2 s 462750 -960 462862 480 0 FreeSans 448 90 0 0 la_data_in[95]
port 265 nsew signal input
flabel metal2 s 466246 -960 466358 480 0 FreeSans 448 90 0 0 la_data_in[96]
port 266 nsew signal input
flabel metal2 s 469834 -960 469946 480 0 FreeSans 448 90 0 0 la_data_in[97]
port 267 nsew signal input
flabel metal2 s 473422 -960 473534 480 0 FreeSans 448 90 0 0 la_data_in[98]
port 268 nsew signal input
flabel metal2 s 476918 -960 477030 480 0 FreeSans 448 90 0 0 la_data_in[99]
port 269 nsew signal input
flabel metal2 s 157770 -960 157882 480 0 FreeSans 448 90 0 0 la_data_in[9]
port 270 nsew signal input
flabel metal2 s 126950 -960 127062 480 0 FreeSans 448 90 0 0 la_data_out[0]
port 271 nsew signal tristate
flabel metal2 s 481702 -960 481814 480 0 FreeSans 448 90 0 0 la_data_out[100]
port 272 nsew signal tristate
flabel metal2 s 485198 -960 485310 480 0 FreeSans 448 90 0 0 la_data_out[101]
port 273 nsew signal tristate
flabel metal2 s 488786 -960 488898 480 0 FreeSans 448 90 0 0 la_data_out[102]
port 274 nsew signal tristate
flabel metal2 s 492282 -960 492394 480 0 FreeSans 448 90 0 0 la_data_out[103]
port 275 nsew signal tristate
flabel metal2 s 495870 -960 495982 480 0 FreeSans 448 90 0 0 la_data_out[104]
port 276 nsew signal tristate
flabel metal2 s 499366 -960 499478 480 0 FreeSans 448 90 0 0 la_data_out[105]
port 277 nsew signal tristate
flabel metal2 s 502954 -960 503066 480 0 FreeSans 448 90 0 0 la_data_out[106]
port 278 nsew signal tristate
flabel metal2 s 506450 -960 506562 480 0 FreeSans 448 90 0 0 la_data_out[107]
port 279 nsew signal tristate
flabel metal2 s 510038 -960 510150 480 0 FreeSans 448 90 0 0 la_data_out[108]
port 280 nsew signal tristate
flabel metal2 s 513534 -960 513646 480 0 FreeSans 448 90 0 0 la_data_out[109]
port 281 nsew signal tristate
flabel metal2 s 162462 -960 162574 480 0 FreeSans 448 90 0 0 la_data_out[10]
port 282 nsew signal tristate
flabel metal2 s 517122 -960 517234 480 0 FreeSans 448 90 0 0 la_data_out[110]
port 283 nsew signal tristate
flabel metal2 s 520710 -960 520822 480 0 FreeSans 448 90 0 0 la_data_out[111]
port 284 nsew signal tristate
flabel metal2 s 524206 -960 524318 480 0 FreeSans 448 90 0 0 la_data_out[112]
port 285 nsew signal tristate
flabel metal2 s 527794 -960 527906 480 0 FreeSans 448 90 0 0 la_data_out[113]
port 286 nsew signal tristate
flabel metal2 s 531290 -960 531402 480 0 FreeSans 448 90 0 0 la_data_out[114]
port 287 nsew signal tristate
flabel metal2 s 534878 -960 534990 480 0 FreeSans 448 90 0 0 la_data_out[115]
port 288 nsew signal tristate
flabel metal2 s 538374 -960 538486 480 0 FreeSans 448 90 0 0 la_data_out[116]
port 289 nsew signal tristate
flabel metal2 s 541962 -960 542074 480 0 FreeSans 448 90 0 0 la_data_out[117]
port 290 nsew signal tristate
flabel metal2 s 545458 -960 545570 480 0 FreeSans 448 90 0 0 la_data_out[118]
port 291 nsew signal tristate
flabel metal2 s 549046 -960 549158 480 0 FreeSans 448 90 0 0 la_data_out[119]
port 292 nsew signal tristate
flabel metal2 s 166050 -960 166162 480 0 FreeSans 448 90 0 0 la_data_out[11]
port 293 nsew signal tristate
flabel metal2 s 552634 -960 552746 480 0 FreeSans 448 90 0 0 la_data_out[120]
port 294 nsew signal tristate
flabel metal2 s 556130 -960 556242 480 0 FreeSans 448 90 0 0 la_data_out[121]
port 295 nsew signal tristate
flabel metal2 s 559718 -960 559830 480 0 FreeSans 448 90 0 0 la_data_out[122]
port 296 nsew signal tristate
flabel metal2 s 563214 -960 563326 480 0 FreeSans 448 90 0 0 la_data_out[123]
port 297 nsew signal tristate
flabel metal2 s 566802 -960 566914 480 0 FreeSans 448 90 0 0 la_data_out[124]
port 298 nsew signal tristate
flabel metal2 s 570298 -960 570410 480 0 FreeSans 448 90 0 0 la_data_out[125]
port 299 nsew signal tristate
flabel metal2 s 573886 -960 573998 480 0 FreeSans 448 90 0 0 la_data_out[126]
port 300 nsew signal tristate
flabel metal2 s 577382 -960 577494 480 0 FreeSans 448 90 0 0 la_data_out[127]
port 301 nsew signal tristate
flabel metal2 s 169546 -960 169658 480 0 FreeSans 448 90 0 0 la_data_out[12]
port 302 nsew signal tristate
flabel metal2 s 173134 -960 173246 480 0 FreeSans 448 90 0 0 la_data_out[13]
port 303 nsew signal tristate
flabel metal2 s 176630 -960 176742 480 0 FreeSans 448 90 0 0 la_data_out[14]
port 304 nsew signal tristate
flabel metal2 s 180218 -960 180330 480 0 FreeSans 448 90 0 0 la_data_out[15]
port 305 nsew signal tristate
flabel metal2 s 183714 -960 183826 480 0 FreeSans 448 90 0 0 la_data_out[16]
port 306 nsew signal tristate
flabel metal2 s 187302 -960 187414 480 0 FreeSans 448 90 0 0 la_data_out[17]
port 307 nsew signal tristate
flabel metal2 s 190798 -960 190910 480 0 FreeSans 448 90 0 0 la_data_out[18]
port 308 nsew signal tristate
flabel metal2 s 194386 -960 194498 480 0 FreeSans 448 90 0 0 la_data_out[19]
port 309 nsew signal tristate
flabel metal2 s 130538 -960 130650 480 0 FreeSans 448 90 0 0 la_data_out[1]
port 310 nsew signal tristate
flabel metal2 s 197882 -960 197994 480 0 FreeSans 448 90 0 0 la_data_out[20]
port 311 nsew signal tristate
flabel metal2 s 201470 -960 201582 480 0 FreeSans 448 90 0 0 la_data_out[21]
port 312 nsew signal tristate
flabel metal2 s 205058 -960 205170 480 0 FreeSans 448 90 0 0 la_data_out[22]
port 313 nsew signal tristate
flabel metal2 s 208554 -960 208666 480 0 FreeSans 448 90 0 0 la_data_out[23]
port 314 nsew signal tristate
flabel metal2 s 212142 -960 212254 480 0 FreeSans 448 90 0 0 la_data_out[24]
port 315 nsew signal tristate
flabel metal2 s 215638 -960 215750 480 0 FreeSans 448 90 0 0 la_data_out[25]
port 316 nsew signal tristate
flabel metal2 s 219226 -960 219338 480 0 FreeSans 448 90 0 0 la_data_out[26]
port 317 nsew signal tristate
flabel metal2 s 222722 -960 222834 480 0 FreeSans 448 90 0 0 la_data_out[27]
port 318 nsew signal tristate
flabel metal2 s 226310 -960 226422 480 0 FreeSans 448 90 0 0 la_data_out[28]
port 319 nsew signal tristate
flabel metal2 s 229806 -960 229918 480 0 FreeSans 448 90 0 0 la_data_out[29]
port 320 nsew signal tristate
flabel metal2 s 134126 -960 134238 480 0 FreeSans 448 90 0 0 la_data_out[2]
port 321 nsew signal tristate
flabel metal2 s 233394 -960 233506 480 0 FreeSans 448 90 0 0 la_data_out[30]
port 322 nsew signal tristate
flabel metal2 s 236982 -960 237094 480 0 FreeSans 448 90 0 0 la_data_out[31]
port 323 nsew signal tristate
flabel metal2 s 240478 -960 240590 480 0 FreeSans 448 90 0 0 la_data_out[32]
port 324 nsew signal tristate
flabel metal2 s 244066 -960 244178 480 0 FreeSans 448 90 0 0 la_data_out[33]
port 325 nsew signal tristate
flabel metal2 s 247562 -960 247674 480 0 FreeSans 448 90 0 0 la_data_out[34]
port 326 nsew signal tristate
flabel metal2 s 251150 -960 251262 480 0 FreeSans 448 90 0 0 la_data_out[35]
port 327 nsew signal tristate
flabel metal2 s 254646 -960 254758 480 0 FreeSans 448 90 0 0 la_data_out[36]
port 328 nsew signal tristate
flabel metal2 s 258234 -960 258346 480 0 FreeSans 448 90 0 0 la_data_out[37]
port 329 nsew signal tristate
flabel metal2 s 261730 -960 261842 480 0 FreeSans 448 90 0 0 la_data_out[38]
port 330 nsew signal tristate
flabel metal2 s 265318 -960 265430 480 0 FreeSans 448 90 0 0 la_data_out[39]
port 331 nsew signal tristate
flabel metal2 s 137622 -960 137734 480 0 FreeSans 448 90 0 0 la_data_out[3]
port 332 nsew signal tristate
flabel metal2 s 268814 -960 268926 480 0 FreeSans 448 90 0 0 la_data_out[40]
port 333 nsew signal tristate
flabel metal2 s 272402 -960 272514 480 0 FreeSans 448 90 0 0 la_data_out[41]
port 334 nsew signal tristate
flabel metal2 s 275990 -960 276102 480 0 FreeSans 448 90 0 0 la_data_out[42]
port 335 nsew signal tristate
flabel metal2 s 279486 -960 279598 480 0 FreeSans 448 90 0 0 la_data_out[43]
port 336 nsew signal tristate
flabel metal2 s 283074 -960 283186 480 0 FreeSans 448 90 0 0 la_data_out[44]
port 337 nsew signal tristate
flabel metal2 s 286570 -960 286682 480 0 FreeSans 448 90 0 0 la_data_out[45]
port 338 nsew signal tristate
flabel metal2 s 290158 -960 290270 480 0 FreeSans 448 90 0 0 la_data_out[46]
port 339 nsew signal tristate
flabel metal2 s 293654 -960 293766 480 0 FreeSans 448 90 0 0 la_data_out[47]
port 340 nsew signal tristate
flabel metal2 s 297242 -960 297354 480 0 FreeSans 448 90 0 0 la_data_out[48]
port 341 nsew signal tristate
flabel metal2 s 300738 -960 300850 480 0 FreeSans 448 90 0 0 la_data_out[49]
port 342 nsew signal tristate
flabel metal2 s 141210 -960 141322 480 0 FreeSans 448 90 0 0 la_data_out[4]
port 343 nsew signal tristate
flabel metal2 s 304326 -960 304438 480 0 FreeSans 448 90 0 0 la_data_out[50]
port 344 nsew signal tristate
flabel metal2 s 307914 -960 308026 480 0 FreeSans 448 90 0 0 la_data_out[51]
port 345 nsew signal tristate
flabel metal2 s 311410 -960 311522 480 0 FreeSans 448 90 0 0 la_data_out[52]
port 346 nsew signal tristate
flabel metal2 s 314998 -960 315110 480 0 FreeSans 448 90 0 0 la_data_out[53]
port 347 nsew signal tristate
flabel metal2 s 318494 -960 318606 480 0 FreeSans 448 90 0 0 la_data_out[54]
port 348 nsew signal tristate
flabel metal2 s 322082 -960 322194 480 0 FreeSans 448 90 0 0 la_data_out[55]
port 349 nsew signal tristate
flabel metal2 s 325578 -960 325690 480 0 FreeSans 448 90 0 0 la_data_out[56]
port 350 nsew signal tristate
flabel metal2 s 329166 -960 329278 480 0 FreeSans 448 90 0 0 la_data_out[57]
port 351 nsew signal tristate
flabel metal2 s 332662 -960 332774 480 0 FreeSans 448 90 0 0 la_data_out[58]
port 352 nsew signal tristate
flabel metal2 s 336250 -960 336362 480 0 FreeSans 448 90 0 0 la_data_out[59]
port 353 nsew signal tristate
flabel metal2 s 144706 -960 144818 480 0 FreeSans 448 90 0 0 la_data_out[5]
port 354 nsew signal tristate
flabel metal2 s 339838 -960 339950 480 0 FreeSans 448 90 0 0 la_data_out[60]
port 355 nsew signal tristate
flabel metal2 s 343334 -960 343446 480 0 FreeSans 448 90 0 0 la_data_out[61]
port 356 nsew signal tristate
flabel metal2 s 346922 -960 347034 480 0 FreeSans 448 90 0 0 la_data_out[62]
port 357 nsew signal tristate
flabel metal2 s 350418 -960 350530 480 0 FreeSans 448 90 0 0 la_data_out[63]
port 358 nsew signal tristate
flabel metal2 s 354006 -960 354118 480 0 FreeSans 448 90 0 0 la_data_out[64]
port 359 nsew signal tristate
flabel metal2 s 357502 -960 357614 480 0 FreeSans 448 90 0 0 la_data_out[65]
port 360 nsew signal tristate
flabel metal2 s 361090 -960 361202 480 0 FreeSans 448 90 0 0 la_data_out[66]
port 361 nsew signal tristate
flabel metal2 s 364586 -960 364698 480 0 FreeSans 448 90 0 0 la_data_out[67]
port 362 nsew signal tristate
flabel metal2 s 368174 -960 368286 480 0 FreeSans 448 90 0 0 la_data_out[68]
port 363 nsew signal tristate
flabel metal2 s 371670 -960 371782 480 0 FreeSans 448 90 0 0 la_data_out[69]
port 364 nsew signal tristate
flabel metal2 s 148294 -960 148406 480 0 FreeSans 448 90 0 0 la_data_out[6]
port 365 nsew signal tristate
flabel metal2 s 375258 -960 375370 480 0 FreeSans 448 90 0 0 la_data_out[70]
port 366 nsew signal tristate
flabel metal2 s 378846 -960 378958 480 0 FreeSans 448 90 0 0 la_data_out[71]
port 367 nsew signal tristate
flabel metal2 s 382342 -960 382454 480 0 FreeSans 448 90 0 0 la_data_out[72]
port 368 nsew signal tristate
flabel metal2 s 385930 -960 386042 480 0 FreeSans 448 90 0 0 la_data_out[73]
port 369 nsew signal tristate
flabel metal2 s 389426 -960 389538 480 0 FreeSans 448 90 0 0 la_data_out[74]
port 370 nsew signal tristate
flabel metal2 s 393014 -960 393126 480 0 FreeSans 448 90 0 0 la_data_out[75]
port 371 nsew signal tristate
flabel metal2 s 396510 -960 396622 480 0 FreeSans 448 90 0 0 la_data_out[76]
port 372 nsew signal tristate
flabel metal2 s 400098 -960 400210 480 0 FreeSans 448 90 0 0 la_data_out[77]
port 373 nsew signal tristate
flabel metal2 s 403594 -960 403706 480 0 FreeSans 448 90 0 0 la_data_out[78]
port 374 nsew signal tristate
flabel metal2 s 407182 -960 407294 480 0 FreeSans 448 90 0 0 la_data_out[79]
port 375 nsew signal tristate
flabel metal2 s 151790 -960 151902 480 0 FreeSans 448 90 0 0 la_data_out[7]
port 376 nsew signal tristate
flabel metal2 s 410770 -960 410882 480 0 FreeSans 448 90 0 0 la_data_out[80]
port 377 nsew signal tristate
flabel metal2 s 414266 -960 414378 480 0 FreeSans 448 90 0 0 la_data_out[81]
port 378 nsew signal tristate
flabel metal2 s 417854 -960 417966 480 0 FreeSans 448 90 0 0 la_data_out[82]
port 379 nsew signal tristate
flabel metal2 s 421350 -960 421462 480 0 FreeSans 448 90 0 0 la_data_out[83]
port 380 nsew signal tristate
flabel metal2 s 424938 -960 425050 480 0 FreeSans 448 90 0 0 la_data_out[84]
port 381 nsew signal tristate
flabel metal2 s 428434 -960 428546 480 0 FreeSans 448 90 0 0 la_data_out[85]
port 382 nsew signal tristate
flabel metal2 s 432022 -960 432134 480 0 FreeSans 448 90 0 0 la_data_out[86]
port 383 nsew signal tristate
flabel metal2 s 435518 -960 435630 480 0 FreeSans 448 90 0 0 la_data_out[87]
port 384 nsew signal tristate
flabel metal2 s 439106 -960 439218 480 0 FreeSans 448 90 0 0 la_data_out[88]
port 385 nsew signal tristate
flabel metal2 s 442602 -960 442714 480 0 FreeSans 448 90 0 0 la_data_out[89]
port 386 nsew signal tristate
flabel metal2 s 155378 -960 155490 480 0 FreeSans 448 90 0 0 la_data_out[8]
port 387 nsew signal tristate
flabel metal2 s 446190 -960 446302 480 0 FreeSans 448 90 0 0 la_data_out[90]
port 388 nsew signal tristate
flabel metal2 s 449778 -960 449890 480 0 FreeSans 448 90 0 0 la_data_out[91]
port 389 nsew signal tristate
flabel metal2 s 453274 -960 453386 480 0 FreeSans 448 90 0 0 la_data_out[92]
port 390 nsew signal tristate
flabel metal2 s 456862 -960 456974 480 0 FreeSans 448 90 0 0 la_data_out[93]
port 391 nsew signal tristate
flabel metal2 s 460358 -960 460470 480 0 FreeSans 448 90 0 0 la_data_out[94]
port 392 nsew signal tristate
flabel metal2 s 463946 -960 464058 480 0 FreeSans 448 90 0 0 la_data_out[95]
port 393 nsew signal tristate
flabel metal2 s 467442 -960 467554 480 0 FreeSans 448 90 0 0 la_data_out[96]
port 394 nsew signal tristate
flabel metal2 s 471030 -960 471142 480 0 FreeSans 448 90 0 0 la_data_out[97]
port 395 nsew signal tristate
flabel metal2 s 474526 -960 474638 480 0 FreeSans 448 90 0 0 la_data_out[98]
port 396 nsew signal tristate
flabel metal2 s 478114 -960 478226 480 0 FreeSans 448 90 0 0 la_data_out[99]
port 397 nsew signal tristate
flabel metal2 s 158874 -960 158986 480 0 FreeSans 448 90 0 0 la_data_out[9]
port 398 nsew signal tristate
flabel metal2 s 128146 -960 128258 480 0 FreeSans 448 90 0 0 la_oenb[0]
port 399 nsew signal input
flabel metal2 s 482806 -960 482918 480 0 FreeSans 448 90 0 0 la_oenb[100]
port 400 nsew signal input
flabel metal2 s 486394 -960 486506 480 0 FreeSans 448 90 0 0 la_oenb[101]
port 401 nsew signal input
flabel metal2 s 489890 -960 490002 480 0 FreeSans 448 90 0 0 la_oenb[102]
port 402 nsew signal input
flabel metal2 s 493478 -960 493590 480 0 FreeSans 448 90 0 0 la_oenb[103]
port 403 nsew signal input
flabel metal2 s 497066 -960 497178 480 0 FreeSans 448 90 0 0 la_oenb[104]
port 404 nsew signal input
flabel metal2 s 500562 -960 500674 480 0 FreeSans 448 90 0 0 la_oenb[105]
port 405 nsew signal input
flabel metal2 s 504150 -960 504262 480 0 FreeSans 448 90 0 0 la_oenb[106]
port 406 nsew signal input
flabel metal2 s 507646 -960 507758 480 0 FreeSans 448 90 0 0 la_oenb[107]
port 407 nsew signal input
flabel metal2 s 511234 -960 511346 480 0 FreeSans 448 90 0 0 la_oenb[108]
port 408 nsew signal input
flabel metal2 s 514730 -960 514842 480 0 FreeSans 448 90 0 0 la_oenb[109]
port 409 nsew signal input
flabel metal2 s 163658 -960 163770 480 0 FreeSans 448 90 0 0 la_oenb[10]
port 410 nsew signal input
flabel metal2 s 518318 -960 518430 480 0 FreeSans 448 90 0 0 la_oenb[110]
port 411 nsew signal input
flabel metal2 s 521814 -960 521926 480 0 FreeSans 448 90 0 0 la_oenb[111]
port 412 nsew signal input
flabel metal2 s 525402 -960 525514 480 0 FreeSans 448 90 0 0 la_oenb[112]
port 413 nsew signal input
flabel metal2 s 528990 -960 529102 480 0 FreeSans 448 90 0 0 la_oenb[113]
port 414 nsew signal input
flabel metal2 s 532486 -960 532598 480 0 FreeSans 448 90 0 0 la_oenb[114]
port 415 nsew signal input
flabel metal2 s 536074 -960 536186 480 0 FreeSans 448 90 0 0 la_oenb[115]
port 416 nsew signal input
flabel metal2 s 539570 -960 539682 480 0 FreeSans 448 90 0 0 la_oenb[116]
port 417 nsew signal input
flabel metal2 s 543158 -960 543270 480 0 FreeSans 448 90 0 0 la_oenb[117]
port 418 nsew signal input
flabel metal2 s 546654 -960 546766 480 0 FreeSans 448 90 0 0 la_oenb[118]
port 419 nsew signal input
flabel metal2 s 550242 -960 550354 480 0 FreeSans 448 90 0 0 la_oenb[119]
port 420 nsew signal input
flabel metal2 s 167154 -960 167266 480 0 FreeSans 448 90 0 0 la_oenb[11]
port 421 nsew signal input
flabel metal2 s 553738 -960 553850 480 0 FreeSans 448 90 0 0 la_oenb[120]
port 422 nsew signal input
flabel metal2 s 557326 -960 557438 480 0 FreeSans 448 90 0 0 la_oenb[121]
port 423 nsew signal input
flabel metal2 s 560822 -960 560934 480 0 FreeSans 448 90 0 0 la_oenb[122]
port 424 nsew signal input
flabel metal2 s 564410 -960 564522 480 0 FreeSans 448 90 0 0 la_oenb[123]
port 425 nsew signal input
flabel metal2 s 567998 -960 568110 480 0 FreeSans 448 90 0 0 la_oenb[124]
port 426 nsew signal input
flabel metal2 s 571494 -960 571606 480 0 FreeSans 448 90 0 0 la_oenb[125]
port 427 nsew signal input
flabel metal2 s 575082 -960 575194 480 0 FreeSans 448 90 0 0 la_oenb[126]
port 428 nsew signal input
flabel metal2 s 578578 -960 578690 480 0 FreeSans 448 90 0 0 la_oenb[127]
port 429 nsew signal input
flabel metal2 s 170742 -960 170854 480 0 FreeSans 448 90 0 0 la_oenb[12]
port 430 nsew signal input
flabel metal2 s 174238 -960 174350 480 0 FreeSans 448 90 0 0 la_oenb[13]
port 431 nsew signal input
flabel metal2 s 177826 -960 177938 480 0 FreeSans 448 90 0 0 la_oenb[14]
port 432 nsew signal input
flabel metal2 s 181414 -960 181526 480 0 FreeSans 448 90 0 0 la_oenb[15]
port 433 nsew signal input
flabel metal2 s 184910 -960 185022 480 0 FreeSans 448 90 0 0 la_oenb[16]
port 434 nsew signal input
flabel metal2 s 188498 -960 188610 480 0 FreeSans 448 90 0 0 la_oenb[17]
port 435 nsew signal input
flabel metal2 s 191994 -960 192106 480 0 FreeSans 448 90 0 0 la_oenb[18]
port 436 nsew signal input
flabel metal2 s 195582 -960 195694 480 0 FreeSans 448 90 0 0 la_oenb[19]
port 437 nsew signal input
flabel metal2 s 131734 -960 131846 480 0 FreeSans 448 90 0 0 la_oenb[1]
port 438 nsew signal input
flabel metal2 s 199078 -960 199190 480 0 FreeSans 448 90 0 0 la_oenb[20]
port 439 nsew signal input
flabel metal2 s 202666 -960 202778 480 0 FreeSans 448 90 0 0 la_oenb[21]
port 440 nsew signal input
flabel metal2 s 206162 -960 206274 480 0 FreeSans 448 90 0 0 la_oenb[22]
port 441 nsew signal input
flabel metal2 s 209750 -960 209862 480 0 FreeSans 448 90 0 0 la_oenb[23]
port 442 nsew signal input
flabel metal2 s 213338 -960 213450 480 0 FreeSans 448 90 0 0 la_oenb[24]
port 443 nsew signal input
flabel metal2 s 216834 -960 216946 480 0 FreeSans 448 90 0 0 la_oenb[25]
port 444 nsew signal input
flabel metal2 s 220422 -960 220534 480 0 FreeSans 448 90 0 0 la_oenb[26]
port 445 nsew signal input
flabel metal2 s 223918 -960 224030 480 0 FreeSans 448 90 0 0 la_oenb[27]
port 446 nsew signal input
flabel metal2 s 227506 -960 227618 480 0 FreeSans 448 90 0 0 la_oenb[28]
port 447 nsew signal input
flabel metal2 s 231002 -960 231114 480 0 FreeSans 448 90 0 0 la_oenb[29]
port 448 nsew signal input
flabel metal2 s 135230 -960 135342 480 0 FreeSans 448 90 0 0 la_oenb[2]
port 449 nsew signal input
flabel metal2 s 234590 -960 234702 480 0 FreeSans 448 90 0 0 la_oenb[30]
port 450 nsew signal input
flabel metal2 s 238086 -960 238198 480 0 FreeSans 448 90 0 0 la_oenb[31]
port 451 nsew signal input
flabel metal2 s 241674 -960 241786 480 0 FreeSans 448 90 0 0 la_oenb[32]
port 452 nsew signal input
flabel metal2 s 245170 -960 245282 480 0 FreeSans 448 90 0 0 la_oenb[33]
port 453 nsew signal input
flabel metal2 s 248758 -960 248870 480 0 FreeSans 448 90 0 0 la_oenb[34]
port 454 nsew signal input
flabel metal2 s 252346 -960 252458 480 0 FreeSans 448 90 0 0 la_oenb[35]
port 455 nsew signal input
flabel metal2 s 255842 -960 255954 480 0 FreeSans 448 90 0 0 la_oenb[36]
port 456 nsew signal input
flabel metal2 s 259430 -960 259542 480 0 FreeSans 448 90 0 0 la_oenb[37]
port 457 nsew signal input
flabel metal2 s 262926 -960 263038 480 0 FreeSans 448 90 0 0 la_oenb[38]
port 458 nsew signal input
flabel metal2 s 266514 -960 266626 480 0 FreeSans 448 90 0 0 la_oenb[39]
port 459 nsew signal input
flabel metal2 s 138818 -960 138930 480 0 FreeSans 448 90 0 0 la_oenb[3]
port 460 nsew signal input
flabel metal2 s 270010 -960 270122 480 0 FreeSans 448 90 0 0 la_oenb[40]
port 461 nsew signal input
flabel metal2 s 273598 -960 273710 480 0 FreeSans 448 90 0 0 la_oenb[41]
port 462 nsew signal input
flabel metal2 s 277094 -960 277206 480 0 FreeSans 448 90 0 0 la_oenb[42]
port 463 nsew signal input
flabel metal2 s 280682 -960 280794 480 0 FreeSans 448 90 0 0 la_oenb[43]
port 464 nsew signal input
flabel metal2 s 284270 -960 284382 480 0 FreeSans 448 90 0 0 la_oenb[44]
port 465 nsew signal input
flabel metal2 s 287766 -960 287878 480 0 FreeSans 448 90 0 0 la_oenb[45]
port 466 nsew signal input
flabel metal2 s 291354 -960 291466 480 0 FreeSans 448 90 0 0 la_oenb[46]
port 467 nsew signal input
flabel metal2 s 294850 -960 294962 480 0 FreeSans 448 90 0 0 la_oenb[47]
port 468 nsew signal input
flabel metal2 s 298438 -960 298550 480 0 FreeSans 448 90 0 0 la_oenb[48]
port 469 nsew signal input
flabel metal2 s 301934 -960 302046 480 0 FreeSans 448 90 0 0 la_oenb[49]
port 470 nsew signal input
flabel metal2 s 142406 -960 142518 480 0 FreeSans 448 90 0 0 la_oenb[4]
port 471 nsew signal input
flabel metal2 s 305522 -960 305634 480 0 FreeSans 448 90 0 0 la_oenb[50]
port 472 nsew signal input
flabel metal2 s 309018 -960 309130 480 0 FreeSans 448 90 0 0 la_oenb[51]
port 473 nsew signal input
flabel metal2 s 312606 -960 312718 480 0 FreeSans 448 90 0 0 la_oenb[52]
port 474 nsew signal input
flabel metal2 s 316194 -960 316306 480 0 FreeSans 448 90 0 0 la_oenb[53]
port 475 nsew signal input
flabel metal2 s 319690 -960 319802 480 0 FreeSans 448 90 0 0 la_oenb[54]
port 476 nsew signal input
flabel metal2 s 323278 -960 323390 480 0 FreeSans 448 90 0 0 la_oenb[55]
port 477 nsew signal input
flabel metal2 s 326774 -960 326886 480 0 FreeSans 448 90 0 0 la_oenb[56]
port 478 nsew signal input
flabel metal2 s 330362 -960 330474 480 0 FreeSans 448 90 0 0 la_oenb[57]
port 479 nsew signal input
flabel metal2 s 333858 -960 333970 480 0 FreeSans 448 90 0 0 la_oenb[58]
port 480 nsew signal input
flabel metal2 s 337446 -960 337558 480 0 FreeSans 448 90 0 0 la_oenb[59]
port 481 nsew signal input
flabel metal2 s 145902 -960 146014 480 0 FreeSans 448 90 0 0 la_oenb[5]
port 482 nsew signal input
flabel metal2 s 340942 -960 341054 480 0 FreeSans 448 90 0 0 la_oenb[60]
port 483 nsew signal input
flabel metal2 s 344530 -960 344642 480 0 FreeSans 448 90 0 0 la_oenb[61]
port 484 nsew signal input
flabel metal2 s 348026 -960 348138 480 0 FreeSans 448 90 0 0 la_oenb[62]
port 485 nsew signal input
flabel metal2 s 351614 -960 351726 480 0 FreeSans 448 90 0 0 la_oenb[63]
port 486 nsew signal input
flabel metal2 s 355202 -960 355314 480 0 FreeSans 448 90 0 0 la_oenb[64]
port 487 nsew signal input
flabel metal2 s 358698 -960 358810 480 0 FreeSans 448 90 0 0 la_oenb[65]
port 488 nsew signal input
flabel metal2 s 362286 -960 362398 480 0 FreeSans 448 90 0 0 la_oenb[66]
port 489 nsew signal input
flabel metal2 s 365782 -960 365894 480 0 FreeSans 448 90 0 0 la_oenb[67]
port 490 nsew signal input
flabel metal2 s 369370 -960 369482 480 0 FreeSans 448 90 0 0 la_oenb[68]
port 491 nsew signal input
flabel metal2 s 372866 -960 372978 480 0 FreeSans 448 90 0 0 la_oenb[69]
port 492 nsew signal input
flabel metal2 s 149490 -960 149602 480 0 FreeSans 448 90 0 0 la_oenb[6]
port 493 nsew signal input
flabel metal2 s 376454 -960 376566 480 0 FreeSans 448 90 0 0 la_oenb[70]
port 494 nsew signal input
flabel metal2 s 379950 -960 380062 480 0 FreeSans 448 90 0 0 la_oenb[71]
port 495 nsew signal input
flabel metal2 s 383538 -960 383650 480 0 FreeSans 448 90 0 0 la_oenb[72]
port 496 nsew signal input
flabel metal2 s 387126 -960 387238 480 0 FreeSans 448 90 0 0 la_oenb[73]
port 497 nsew signal input
flabel metal2 s 390622 -960 390734 480 0 FreeSans 448 90 0 0 la_oenb[74]
port 498 nsew signal input
flabel metal2 s 394210 -960 394322 480 0 FreeSans 448 90 0 0 la_oenb[75]
port 499 nsew signal input
flabel metal2 s 397706 -960 397818 480 0 FreeSans 448 90 0 0 la_oenb[76]
port 500 nsew signal input
flabel metal2 s 401294 -960 401406 480 0 FreeSans 448 90 0 0 la_oenb[77]
port 501 nsew signal input
flabel metal2 s 404790 -960 404902 480 0 FreeSans 448 90 0 0 la_oenb[78]
port 502 nsew signal input
flabel metal2 s 408378 -960 408490 480 0 FreeSans 448 90 0 0 la_oenb[79]
port 503 nsew signal input
flabel metal2 s 152986 -960 153098 480 0 FreeSans 448 90 0 0 la_oenb[7]
port 504 nsew signal input
flabel metal2 s 411874 -960 411986 480 0 FreeSans 448 90 0 0 la_oenb[80]
port 505 nsew signal input
flabel metal2 s 415462 -960 415574 480 0 FreeSans 448 90 0 0 la_oenb[81]
port 506 nsew signal input
flabel metal2 s 418958 -960 419070 480 0 FreeSans 448 90 0 0 la_oenb[82]
port 507 nsew signal input
flabel metal2 s 422546 -960 422658 480 0 FreeSans 448 90 0 0 la_oenb[83]
port 508 nsew signal input
flabel metal2 s 426134 -960 426246 480 0 FreeSans 448 90 0 0 la_oenb[84]
port 509 nsew signal input
flabel metal2 s 429630 -960 429742 480 0 FreeSans 448 90 0 0 la_oenb[85]
port 510 nsew signal input
flabel metal2 s 433218 -960 433330 480 0 FreeSans 448 90 0 0 la_oenb[86]
port 511 nsew signal input
flabel metal2 s 436714 -960 436826 480 0 FreeSans 448 90 0 0 la_oenb[87]
port 512 nsew signal input
flabel metal2 s 440302 -960 440414 480 0 FreeSans 448 90 0 0 la_oenb[88]
port 513 nsew signal input
flabel metal2 s 443798 -960 443910 480 0 FreeSans 448 90 0 0 la_oenb[89]
port 514 nsew signal input
flabel metal2 s 156574 -960 156686 480 0 FreeSans 448 90 0 0 la_oenb[8]
port 515 nsew signal input
flabel metal2 s 447386 -960 447498 480 0 FreeSans 448 90 0 0 la_oenb[90]
port 516 nsew signal input
flabel metal2 s 450882 -960 450994 480 0 FreeSans 448 90 0 0 la_oenb[91]
port 517 nsew signal input
flabel metal2 s 454470 -960 454582 480 0 FreeSans 448 90 0 0 la_oenb[92]
port 518 nsew signal input
flabel metal2 s 458058 -960 458170 480 0 FreeSans 448 90 0 0 la_oenb[93]
port 519 nsew signal input
flabel metal2 s 461554 -960 461666 480 0 FreeSans 448 90 0 0 la_oenb[94]
port 520 nsew signal input
flabel metal2 s 465142 -960 465254 480 0 FreeSans 448 90 0 0 la_oenb[95]
port 521 nsew signal input
flabel metal2 s 468638 -960 468750 480 0 FreeSans 448 90 0 0 la_oenb[96]
port 522 nsew signal input
flabel metal2 s 472226 -960 472338 480 0 FreeSans 448 90 0 0 la_oenb[97]
port 523 nsew signal input
flabel metal2 s 475722 -960 475834 480 0 FreeSans 448 90 0 0 la_oenb[98]
port 524 nsew signal input
flabel metal2 s 479310 -960 479422 480 0 FreeSans 448 90 0 0 la_oenb[99]
port 525 nsew signal input
flabel metal2 s 160070 -960 160182 480 0 FreeSans 448 90 0 0 la_oenb[9]
port 526 nsew signal input
flabel metal2 s 579774 -960 579886 480 0 FreeSans 448 90 0 0 user_clock2
port 527 nsew signal input
flabel metal2 s 580970 -960 581082 480 0 FreeSans 448 90 0 0 user_irq[0]
port 528 nsew signal tristate
flabel metal2 s 582166 -960 582278 480 0 FreeSans 448 90 0 0 user_irq[1]
port 529 nsew signal tristate
flabel metal2 s 583362 -960 583474 480 0 FreeSans 448 90 0 0 user_irq[2]
port 530 nsew signal tristate
flabel metal4 s -2006 -934 -1386 704870 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -2006 -934 585930 -314 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -2006 704250 585930 704870 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 585310 -934 585930 704870 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 1794 -7654 2414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 37794 -7654 38414 24559 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 37794 133057 38414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 73794 -7654 74414 24068 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 73794 320601 74414 447495 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 73794 595705 74414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 109794 -7654 110414 24559 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 109794 133057 110414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 145794 -7654 146414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 181794 -7654 182414 50791 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 181794 131409 182414 270287 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 181794 423529 182414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 217794 -7654 218414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 253794 -7654 254414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 289794 -7654 290414 43007 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 289794 320417 290414 380831 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 289794 648313 290414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 325794 -7654 326414 40068 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 325794 320417 326414 380831 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 325794 648313 326414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 361794 -7654 362414 43007 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 361794 320417 362414 380831 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 361794 648313 362414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 397794 -7654 398414 43007 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 397794 320417 398414 380831 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 397794 648313 398414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 433794 -7654 434414 43007 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 433794 320417 434414 380831 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 433794 648313 434414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 469794 -7654 470414 43007 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 469794 320417 470414 380831 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 469794 648313 470414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 505794 -7654 506414 43007 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 505794 320417 506414 380831 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 505794 648313 506414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 541794 -7654 542414 43007 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 541794 320417 542414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 577794 -7654 578414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 2866 592650 3486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 38866 592650 39486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 74866 592650 75486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 110866 592650 111486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 146866 592650 147486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 182866 592650 183486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 218866 592650 219486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 254866 592650 255486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 290866 592650 291486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 326866 592650 327486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 362866 592650 363486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 398866 592650 399486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 434866 592650 435486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 470866 592650 471486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 506866 592650 507486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 542866 592650 543486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 578866 592650 579486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 614866 592650 615486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 650866 592650 651486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 686866 592650 687486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s -3926 -2854 -3306 706790 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -3926 -2854 587850 -2234 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -3926 706170 587850 706790 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 587230 -2854 587850 706790 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 9234 -7654 9854 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 45234 -7654 45854 24559 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 45234 133057 45854 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 81234 -7654 81854 24559 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 81234 320601 81854 447495 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 81234 595705 81854 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 117234 -7654 117854 24559 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 117234 133057 117854 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 153234 -7654 153854 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 189234 -7654 189854 50791 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 189234 131409 189854 270287 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 189234 423529 189854 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 225234 -7654 225854 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 261234 -7654 261854 43007 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 261234 320417 261854 380831 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 261234 648313 261854 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 297234 -7654 297854 43007 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 297234 320417 297854 380831 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 297234 648313 297854 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 333234 -7654 333854 43007 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 333234 320417 333854 380831 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 333234 648313 333854 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 369234 -7654 369854 43007 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 369234 320417 369854 380831 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 369234 648313 369854 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 405234 -7654 405854 43007 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 405234 320417 405854 380831 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 405234 648313 405854 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 441234 -7654 441854 43007 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 441234 320417 441854 380831 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 441234 648313 441854 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 477234 -7654 477854 43007 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 477234 320417 477854 380831 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 477234 648313 477854 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 513234 -7654 513854 43007 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 513234 320417 513854 380831 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 513234 648313 513854 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 549234 -7654 549854 43007 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 549234 320417 549854 380068 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 549234 649212 549854 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 10306 592650 10926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 46306 592650 46926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 82306 592650 82926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 118306 592650 118926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 154306 592650 154926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 190306 592650 190926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 226306 592650 226926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 262306 592650 262926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 298306 592650 298926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 334306 592650 334926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 370306 592650 370926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 406306 592650 406926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 442306 592650 442926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 478306 592650 478926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 514306 592650 514926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 550306 592650 550926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 586306 592650 586926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 622306 592650 622926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 658306 592650 658926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 694306 592650 694926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s -5846 -4774 -5226 708710 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -5846 -4774 589770 -4154 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -5846 708090 589770 708710 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 589150 -4774 589770 708710 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 16674 -7654 17294 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 52674 -7654 53294 24559 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 52674 133057 53294 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 88674 -7654 89294 24559 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 88674 133057 89294 167495 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 88674 320601 89294 447495 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 88674 595705 89294 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 124674 -7654 125294 24559 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 124674 133057 125294 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 160674 -7654 161294 50791 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 160674 131409 161294 270287 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 160674 423529 161294 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 196674 -7654 197294 270287 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 196674 423529 197294 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 232674 -7654 233294 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 268674 -7654 269294 43007 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 268674 320417 269294 380831 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 268674 648313 269294 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 304674 -7654 305294 43007 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 304674 320417 305294 380831 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 304674 648313 305294 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 340674 -7654 341294 40068 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 340674 320417 341294 380831 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 340674 648313 341294 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 376674 -7654 377294 43007 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 376674 320417 377294 380831 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 376674 648313 377294 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 412674 -7654 413294 43007 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 412674 320417 413294 380831 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 412674 648313 413294 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 448674 -7654 449294 40068 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 448674 320417 449294 380831 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 448674 648313 449294 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 484674 -7654 485294 43007 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 484674 320417 485294 380831 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 484674 648313 485294 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 520674 -7654 521294 43007 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 520674 320417 521294 380831 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 520674 648313 521294 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 556674 -7654 557294 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 17746 592650 18366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 53746 592650 54366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 89746 592650 90366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 125746 592650 126366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 161746 592650 162366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 197746 592650 198366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 233746 592650 234366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 269746 592650 270366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 305746 592650 306366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 341746 592650 342366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 377746 592650 378366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 413746 592650 414366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 449746 592650 450366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 485746 592650 486366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 521746 592650 522366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 557746 592650 558366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 593746 592650 594366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 629746 592650 630366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 665746 592650 666366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s -7766 -6694 -7146 710630 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -7766 -6694 591690 -6074 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -7766 710010 591690 710630 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 591070 -6694 591690 710630 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 24114 -7654 24734 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 60114 133057 60734 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 96114 133057 96734 167495 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 96114 320601 96734 447495 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 96114 595705 96734 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 132114 133057 132734 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 168114 -7654 168734 50791 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 168114 131409 168734 270287 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 168114 423529 168734 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 204114 -7654 204734 270287 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 204114 423529 204734 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 240114 -7654 240734 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 276114 -7654 276734 43007 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 276114 498713 276734 530431 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 276114 648313 276734 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 312114 -7654 312734 43007 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 312114 498713 312734 530431 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 312114 648313 312734 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 348114 -7654 348734 43007 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 348114 498713 348734 530431 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 348114 648313 348734 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 384114 -7654 384734 43007 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 384114 498713 384734 530431 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 384114 648313 384734 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 420114 -7654 420734 43007 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 420114 498713 420734 530431 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 420114 648313 420734 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 456114 -7654 456734 43007 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 456114 498713 456734 530431 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 456114 648313 456734 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 492114 -7654 492734 43007 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 492114 498713 492734 530431 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 492114 648313 492734 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 528114 -7654 528734 43007 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 528114 498713 528734 530431 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 528114 648313 528734 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 564114 -7654 564734 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 25186 592650 25806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 61186 592650 61806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 97186 592650 97806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 133186 592650 133806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 169186 592650 169806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 205186 592650 205806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 241186 592650 241806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 277186 592650 277806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 313186 592650 313806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 349186 592650 349806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 385186 592650 385806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 421186 592650 421806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 457186 592650 457806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 493186 592650 493806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 529186 592650 529806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 565186 592650 565806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 601186 592650 601806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 637186 592650 637806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 673186 592650 673806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s -6806 -5734 -6186 709670 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -6806 -5734 590730 -5114 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -6806 709050 590730 709670 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 590110 -5734 590730 709670 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 20394 -7654 21014 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 56394 -7654 57014 24559 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 56394 133057 57014 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 92394 -7654 93014 24559 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 92394 133057 93014 167495 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 92394 320601 93014 447495 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 92394 595705 93014 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 128394 -7654 129014 24559 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 128394 133057 129014 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 164394 -7654 165014 50791 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 164394 131409 165014 270287 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 164394 423529 165014 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 200394 -7654 201014 270287 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 200394 423529 201014 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 236394 -7654 237014 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 272394 -7654 273014 43007 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 272394 648313 273014 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 308394 -7654 309014 43007 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 308394 648313 309014 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 344394 -7654 345014 43007 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 344394 648313 345014 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 380394 -7654 381014 43007 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 380394 649212 381014 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 416394 -7654 417014 43007 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 416394 648313 417014 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 452394 -7654 453014 43007 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 452394 648313 453014 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 488394 -7654 489014 43007 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 488394 649212 489014 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 524394 -7654 525014 43007 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 524394 648313 525014 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 560394 -7654 561014 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 21466 592650 22086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 57466 592650 58086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 93466 592650 94086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 129466 592650 130086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 165466 592650 166086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 201466 592650 202086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 237466 592650 238086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 273466 592650 274086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 309466 592650 310086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 345466 592650 346086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 381466 592650 382086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 417466 592650 418086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 453466 592650 454086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 489466 592650 490086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 525466 592650 526086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 561466 592650 562086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 597466 592650 598086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 633466 592650 634086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 669466 592650 670086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s -8726 -7654 -8106 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 -7654 592650 -7034 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 710970 592650 711590 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 592030 -7654 592650 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 27834 133820 28454 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 63834 320601 64454 447495 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 63834 595705 64454 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 99834 320601 100454 447495 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 99834 595705 100454 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 135834 -7654 136454 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 171834 -7654 172454 50791 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 171834 131409 172454 270287 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 171834 423529 172454 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 207834 -7654 208454 52068 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 207834 131900 208454 270068 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 207834 429868 208454 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 243834 -7654 244454 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 279834 -7654 280454 40068 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 279834 648313 280454 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 315834 -7654 316454 43007 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 315834 648313 316454 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 351834 -7654 352454 43007 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 351834 648313 352454 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 387834 -7654 388454 43007 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 387834 648313 388454 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 423834 -7654 424454 43007 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 423834 648313 424454 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 459834 -7654 460454 43007 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 459834 648313 460454 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 495834 -7654 496454 43007 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 495834 648313 496454 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 531834 -7654 532454 43007 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 531834 648313 532454 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 567834 -7654 568454 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 28906 592650 29526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 64906 592650 65526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 100906 592650 101526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 136906 592650 137526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 172906 592650 173526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 208906 592650 209526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 244906 592650 245526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 280906 592650 281526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 316906 592650 317526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 352906 592650 353526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 388906 592650 389526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 424906 592650 425526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 460906 592650 461526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 496906 592650 497526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 532906 592650 533526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 568906 592650 569526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 604906 592650 605526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 640906 592650 641526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 676906 592650 677526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s -2966 -1894 -2346 705830 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -2966 -1894 586890 -1274 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -2966 705210 586890 705830 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 586270 -1894 586890 705830 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 5514 -7654 6134 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 41514 -7654 42134 24559 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 41514 133057 42134 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 77514 -7654 78134 24559 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 77514 320601 78134 447495 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 77514 595705 78134 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 113514 -7654 114134 24559 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 113514 133057 114134 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 149514 -7654 150134 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 185514 -7654 186134 50791 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 185514 131409 186134 270287 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 185514 423529 186134 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 221514 -7654 222134 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 257514 -7654 258134 380068 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 257514 649212 258134 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 293514 -7654 294134 43007 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 293514 320417 294134 380831 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 293514 648313 294134 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 329514 -7654 330134 43007 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 329514 320417 330134 380831 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 329514 648313 330134 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 365514 -7654 366134 43007 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 365514 320417 366134 380068 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 365514 649212 366134 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 401514 -7654 402134 43007 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 401514 320417 402134 380831 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 401514 648313 402134 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 437514 -7654 438134 43007 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 437514 320417 438134 380831 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 437514 648313 438134 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 473514 -7654 474134 43007 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 473514 320417 474134 380831 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 473514 648313 474134 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 509514 -7654 510134 40068 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 509514 320417 510134 380831 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 509514 648313 510134 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 545514 -7654 546134 43007 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 545514 320417 546134 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 581514 -7654 582134 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 6586 592650 7206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 42586 592650 43206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 78586 592650 79206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 114586 592650 115206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 150586 592650 151206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 186586 592650 187206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 222586 592650 223206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 258586 592650 259206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 294586 592650 295206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 330586 592650 331206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 366586 592650 367206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 402586 592650 403206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 438586 592650 439206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 474586 592650 475206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 510586 592650 511206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 546586 592650 547206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 582586 592650 583206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 618586 592650 619206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 654586 592650 655206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 690586 592650 691206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s -4886 -3814 -4266 707750 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -4886 -3814 588810 -3194 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -4886 707130 588810 707750 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 588190 -3814 588810 707750 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 12954 -7654 13574 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 48954 -7654 49574 24559 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 48954 323676 49574 440068 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 48954 599868 49574 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 84954 -7654 85574 24559 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 84954 320601 85574 447495 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 84954 595705 85574 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 120954 -7654 121574 24559 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 120954 133057 121574 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 156954 -7654 157574 270287 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 156954 423529 157574 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 192954 -7654 193574 52068 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 192954 131900 193574 270068 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 192954 429868 193574 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 228954 -7654 229574 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 264954 -7654 265574 43007 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 264954 320417 265574 380831 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 264954 648313 265574 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 300954 -7654 301574 43007 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 300954 320417 301574 380831 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 300954 648313 301574 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 336954 -7654 337574 43007 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 336954 320417 337574 380831 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 336954 648313 337574 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 372954 -7654 373574 43007 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 372954 320417 373574 380831 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 372954 648313 373574 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 408954 -7654 409574 43007 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 408954 320417 409574 380831 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 408954 648313 409574 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 444954 -7654 445574 43007 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 444954 320417 445574 380831 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 444954 648313 445574 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 480954 -7654 481574 43007 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 480954 320417 481574 380831 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 480954 648313 481574 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 516954 -7654 517574 43007 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 516954 320417 517574 380831 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 516954 648313 517574 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 552954 -7654 553574 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 14026 592650 14646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 50026 592650 50646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 86026 592650 86646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 122026 592650 122646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 158026 592650 158646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 194026 592650 194646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 230026 592650 230646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 266026 592650 266646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 302026 592650 302646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 338026 592650 338646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 374026 592650 374646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 410026 592650 410646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 446026 592650 446646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 482026 592650 482646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 518026 592650 518646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 554026 592650 554646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 590026 592650 590646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 626026 592650 626646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 662026 592650 662646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 698026 592650 698646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal2 s 542 -960 654 480 0 FreeSans 448 90 0 0 wb_clk_i
port 539 nsew signal input
flabel metal2 s 1646 -960 1758 480 0 FreeSans 448 90 0 0 wb_rst_i
port 540 nsew signal input
flabel metal2 s 2842 -960 2954 480 0 FreeSans 448 90 0 0 wbs_ack_o
port 541 nsew signal tristate
flabel metal2 s 7626 -960 7738 480 0 FreeSans 448 90 0 0 wbs_adr_i[0]
port 542 nsew signal input
flabel metal2 s 47830 -960 47942 480 0 FreeSans 448 90 0 0 wbs_adr_i[10]
port 543 nsew signal input
flabel metal2 s 51326 -960 51438 480 0 FreeSans 448 90 0 0 wbs_adr_i[11]
port 544 nsew signal input
flabel metal2 s 54914 -960 55026 480 0 FreeSans 448 90 0 0 wbs_adr_i[12]
port 545 nsew signal input
flabel metal2 s 58410 -960 58522 480 0 FreeSans 448 90 0 0 wbs_adr_i[13]
port 546 nsew signal input
flabel metal2 s 61998 -960 62110 480 0 FreeSans 448 90 0 0 wbs_adr_i[14]
port 547 nsew signal input
flabel metal2 s 65494 -960 65606 480 0 FreeSans 448 90 0 0 wbs_adr_i[15]
port 548 nsew signal input
flabel metal2 s 69082 -960 69194 480 0 FreeSans 448 90 0 0 wbs_adr_i[16]
port 549 nsew signal input
flabel metal2 s 72578 -960 72690 480 0 FreeSans 448 90 0 0 wbs_adr_i[17]
port 550 nsew signal input
flabel metal2 s 76166 -960 76278 480 0 FreeSans 448 90 0 0 wbs_adr_i[18]
port 551 nsew signal input
flabel metal2 s 79662 -960 79774 480 0 FreeSans 448 90 0 0 wbs_adr_i[19]
port 552 nsew signal input
flabel metal2 s 12318 -960 12430 480 0 FreeSans 448 90 0 0 wbs_adr_i[1]
port 553 nsew signal input
flabel metal2 s 83250 -960 83362 480 0 FreeSans 448 90 0 0 wbs_adr_i[20]
port 554 nsew signal input
flabel metal2 s 86838 -960 86950 480 0 FreeSans 448 90 0 0 wbs_adr_i[21]
port 555 nsew signal input
flabel metal2 s 90334 -960 90446 480 0 FreeSans 448 90 0 0 wbs_adr_i[22]
port 556 nsew signal input
flabel metal2 s 93922 -960 94034 480 0 FreeSans 448 90 0 0 wbs_adr_i[23]
port 557 nsew signal input
flabel metal2 s 97418 -960 97530 480 0 FreeSans 448 90 0 0 wbs_adr_i[24]
port 558 nsew signal input
flabel metal2 s 101006 -960 101118 480 0 FreeSans 448 90 0 0 wbs_adr_i[25]
port 559 nsew signal input
flabel metal2 s 104502 -960 104614 480 0 FreeSans 448 90 0 0 wbs_adr_i[26]
port 560 nsew signal input
flabel metal2 s 108090 -960 108202 480 0 FreeSans 448 90 0 0 wbs_adr_i[27]
port 561 nsew signal input
flabel metal2 s 111586 -960 111698 480 0 FreeSans 448 90 0 0 wbs_adr_i[28]
port 562 nsew signal input
flabel metal2 s 115174 -960 115286 480 0 FreeSans 448 90 0 0 wbs_adr_i[29]
port 563 nsew signal input
flabel metal2 s 17010 -960 17122 480 0 FreeSans 448 90 0 0 wbs_adr_i[2]
port 564 nsew signal input
flabel metal2 s 118762 -960 118874 480 0 FreeSans 448 90 0 0 wbs_adr_i[30]
port 565 nsew signal input
flabel metal2 s 122258 -960 122370 480 0 FreeSans 448 90 0 0 wbs_adr_i[31]
port 566 nsew signal input
flabel metal2 s 21794 -960 21906 480 0 FreeSans 448 90 0 0 wbs_adr_i[3]
port 567 nsew signal input
flabel metal2 s 26486 -960 26598 480 0 FreeSans 448 90 0 0 wbs_adr_i[4]
port 568 nsew signal input
flabel metal2 s 30074 -960 30186 480 0 FreeSans 448 90 0 0 wbs_adr_i[5]
port 569 nsew signal input
flabel metal2 s 33570 -960 33682 480 0 FreeSans 448 90 0 0 wbs_adr_i[6]
port 570 nsew signal input
flabel metal2 s 37158 -960 37270 480 0 FreeSans 448 90 0 0 wbs_adr_i[7]
port 571 nsew signal input
flabel metal2 s 40654 -960 40766 480 0 FreeSans 448 90 0 0 wbs_adr_i[8]
port 572 nsew signal input
flabel metal2 s 44242 -960 44354 480 0 FreeSans 448 90 0 0 wbs_adr_i[9]
port 573 nsew signal input
flabel metal2 s 4038 -960 4150 480 0 FreeSans 448 90 0 0 wbs_cyc_i
port 574 nsew signal input
flabel metal2 s 8730 -960 8842 480 0 FreeSans 448 90 0 0 wbs_dat_i[0]
port 575 nsew signal input
flabel metal2 s 48934 -960 49046 480 0 FreeSans 448 90 0 0 wbs_dat_i[10]
port 576 nsew signal input
flabel metal2 s 52522 -960 52634 480 0 FreeSans 448 90 0 0 wbs_dat_i[11]
port 577 nsew signal input
flabel metal2 s 56018 -960 56130 480 0 FreeSans 448 90 0 0 wbs_dat_i[12]
port 578 nsew signal input
flabel metal2 s 59606 -960 59718 480 0 FreeSans 448 90 0 0 wbs_dat_i[13]
port 579 nsew signal input
flabel metal2 s 63194 -960 63306 480 0 FreeSans 448 90 0 0 wbs_dat_i[14]
port 580 nsew signal input
flabel metal2 s 66690 -960 66802 480 0 FreeSans 448 90 0 0 wbs_dat_i[15]
port 581 nsew signal input
flabel metal2 s 70278 -960 70390 480 0 FreeSans 448 90 0 0 wbs_dat_i[16]
port 582 nsew signal input
flabel metal2 s 73774 -960 73886 480 0 FreeSans 448 90 0 0 wbs_dat_i[17]
port 583 nsew signal input
flabel metal2 s 77362 -960 77474 480 0 FreeSans 448 90 0 0 wbs_dat_i[18]
port 584 nsew signal input
flabel metal2 s 80858 -960 80970 480 0 FreeSans 448 90 0 0 wbs_dat_i[19]
port 585 nsew signal input
flabel metal2 s 13514 -960 13626 480 0 FreeSans 448 90 0 0 wbs_dat_i[1]
port 586 nsew signal input
flabel metal2 s 84446 -960 84558 480 0 FreeSans 448 90 0 0 wbs_dat_i[20]
port 587 nsew signal input
flabel metal2 s 87942 -960 88054 480 0 FreeSans 448 90 0 0 wbs_dat_i[21]
port 588 nsew signal input
flabel metal2 s 91530 -960 91642 480 0 FreeSans 448 90 0 0 wbs_dat_i[22]
port 589 nsew signal input
flabel metal2 s 95118 -960 95230 480 0 FreeSans 448 90 0 0 wbs_dat_i[23]
port 590 nsew signal input
flabel metal2 s 98614 -960 98726 480 0 FreeSans 448 90 0 0 wbs_dat_i[24]
port 591 nsew signal input
flabel metal2 s 102202 -960 102314 480 0 FreeSans 448 90 0 0 wbs_dat_i[25]
port 592 nsew signal input
flabel metal2 s 105698 -960 105810 480 0 FreeSans 448 90 0 0 wbs_dat_i[26]
port 593 nsew signal input
flabel metal2 s 109286 -960 109398 480 0 FreeSans 448 90 0 0 wbs_dat_i[27]
port 594 nsew signal input
flabel metal2 s 112782 -960 112894 480 0 FreeSans 448 90 0 0 wbs_dat_i[28]
port 595 nsew signal input
flabel metal2 s 116370 -960 116482 480 0 FreeSans 448 90 0 0 wbs_dat_i[29]
port 596 nsew signal input
flabel metal2 s 18206 -960 18318 480 0 FreeSans 448 90 0 0 wbs_dat_i[2]
port 597 nsew signal input
flabel metal2 s 119866 -960 119978 480 0 FreeSans 448 90 0 0 wbs_dat_i[30]
port 598 nsew signal input
flabel metal2 s 123454 -960 123566 480 0 FreeSans 448 90 0 0 wbs_dat_i[31]
port 599 nsew signal input
flabel metal2 s 22990 -960 23102 480 0 FreeSans 448 90 0 0 wbs_dat_i[3]
port 600 nsew signal input
flabel metal2 s 27682 -960 27794 480 0 FreeSans 448 90 0 0 wbs_dat_i[4]
port 601 nsew signal input
flabel metal2 s 31270 -960 31382 480 0 FreeSans 448 90 0 0 wbs_dat_i[5]
port 602 nsew signal input
flabel metal2 s 34766 -960 34878 480 0 FreeSans 448 90 0 0 wbs_dat_i[6]
port 603 nsew signal input
flabel metal2 s 38354 -960 38466 480 0 FreeSans 448 90 0 0 wbs_dat_i[7]
port 604 nsew signal input
flabel metal2 s 41850 -960 41962 480 0 FreeSans 448 90 0 0 wbs_dat_i[8]
port 605 nsew signal input
flabel metal2 s 45438 -960 45550 480 0 FreeSans 448 90 0 0 wbs_dat_i[9]
port 606 nsew signal input
flabel metal2 s 9926 -960 10038 480 0 FreeSans 448 90 0 0 wbs_dat_o[0]
port 607 nsew signal tristate
flabel metal2 s 50130 -960 50242 480 0 FreeSans 448 90 0 0 wbs_dat_o[10]
port 608 nsew signal tristate
flabel metal2 s 53718 -960 53830 480 0 FreeSans 448 90 0 0 wbs_dat_o[11]
port 609 nsew signal tristate
flabel metal2 s 57214 -960 57326 480 0 FreeSans 448 90 0 0 wbs_dat_o[12]
port 610 nsew signal tristate
flabel metal2 s 60802 -960 60914 480 0 FreeSans 448 90 0 0 wbs_dat_o[13]
port 611 nsew signal tristate
flabel metal2 s 64298 -960 64410 480 0 FreeSans 448 90 0 0 wbs_dat_o[14]
port 612 nsew signal tristate
flabel metal2 s 67886 -960 67998 480 0 FreeSans 448 90 0 0 wbs_dat_o[15]
port 613 nsew signal tristate
flabel metal2 s 71474 -960 71586 480 0 FreeSans 448 90 0 0 wbs_dat_o[16]
port 614 nsew signal tristate
flabel metal2 s 74970 -960 75082 480 0 FreeSans 448 90 0 0 wbs_dat_o[17]
port 615 nsew signal tristate
flabel metal2 s 78558 -960 78670 480 0 FreeSans 448 90 0 0 wbs_dat_o[18]
port 616 nsew signal tristate
flabel metal2 s 82054 -960 82166 480 0 FreeSans 448 90 0 0 wbs_dat_o[19]
port 617 nsew signal tristate
flabel metal2 s 14710 -960 14822 480 0 FreeSans 448 90 0 0 wbs_dat_o[1]
port 618 nsew signal tristate
flabel metal2 s 85642 -960 85754 480 0 FreeSans 448 90 0 0 wbs_dat_o[20]
port 619 nsew signal tristate
flabel metal2 s 89138 -960 89250 480 0 FreeSans 448 90 0 0 wbs_dat_o[21]
port 620 nsew signal tristate
flabel metal2 s 92726 -960 92838 480 0 FreeSans 448 90 0 0 wbs_dat_o[22]
port 621 nsew signal tristate
flabel metal2 s 96222 -960 96334 480 0 FreeSans 448 90 0 0 wbs_dat_o[23]
port 622 nsew signal tristate
flabel metal2 s 99810 -960 99922 480 0 FreeSans 448 90 0 0 wbs_dat_o[24]
port 623 nsew signal tristate
flabel metal2 s 103306 -960 103418 480 0 FreeSans 448 90 0 0 wbs_dat_o[25]
port 624 nsew signal tristate
flabel metal2 s 106894 -960 107006 480 0 FreeSans 448 90 0 0 wbs_dat_o[26]
port 625 nsew signal tristate
flabel metal2 s 110482 -960 110594 480 0 FreeSans 448 90 0 0 wbs_dat_o[27]
port 626 nsew signal tristate
flabel metal2 s 113978 -960 114090 480 0 FreeSans 448 90 0 0 wbs_dat_o[28]
port 627 nsew signal tristate
flabel metal2 s 117566 -960 117678 480 0 FreeSans 448 90 0 0 wbs_dat_o[29]
port 628 nsew signal tristate
flabel metal2 s 19402 -960 19514 480 0 FreeSans 448 90 0 0 wbs_dat_o[2]
port 629 nsew signal tristate
flabel metal2 s 121062 -960 121174 480 0 FreeSans 448 90 0 0 wbs_dat_o[30]
port 630 nsew signal tristate
flabel metal2 s 124650 -960 124762 480 0 FreeSans 448 90 0 0 wbs_dat_o[31]
port 631 nsew signal tristate
flabel metal2 s 24186 -960 24298 480 0 FreeSans 448 90 0 0 wbs_dat_o[3]
port 632 nsew signal tristate
flabel metal2 s 28878 -960 28990 480 0 FreeSans 448 90 0 0 wbs_dat_o[4]
port 633 nsew signal tristate
flabel metal2 s 32374 -960 32486 480 0 FreeSans 448 90 0 0 wbs_dat_o[5]
port 634 nsew signal tristate
flabel metal2 s 35962 -960 36074 480 0 FreeSans 448 90 0 0 wbs_dat_o[6]
port 635 nsew signal tristate
flabel metal2 s 39550 -960 39662 480 0 FreeSans 448 90 0 0 wbs_dat_o[7]
port 636 nsew signal tristate
flabel metal2 s 43046 -960 43158 480 0 FreeSans 448 90 0 0 wbs_dat_o[8]
port 637 nsew signal tristate
flabel metal2 s 46634 -960 46746 480 0 FreeSans 448 90 0 0 wbs_dat_o[9]
port 638 nsew signal tristate
flabel metal2 s 11122 -960 11234 480 0 FreeSans 448 90 0 0 wbs_sel_i[0]
port 639 nsew signal input
flabel metal2 s 15906 -960 16018 480 0 FreeSans 448 90 0 0 wbs_sel_i[1]
port 640 nsew signal input
flabel metal2 s 20598 -960 20710 480 0 FreeSans 448 90 0 0 wbs_sel_i[2]
port 641 nsew signal input
flabel metal2 s 25290 -960 25402 480 0 FreeSans 448 90 0 0 wbs_sel_i[3]
port 642 nsew signal input
flabel metal2 s 5234 -960 5346 480 0 FreeSans 448 90 0 0 wbs_stb_i
port 643 nsew signal input
flabel metal2 s 6430 -960 6542 480 0 FreeSans 448 90 0 0 wbs_we_i
port 644 nsew signal input
rlabel via4 218264 111336 218264 111336 0 vccd1
rlabel via4 81704 442776 81704 442776 0 vccd2
rlabel via4 197144 126216 197144 126216 0 vdda1
rlabel via4 204584 97656 204584 97656 0 vdda2
rlabel via4 200864 129936 200864 129936 0 vssa1
rlabel via4 172304 425376 172304 425376 0 vssa2
rlabel via4 208448 115056 208448 115056 0 vssd1
rlabel via4 553424 626496 553424 626496 0 vssd2
rlabel metal2 580198 6715 580198 6715 0 io_in[0]
rlabel metal2 580198 457453 580198 457453 0 io_in[10]
rlabel metal2 234094 280585 234094 280585 0 io_in[11]
rlabel metal3 582092 564332 582092 564332 0 io_in[12]
rlabel metal2 580198 617185 580198 617185 0 io_in[13]
rlabel metal4 251804 361692 251804 361692 0 io_in[14]
rlabel metal2 559682 701957 559682 701957 0 io_in[15]
rlabel metal1 369196 700434 369196 700434 0 io_in[16]
rlabel metal2 253322 375887 253322 375887 0 io_in[17]
rlabel metal2 365010 702212 365010 702212 0 io_in[18]
rlabel metal2 253230 375700 253230 375700 0 io_in[19]
rlabel metal3 582184 46308 582184 46308 0 io_in[1]
rlabel metal2 234830 703596 234830 703596 0 io_in[20]
rlabel metal1 164128 429862 164128 429862 0 io_in[21]
rlabel metal1 124154 700570 124154 700570 0 io_in[22]
rlabel metal2 40526 701940 40526 701940 0 io_in[23]
rlabel metal3 1878 684284 1878 684284 0 io_in[24]
rlabel metal3 1878 632060 1878 632060 0 io_in[25]
rlabel metal3 1832 579972 1832 579972 0 io_in[26]
rlabel metal3 1648 527884 1648 527884 0 io_in[27]
rlabel metal3 1970 475660 1970 475660 0 io_in[28]
rlabel metal3 1832 423572 1832 423572 0 io_in[29]
rlabel metal3 582230 86156 582230 86156 0 io_in[2]
rlabel metal3 1832 371348 1832 371348 0 io_in[30]
rlabel metal3 1878 319260 1878 319260 0 io_in[31]
rlabel metal3 1694 267172 1694 267172 0 io_in[32]
rlabel metal3 1832 214948 1832 214948 0 io_in[33]
rlabel metal3 1832 162860 1832 162860 0 io_in[34]
rlabel metal3 1878 110636 1878 110636 0 io_in[35]
rlabel metal3 1924 71604 1924 71604 0 io_in[36]
rlabel metal3 2062 32436 2062 32436 0 io_in[37]
rlabel metal3 582138 126004 582138 126004 0 io_in[3]
rlabel metal3 582092 165852 582092 165852 0 io_in[4]
rlabel metal3 582000 205700 582000 205700 0 io_in[5]
rlabel metal3 581954 245548 581954 245548 0 io_in[6]
rlabel metal3 581908 298724 581908 298724 0 io_in[7]
rlabel via2 580198 351917 580198 351917 0 io_in[8]
rlabel metal3 582230 404940 582230 404940 0 io_in[9]
rlabel metal3 581954 33116 581954 33116 0 io_oeb[0]
rlabel metal3 582046 484636 582046 484636 0 io_oeb[10]
rlabel metal2 580198 533545 580198 533545 0 io_oeb[11]
rlabel metal3 582000 590988 582000 590988 0 io_oeb[12]
rlabel metal3 582046 644028 582046 644028 0 io_oeb[13]
rlabel metal2 580198 697085 580198 697085 0 io_oeb[14]
rlabel metal2 527206 701974 527206 701974 0 io_oeb[15]
rlabel metal2 249090 375683 249090 375683 0 io_oeb[16]
rlabel metal1 319148 700774 319148 700774 0 io_oeb[17]
rlabel metal2 332534 702280 332534 702280 0 io_oeb[18]
rlabel metal2 238050 375666 238050 375666 0 io_oeb[19]
rlabel metal3 581862 72964 581862 72964 0 io_oeb[1]
rlabel metal1 210496 700298 210496 700298 0 io_oeb[20]
rlabel metal2 137172 703596 137172 703596 0 io_oeb[21]
rlabel metal1 110676 700434 110676 700434 0 io_oeb[22]
rlabel metal2 153962 91035 153962 91035 0 io_oeb[23]
rlabel metal3 1878 658172 1878 658172 0 io_oeb[24]
rlabel metal3 1786 606084 1786 606084 0 io_oeb[25]
rlabel metal3 1878 553860 1878 553860 0 io_oeb[26]
rlabel metal3 1924 501772 1924 501772 0 io_oeb[27]
rlabel metal3 2062 449548 2062 449548 0 io_oeb[28]
rlabel metal3 1832 397460 1832 397460 0 io_oeb[29]
rlabel metal2 580198 112319 580198 112319 0 io_oeb[2]
rlabel metal3 1694 345372 1694 345372 0 io_oeb[30]
rlabel metal3 1878 293148 1878 293148 0 io_oeb[31]
rlabel metal3 1924 241060 1924 241060 0 io_oeb[32]
rlabel metal3 1970 188836 1970 188836 0 io_oeb[33]
rlabel metal3 1878 136748 1878 136748 0 io_oeb[34]
rlabel metal3 1878 84660 1878 84660 0 io_oeb[35]
rlabel metal3 2016 45492 2016 45492 0 io_oeb[36]
rlabel metal3 1878 6460 1878 6460 0 io_oeb[37]
rlabel metal2 580014 152235 580014 152235 0 io_oeb[3]
rlabel metal3 582046 192508 582046 192508 0 io_oeb[4]
rlabel metal2 579646 232101 579646 232101 0 io_oeb[5]
rlabel metal2 580198 272051 580198 272051 0 io_oeb[6]
rlabel metal2 580198 324785 580198 324785 0 io_oeb[7]
rlabel metal2 579830 378301 579830 378301 0 io_oeb[8]
rlabel metal3 582138 431596 582138 431596 0 io_oeb[9]
rlabel metal3 581908 19788 581908 19788 0 io_out[0]
rlabel metal3 582092 471444 582092 471444 0 io_out[10]
rlabel via2 580198 524467 580198 524467 0 io_out[11]
rlabel metal3 581954 577660 581954 577660 0 io_out[12]
rlabel metal2 229770 184195 229770 184195 0 io_out[13]
rlabel metal2 580198 683519 580198 683519 0 io_out[14]
rlabel metal2 232530 375887 232530 375887 0 io_out[15]
rlabel metal2 233910 375445 233910 375445 0 io_out[16]
rlabel metal1 316204 700638 316204 700638 0 io_out[17]
rlabel metal2 348818 702246 348818 702246 0 io_out[18]
rlabel metal2 251850 374204 251850 374204 0 io_out[19]
rlabel metal2 580106 59517 580106 59517 0 io_out[1]
rlabel metal2 218454 703596 218454 703596 0 io_out[20]
rlabel metal2 153686 702420 153686 702420 0 io_out[21]
rlabel metal1 120152 700502 120152 700502 0 io_out[22]
rlabel metal2 24334 701974 24334 701974 0 io_out[23]
rlabel metal3 1924 671228 1924 671228 0 io_out[24]
rlabel metal3 1740 619140 1740 619140 0 io_out[25]
rlabel metal3 1878 566916 1878 566916 0 io_out[26]
rlabel metal3 1924 514828 1924 514828 0 io_out[27]
rlabel metal3 2016 462604 2016 462604 0 io_out[28]
rlabel metal3 1832 410516 1832 410516 0 io_out[29]
rlabel metal3 582184 99484 582184 99484 0 io_out[2]
rlabel metal3 1648 358428 1648 358428 0 io_out[30]
rlabel metal3 1786 306204 1786 306204 0 io_out[31]
rlabel metal3 1924 254116 1924 254116 0 io_out[32]
rlabel metal3 1786 201892 1786 201892 0 io_out[33]
rlabel metal3 1878 149804 1878 149804 0 io_out[34]
rlabel metal3 1878 97580 1878 97580 0 io_out[35]
rlabel metal3 1970 58548 1970 58548 0 io_out[36]
rlabel metal3 1878 19380 1878 19380 0 io_out[37]
rlabel metal2 580198 138669 580198 138669 0 io_out[3]
rlabel metal2 580198 178619 580198 178619 0 io_out[4]
rlabel metal2 580198 218535 580198 218535 0 io_out[5]
rlabel metal2 580198 258485 580198 258485 0 io_out[6]
rlabel metal3 582000 312052 582000 312052 0 io_out[7]
rlabel metal2 580014 364735 580014 364735 0 io_out[8]
rlabel metal3 582184 418268 582184 418268 0 io_out[9]
rlabel metal2 125757 340 125757 340 0 la_data_in[0]
rlabel metal2 480562 2098 480562 2098 0 la_data_in[100]
rlabel metal2 484058 2030 484058 2030 0 la_data_in[101]
rlabel metal2 487646 2166 487646 2166 0 la_data_in[102]
rlabel metal2 490951 340 490951 340 0 la_data_in[103]
rlabel metal2 494408 16560 494408 16560 0 la_data_in[104]
rlabel metal3 353671 35292 353671 35292 0 la_data_in[105]
rlabel metal2 501814 1962 501814 1962 0 la_data_in[106]
rlabel metal2 505264 16560 505264 16560 0 la_data_in[107]
rlabel metal2 508392 16560 508392 16560 0 la_data_in[108]
rlabel metal2 512249 340 512249 340 0 la_data_in[109]
rlabel metal2 161322 1928 161322 1928 0 la_data_in[10]
rlabel metal2 515791 340 515791 340 0 la_data_in[110]
rlabel metal2 519570 1911 519570 1911 0 la_data_in[111]
rlabel metal2 523066 1996 523066 1996 0 la_data_in[112]
rlabel metal2 526654 2064 526654 2064 0 la_data_in[113]
rlabel metal2 530051 340 530051 340 0 la_data_in[114]
rlabel metal2 533232 16560 533232 16560 0 la_data_in[115]
rlabel metal1 398544 18598 398544 18598 0 la_data_in[116]
rlabel metal2 540631 340 540631 340 0 la_data_in[117]
rlabel metal2 544088 16560 544088 16560 0 la_data_in[118]
rlabel metal1 380558 36822 380558 36822 0 la_data_in[119]
rlabel metal2 164910 1962 164910 1962 0 la_data_in[11]
rlabel metal2 551257 340 551257 340 0 la_data_in[120]
rlabel metal2 554891 340 554891 340 0 la_data_in[121]
rlabel metal2 558072 16560 558072 16560 0 la_data_in[122]
rlabel metal2 561890 16560 561890 16560 0 la_data_in[123]
rlabel metal2 565425 340 565425 340 0 la_data_in[124]
rlabel metal2 568921 340 568921 340 0 la_data_in[125]
rlabel metal2 572746 1843 572746 1843 0 la_data_in[126]
rlabel metal2 576334 2574 576334 2574 0 la_data_in[127]
rlabel metal2 168406 1231 168406 1231 0 la_data_in[12]
rlabel metal2 171580 16560 171580 16560 0 la_data_in[13]
rlabel metal2 175398 16560 175398 16560 0 la_data_in[14]
rlabel metal2 178841 340 178841 340 0 la_data_in[15]
rlabel metal2 182475 340 182475 340 0 la_data_in[16]
rlabel metal2 186162 1911 186162 1911 0 la_data_in[17]
rlabel metal2 189750 1826 189750 1826 0 la_data_in[18]
rlabel metal2 193246 1758 193246 1758 0 la_data_in[19]
rlabel metal2 129161 340 129161 340 0 la_data_in[1]
rlabel metal2 196834 3627 196834 3627 0 la_data_in[20]
rlabel metal2 200330 2132 200330 2132 0 la_data_in[21]
rlabel metal2 203918 2030 203918 2030 0 la_data_in[22]
rlabel metal2 207414 2064 207414 2064 0 la_data_in[23]
rlabel metal2 211002 2098 211002 2098 0 la_data_in[24]
rlabel metal2 214498 1622 214498 1622 0 la_data_in[25]
rlabel metal2 218086 3627 218086 3627 0 la_data_in[26]
rlabel metal2 221345 340 221345 340 0 la_data_in[27]
rlabel metal2 213210 18156 213210 18156 0 la_data_in[28]
rlabel metal2 228521 340 228521 340 0 la_data_in[29]
rlabel metal2 132986 1724 132986 1724 0 la_data_in[2]
rlabel metal2 232063 340 232063 340 0 la_data_in[30]
rlabel metal2 235290 16560 235290 16560 0 la_data_in[31]
rlabel metal2 239062 16560 239062 16560 0 la_data_in[32]
rlabel metal2 242926 25932 242926 25932 0 la_data_in[33]
rlabel metal2 246422 2030 246422 2030 0 la_data_in[34]
rlabel metal2 249918 16560 249918 16560 0 la_data_in[35]
rlabel metal2 253506 1911 253506 1911 0 la_data_in[36]
rlabel metal2 257094 1860 257094 1860 0 la_data_in[37]
rlabel metal2 260682 2183 260682 2183 0 la_data_in[38]
rlabel metal2 264178 2115 264178 2115 0 la_data_in[39]
rlabel metal2 136482 2030 136482 2030 0 la_data_in[3]
rlabel metal2 267766 2047 267766 2047 0 la_data_in[40]
rlabel metal2 271262 1758 271262 1758 0 la_data_in[41]
rlabel metal2 274850 1792 274850 1792 0 la_data_in[42]
rlabel metal2 278346 1979 278346 1979 0 la_data_in[43]
rlabel metal2 281743 340 281743 340 0 la_data_in[44]
rlabel metal2 285239 340 285239 340 0 la_data_in[45]
rlabel metal2 289018 1826 289018 1826 0 la_data_in[46]
rlabel metal2 292606 1860 292606 1860 0 la_data_in[47]
rlabel metal2 296102 2234 296102 2234 0 la_data_in[48]
rlabel metal2 299690 3458 299690 3458 0 la_data_in[49]
rlabel metal2 139833 340 139833 340 0 la_data_in[4]
rlabel metal2 303186 3543 303186 3543 0 la_data_in[50]
rlabel metal2 306774 3220 306774 3220 0 la_data_in[51]
rlabel metal2 310033 340 310033 340 0 la_data_in[52]
rlabel metal2 313582 16560 313582 16560 0 la_data_in[53]
rlabel metal2 317354 1860 317354 1860 0 la_data_in[54]
rlabel metal2 320705 340 320705 340 0 la_data_in[55]
rlabel metal2 324438 1775 324438 1775 0 la_data_in[56]
rlabel metal2 328026 3560 328026 3560 0 la_data_in[57]
rlabel metal2 331423 340 331423 340 0 la_data_in[58]
rlabel metal2 334873 340 334873 340 0 la_data_in[59]
rlabel metal2 143566 3627 143566 3627 0 la_data_in[5]
rlabel metal2 338422 16560 338422 16560 0 la_data_in[60]
rlabel metal2 256634 28526 256634 28526 0 la_data_in[61]
rlabel metal2 345545 340 345545 340 0 la_data_in[62]
rlabel metal2 349186 19891 349186 19891 0 la_data_in[63]
rlabel metal2 352866 4104 352866 4104 0 la_data_in[64]
rlabel metal2 356362 3475 356362 3475 0 la_data_in[65]
rlabel metal2 359713 340 359713 340 0 la_data_in[66]
rlabel metal1 281014 24378 281014 24378 0 la_data_in[67]
rlabel metal2 367034 4070 367034 4070 0 la_data_in[68]
rlabel metal2 370622 3407 370622 3407 0 la_data_in[69]
rlabel metal2 146740 16560 146740 16560 0 la_data_in[6]
rlabel metal3 286925 21556 286925 21556 0 la_data_in[70]
rlabel metal2 256358 28934 256358 28934 0 la_data_in[71]
rlabel metal2 253322 29682 253322 29682 0 la_data_in[72]
rlabel metal2 384553 340 384553 340 0 la_data_in[73]
rlabel metal2 388286 4818 388286 4818 0 la_data_in[74]
rlabel metal2 391874 4784 391874 4784 0 la_data_in[75]
rlabel metal2 395048 16560 395048 16560 0 la_data_in[76]
rlabel metal2 398958 1775 398958 1775 0 la_data_in[77]
rlabel metal2 402546 2642 402546 2642 0 la_data_in[78]
rlabel metal2 406042 4036 406042 4036 0 la_data_in[79]
rlabel metal2 150650 2098 150650 2098 0 la_data_in[7]
rlabel metal2 409630 3339 409630 3339 0 la_data_in[80]
rlabel metal2 253506 30600 253506 30600 0 la_data_in[81]
rlabel metal2 416714 1860 416714 1860 0 la_data_in[82]
rlabel metal1 311558 9146 311558 9146 0 la_data_in[83]
rlabel metal2 423798 2659 423798 2659 0 la_data_in[84]
rlabel metal2 427057 340 427057 340 0 la_data_in[85]
rlabel metal2 253598 30600 253598 30600 0 la_data_in[86]
rlabel metal2 253230 29988 253230 29988 0 la_data_in[87]
rlabel metal2 437966 3322 437966 3322 0 la_data_in[88]
rlabel metal2 441554 1860 441554 1860 0 la_data_in[89]
rlabel metal2 154001 340 154001 340 0 la_data_in[8]
rlabel metal2 445050 4699 445050 4699 0 la_data_in[90]
rlabel metal2 448638 1163 448638 1163 0 la_data_in[91]
rlabel metal2 451897 340 451897 340 0 la_data_in[92]
rlabel metal1 330740 12070 330740 12070 0 la_data_in[93]
rlabel metal1 332534 12002 332534 12002 0 la_data_in[94]
rlabel metal2 462569 340 462569 340 0 la_data_in[95]
rlabel metal2 466065 340 466065 340 0 la_data_in[96]
rlabel metal2 469890 7504 469890 7504 0 la_data_in[97]
rlabel metal1 340400 14586 340400 14586 0 la_data_in[98]
rlabel metal2 476737 340 476737 340 0 la_data_in[99]
rlabel metal2 157596 16560 157596 16560 0 la_data_in[9]
rlabel metal1 153640 17510 153640 17510 0 la_data_out[0]
rlabel metal2 481758 3271 481758 3271 0 la_data_out[100]
rlabel metal2 485254 4648 485254 4648 0 la_data_out[101]
rlabel metal2 488566 20401 488566 20401 0 la_data_out[102]
rlabel metal1 339503 4862 339503 4862 0 la_data_out[103]
rlabel metal2 495689 340 495689 340 0 la_data_out[104]
rlabel metal2 499185 340 499185 340 0 la_data_out[105]
rlabel metal2 503010 3288 503010 3288 0 la_data_out[106]
rlabel metal2 506506 11618 506506 11618 0 la_data_out[107]
rlabel metal1 359996 7650 359996 7650 0 la_data_out[108]
rlabel metal2 513491 340 513491 340 0 la_data_out[109]
rlabel metal2 162518 3356 162518 3356 0 la_data_out[10]
rlabel metal2 516672 16560 516672 16560 0 la_data_out[110]
rlabel metal2 520529 340 520529 340 0 la_data_out[111]
rlabel metal2 524025 340 524025 340 0 la_data_out[112]
rlabel metal2 527850 6042 527850 6042 0 la_data_out[113]
rlabel metal2 531346 1911 531346 1911 0 la_data_out[114]
rlabel metal2 534697 340 534697 340 0 la_data_out[115]
rlabel metal2 538331 340 538331 340 0 la_data_out[116]
rlabel metal2 541006 18973 541006 18973 0 la_data_out[117]
rlabel metal2 545146 21047 545146 21047 0 la_data_out[118]
rlabel metal3 381409 8908 381409 8908 0 la_data_out[119]
rlabel metal2 166106 6076 166106 6076 0 la_data_out[11]
rlabel metal2 552368 16560 552368 16560 0 la_data_out[120]
rlabel metal2 487830 17306 487830 17306 0 la_data_out[121]
rlabel metal2 559537 340 559537 340 0 la_data_out[122]
rlabel metal2 563171 340 563171 340 0 la_data_out[123]
rlabel metal2 566858 2591 566858 2591 0 la_data_out[124]
rlabel metal3 392311 25636 392311 25636 0 la_data_out[125]
rlabel metal2 573751 340 573751 340 0 la_data_out[126]
rlabel metal2 577201 340 577201 340 0 la_data_out[127]
rlabel metal2 169602 1894 169602 1894 0 la_data_out[12]
rlabel metal2 173190 1928 173190 1928 0 la_data_out[13]
rlabel metal2 176686 3627 176686 3627 0 la_data_out[14]
rlabel metal2 179446 19653 179446 19653 0 la_data_out[15]
rlabel metal2 183678 16560 183678 16560 0 la_data_out[16]
rlabel metal2 187121 340 187121 340 0 la_data_out[17]
rlabel metal2 190854 2234 190854 2234 0 la_data_out[18]
rlabel metal2 193706 19653 193706 19653 0 la_data_out[19]
rlabel metal3 155365 18700 155365 18700 0 la_data_out[1]
rlabel metal2 197938 1792 197938 1792 0 la_data_out[20]
rlabel metal2 201526 2200 201526 2200 0 la_data_out[21]
rlabel metal2 205114 2166 205114 2166 0 la_data_out[22]
rlabel metal2 208610 1758 208610 1758 0 la_data_out[23]
rlabel metal2 212198 1860 212198 1860 0 la_data_out[24]
rlabel metal2 215694 1894 215694 1894 0 la_data_out[25]
rlabel metal2 219282 1996 219282 1996 0 la_data_out[26]
rlabel metal2 222778 3560 222778 3560 0 la_data_out[27]
rlabel metal2 226366 1843 226366 1843 0 la_data_out[28]
rlabel metal2 229862 3390 229862 3390 0 la_data_out[29]
rlabel metal2 134182 2132 134182 2132 0 la_data_out[2]
rlabel metal2 233450 3203 233450 3203 0 la_data_out[30]
rlabel metal2 236801 340 236801 340 0 la_data_out[31]
rlabel metal2 240343 340 240343 340 0 la_data_out[32]
rlabel metal2 243570 16560 243570 16560 0 la_data_out[33]
rlabel metal2 247342 16560 247342 16560 0 la_data_out[34]
rlabel metal2 251206 1843 251206 1843 0 la_data_out[35]
rlabel metal2 254465 340 254465 340 0 la_data_out[36]
rlabel metal2 258198 16560 258198 16560 0 la_data_out[37]
rlabel metal1 225860 21658 225860 21658 0 la_data_out[38]
rlabel metal2 265183 340 265183 340 0 la_data_out[39]
rlabel metal2 137441 340 137441 340 0 la_data_out[3]
rlabel metal2 268633 340 268633 340 0 la_data_out[40]
rlabel metal2 272458 6824 272458 6824 0 la_data_out[41]
rlabel metal2 276046 1911 276046 1911 0 la_data_out[42]
rlabel metal2 279305 340 279305 340 0 la_data_out[43]
rlabel metal3 237935 13260 237935 13260 0 la_data_out[44]
rlabel metal2 286166 16560 286166 16560 0 la_data_out[45]
rlabel metal2 290214 3186 290214 3186 0 la_data_out[46]
rlabel metal2 293473 340 293473 340 0 la_data_out[47]
rlabel metal1 245916 10506 245916 10506 0 la_data_out[48]
rlabel metal2 300794 1860 300794 1860 0 la_data_out[49]
rlabel metal2 141036 16560 141036 16560 0 la_data_out[4]
rlabel metal2 304145 340 304145 340 0 la_data_out[50]
rlabel metal2 307970 2744 307970 2744 0 la_data_out[51]
rlabel metal2 311466 3424 311466 3424 0 la_data_out[52]
rlabel metal2 315054 4172 315054 4172 0 la_data_out[53]
rlabel metal2 318313 340 318313 340 0 la_data_out[54]
rlabel metal3 258911 14620 258911 14620 0 la_data_out[55]
rlabel metal2 325634 1860 325634 1860 0 la_data_out[56]
rlabel metal2 328985 340 328985 340 0 la_data_out[57]
rlabel metal2 332718 7368 332718 7368 0 la_data_out[58]
rlabel metal1 266248 15062 266248 15062 0 la_data_out[59]
rlabel metal1 144164 11662 144164 11662 0 la_data_out[5]
rlabel metal2 339703 340 339703 340 0 la_data_out[60]
rlabel metal2 343153 340 343153 340 0 la_data_out[61]
rlabel metal2 346978 7640 346978 7640 0 la_data_out[62]
rlabel metal2 350474 4138 350474 4138 0 la_data_out[63]
rlabel metal2 353825 340 353825 340 0 la_data_out[64]
rlabel metal3 277817 32708 277817 32708 0 la_data_out[65]
rlabel metal1 280048 9486 280048 9486 0 la_data_out[66]
rlabel metal2 364504 16560 364504 16560 0 la_data_out[67]
rlabel metal2 368230 2676 368230 2676 0 la_data_out[68]
rlabel metal2 371489 340 371489 340 0 la_data_out[69]
rlabel metal2 148113 340 148113 340 0 la_data_out[6]
rlabel metal2 375314 1860 375314 1860 0 la_data_out[70]
rlabel metal2 378665 340 378665 340 0 la_data_out[71]
rlabel metal1 291456 24310 291456 24310 0 la_data_out[72]
rlabel metal2 385526 16560 385526 16560 0 la_data_out[73]
rlabel metal2 389482 6314 389482 6314 0 la_data_out[74]
rlabel metal2 392833 340 392833 340 0 la_data_out[75]
rlabel metal2 396329 340 396329 340 0 la_data_out[76]
rlabel metal2 400154 1860 400154 1860 0 la_data_out[77]
rlabel metal2 403650 3356 403650 3356 0 la_data_out[78]
rlabel metal2 407238 1775 407238 1775 0 la_data_out[79]
rlabel metal2 151846 21920 151846 21920 0 la_data_out[7]
rlabel metal2 410826 7419 410826 7419 0 la_data_out[80]
rlabel metal1 308660 16354 308660 16354 0 la_data_out[81]
rlabel metal2 417673 340 417673 340 0 la_data_out[82]
rlabel metal2 421169 340 421169 340 0 la_data_out[83]
rlabel metal2 424994 1860 424994 1860 0 la_data_out[84]
rlabel metal2 428490 8099 428490 8099 0 la_data_out[85]
rlabel metal1 318320 16150 318320 16150 0 la_data_out[86]
rlabel metal2 435337 340 435337 340 0 la_data_out[87]
rlabel metal1 321770 16014 321770 16014 0 la_data_out[88]
rlabel metal2 441646 19041 441646 19041 0 la_data_out[89]
rlabel metal2 155020 16560 155020 16560 0 la_data_out[8]
rlabel metal2 446009 340 446009 340 0 la_data_out[90]
rlabel metal2 449834 1860 449834 1860 0 la_data_out[91]
rlabel metal1 329774 14790 329774 14790 0 la_data_out[92]
rlabel metal1 331522 14722 331522 14722 0 la_data_out[93]
rlabel metal1 333592 9078 333592 9078 0 la_data_out[94]
rlabel metal2 463726 17018 463726 17018 0 la_data_out[95]
rlabel metal2 466486 17171 466486 17171 0 la_data_out[96]
rlabel metal2 470849 340 470849 340 0 la_data_out[97]
rlabel metal2 474391 340 474391 340 0 la_data_out[98]
rlabel metal3 342401 17340 342401 17340 0 la_data_out[99]
rlabel metal2 158930 1894 158930 1894 0 la_data_out[9]
rlabel metal3 154215 17340 154215 17340 0 la_oenb[0]
rlabel metal2 482862 4682 482862 4682 0 la_oenb[100]
rlabel metal2 486450 5362 486450 5362 0 la_oenb[101]
rlabel metal2 489946 1775 489946 1775 0 la_oenb[102]
rlabel metal2 493297 340 493297 340 0 la_oenb[103]
rlabel metal3 353165 24276 353165 24276 0 la_oenb[104]
rlabel metal2 500618 6756 500618 6756 0 la_oenb[105]
rlabel metal2 503969 340 503969 340 0 la_oenb[106]
rlabel metal2 507465 340 507465 340 0 la_oenb[107]
rlabel metal2 468510 10880 468510 10880 0 la_oenb[108]
rlabel metal2 514786 1911 514786 1911 0 la_oenb[109]
rlabel metal2 163714 3271 163714 3271 0 la_oenb[10]
rlabel metal2 518137 340 518137 340 0 la_oenb[110]
rlabel metal2 521771 340 521771 340 0 la_oenb[111]
rlabel metal2 524446 17035 524446 17035 0 la_oenb[112]
rlabel metal2 528809 340 528809 340 0 la_oenb[113]
rlabel metal2 532351 340 532351 340 0 la_oenb[114]
rlabel metal1 374118 17374 374118 17374 0 la_oenb[115]
rlabel metal2 539626 1911 539626 1911 0 la_oenb[116]
rlabel metal2 542977 340 542977 340 0 la_oenb[117]
rlabel metal2 546611 340 546611 340 0 la_oenb[118]
rlabel metal2 549792 16560 549792 16560 0 la_oenb[119]
rlabel metal2 167210 2591 167210 2591 0 la_oenb[11]
rlabel metal2 553794 3254 553794 3254 0 la_oenb[120]
rlabel metal2 557145 340 557145 340 0 la_oenb[121]
rlabel metal2 560641 340 560641 340 0 la_oenb[122]
rlabel metal2 564466 17058 564466 17058 0 la_oenb[123]
rlabel metal2 567817 340 567817 340 0 la_oenb[124]
rlabel metal1 393484 7582 393484 7582 0 la_oenb[125]
rlabel metal1 395324 10302 395324 10302 0 la_oenb[126]
rlabel metal2 578634 6722 578634 6722 0 la_oenb[127]
rlabel metal2 170561 340 170561 340 0 la_oenb[12]
rlabel metal2 174294 1894 174294 1894 0 la_oenb[13]
rlabel metal1 177284 11730 177284 11730 0 la_oenb[14]
rlabel metal2 181233 340 181233 340 0 la_oenb[15]
rlabel metal2 184966 1962 184966 1962 0 la_oenb[16]
rlabel metal2 188554 2948 188554 2948 0 la_oenb[17]
rlabel metal2 192050 6382 192050 6382 0 la_oenb[18]
rlabel metal2 195401 340 195401 340 0 la_oenb[19]
rlabel metal2 131553 340 131553 340 0 la_oenb[1]
rlabel metal2 199134 1826 199134 1826 0 la_oenb[20]
rlabel metal2 202722 1860 202722 1860 0 la_oenb[21]
rlabel metal1 196420 10302 196420 10302 0 la_oenb[22]
rlabel metal2 209806 1588 209806 1588 0 la_oenb[23]
rlabel metal2 213394 1928 213394 1928 0 la_oenb[24]
rlabel metal2 216890 3594 216890 3594 0 la_oenb[25]
rlabel metal1 204332 9418 204332 9418 0 la_oenb[26]
rlabel metal2 223783 340 223783 340 0 la_oenb[27]
rlabel metal2 227562 1894 227562 1894 0 la_oenb[28]
rlabel metal2 230782 16560 230782 16560 0 la_oenb[29]
rlabel metal2 135286 13624 135286 13624 0 la_oenb[2]
rlabel metal2 234646 1962 234646 1962 0 la_oenb[30]
rlabel metal2 237905 340 237905 340 0 la_oenb[31]
rlabel metal1 215464 9350 215464 9350 0 la_oenb[32]
rlabel metal2 244766 16560 244766 16560 0 la_oenb[33]
rlabel metal2 248623 340 248623 340 0 la_oenb[34]
rlabel metal2 252402 1894 252402 1894 0 la_oenb[35]
rlabel metal2 255622 16560 255622 16560 0 la_oenb[36]
rlabel metal2 259486 23280 259486 23280 0 la_oenb[37]
rlabel metal2 262745 340 262745 340 0 la_oenb[38]
rlabel metal3 228735 36516 228735 36516 0 la_oenb[39]
rlabel metal2 138874 1911 138874 1911 0 la_oenb[3]
rlabel metal2 270066 3526 270066 3526 0 la_oenb[40]
rlabel metal2 273463 340 273463 340 0 la_oenb[41]
rlabel metal2 276959 340 276959 340 0 la_oenb[42]
rlabel metal1 236256 19074 236256 19074 0 la_oenb[43]
rlabel metal2 284326 1911 284326 1911 0 la_oenb[44]
rlabel metal2 287585 340 287585 340 0 la_oenb[45]
rlabel metal2 291226 17783 291226 17783 0 la_oenb[46]
rlabel metal2 293986 17749 293986 17749 0 la_oenb[47]
rlabel metal2 298303 340 298303 340 0 la_oenb[48]
rlabel metal2 301753 340 301753 340 0 la_oenb[49]
rlabel metal2 142462 1996 142462 1996 0 la_oenb[4]
rlabel metal1 250010 18870 250010 18870 0 la_oenb[50]
rlabel metal2 309074 1860 309074 1860 0 la_oenb[51]
rlabel metal2 312425 340 312425 340 0 la_oenb[52]
rlabel metal1 255530 17170 255530 17170 0 la_oenb[53]
rlabel metal3 257071 37876 257071 37876 0 la_oenb[54]
rlabel metal2 323334 2710 323334 2710 0 la_oenb[55]
rlabel metal2 326593 340 326593 340 0 la_oenb[56]
rlabel metal2 329866 17681 329866 17681 0 la_oenb[57]
rlabel metal2 333914 1860 333914 1860 0 la_oenb[58]
rlabel metal2 337265 340 337265 340 0 la_oenb[59]
rlabel metal2 145721 340 145721 340 0 la_oenb[5]
rlabel metal2 340952 16560 340952 16560 0 la_oenb[60]
rlabel metal1 271078 9622 271078 9622 0 la_oenb[61]
rlabel metal2 347944 16560 347944 16560 0 la_oenb[62]
rlabel metal2 351433 340 351433 340 0 la_oenb[63]
rlabel metal3 276851 15980 276851 15980 0 la_oenb[64]
rlabel metal2 358754 1860 358754 1860 0 la_oenb[65]
rlabel metal2 362105 340 362105 340 0 la_oenb[66]
rlabel metal2 365792 16560 365792 16560 0 la_oenb[67]
rlabel metal2 368506 21115 368506 21115 0 la_oenb[68]
rlabel metal2 372784 16560 372784 16560 0 la_oenb[69]
rlabel metal2 149316 16560 149316 16560 0 la_oenb[6]
rlabel metal2 376273 340 376273 340 0 la_oenb[70]
rlabel metal2 379769 340 379769 340 0 la_oenb[71]
rlabel metal2 383594 1860 383594 1860 0 la_oenb[72]
rlabel metal2 386945 340 386945 340 0 la_oenb[73]
rlabel metal2 390632 16560 390632 16560 0 la_oenb[74]
rlabel metal2 253690 30260 253690 30260 0 la_oenb[75]
rlabel metal2 255898 35224 255898 35224 0 la_oenb[76]
rlabel metal2 401113 340 401113 340 0 la_oenb[77]
rlabel metal2 404609 340 404609 340 0 la_oenb[78]
rlabel metal2 408434 1860 408434 1860 0 la_oenb[79]
rlabel metal2 152490 16560 152490 16560 0 la_oenb[7]
rlabel metal2 253782 33966 253782 33966 0 la_oenb[80]
rlabel metal1 310362 20162 310362 20162 0 la_oenb[81]
rlabel metal2 418777 340 418777 340 0 la_oenb[82]
rlabel metal2 422326 18327 422326 18327 0 la_oenb[83]
rlabel metal2 425953 340 425953 340 0 la_oenb[84]
rlabel metal2 429449 340 429449 340 0 la_oenb[85]
rlabel metal2 433274 2064 433274 2064 0 la_oenb[86]
rlabel metal1 326048 18666 326048 18666 0 la_oenb[87]
rlabel metal2 440358 1231 440358 1231 0 la_oenb[88]
rlabel metal2 443617 340 443617 340 0 la_oenb[89]
rlabel metal2 156393 340 156393 340 0 la_oenb[8]
rlabel metal2 447442 7606 447442 7606 0 la_oenb[90]
rlabel metal2 450938 1588 450938 1588 0 la_oenb[91]
rlabel metal2 454289 340 454289 340 0 la_oenb[92]
rlabel metal2 458114 1860 458114 1860 0 la_oenb[93]
rlabel metal2 461610 2132 461610 2132 0 la_oenb[94]
rlabel metal2 465198 6790 465198 6790 0 la_oenb[95]
rlabel metal2 468694 1843 468694 1843 0 la_oenb[96]
rlabel metal1 365332 21590 365332 21590 0 la_oenb[97]
rlabel metal1 341228 38114 341228 38114 0 la_oenb[98]
rlabel metal2 479366 1860 479366 1860 0 la_oenb[99]
rlabel metal2 160126 2574 160126 2574 0 la_oenb[9]
rlabel metal3 156730 292332 156730 292332 0 mprj/c0_clk
rlabel metal2 137310 236980 137310 236980 0 mprj/c0_dbg_pc\[0\]
rlabel metal3 156638 329324 156638 329324 0 mprj/c0_dbg_pc\[10\]
rlabel metal2 154974 331755 154974 331755 0 mprj/c0_dbg_pc\[11\]
rlabel metal2 154790 334407 154790 334407 0 mprj/c0_dbg_pc\[12\]
rlabel metal2 155066 337127 155066 337127 0 mprj/c0_dbg_pc\[13\]
rlabel metal2 154974 339983 154974 339983 0 mprj/c0_dbg_pc\[14\]
rlabel metal2 154882 342669 154882 342669 0 mprj/c0_dbg_pc\[15\]
rlabel metal2 133262 236946 133262 236946 0 mprj/c0_dbg_pc\[1\]
rlabel metal1 154100 303654 154100 303654 0 mprj/c0_dbg_pc\[2\]
rlabel metal2 155066 307105 155066 307105 0 mprj/c0_dbg_pc\[3\]
rlabel metal2 154974 310777 154974 310777 0 mprj/c0_dbg_pc\[4\]
rlabel metal1 155388 306510 155388 306510 0 mprj/c0_dbg_pc\[5\]
rlabel metal2 154790 316795 154790 316795 0 mprj/c0_dbg_pc\[6\]
rlabel metal2 154882 320501 154882 320501 0 mprj/c0_dbg_pc\[7\]
rlabel metal3 156040 323884 156040 323884 0 mprj/c0_dbg_pc\[8\]
rlabel metal2 154974 326247 154974 326247 0 mprj/c0_dbg_pc\[9\]
rlabel metal2 138874 248812 138874 248812 0 mprj/c0_dbg_r0\[0\]
rlabel metal2 154882 329103 154882 329103 0 mprj/c0_dbg_r0\[10\]
rlabel metal3 156960 332316 156960 332316 0 mprj/c0_dbg_r0\[11\]
rlabel metal3 157006 335036 157006 335036 0 mprj/c0_dbg_r0\[12\]
rlabel metal2 154882 337365 154882 337365 0 mprj/c0_dbg_r0\[13\]
rlabel metal2 133262 315282 133262 315282 0 mprj/c0_dbg_r0\[14\]
rlabel metal2 115138 316268 115138 316268 0 mprj/c0_dbg_r0\[15\]
rlabel metal3 109940 192285 109940 192285 0 mprj/c0_dbg_r0\[1\]
rlabel metal2 115322 252620 115322 252620 0 mprj/c0_dbg_r0\[2\]
rlabel metal2 154974 307921 154974 307921 0 mprj/c0_dbg_r0\[3\]
rlabel metal2 155066 310811 155066 310811 0 mprj/c0_dbg_r0\[4\]
rlabel metal2 154882 313871 154882 313871 0 mprj/c0_dbg_r0\[5\]
rlabel via2 154974 317645 154974 317645 0 mprj/c0_dbg_r0\[6\]
rlabel metal2 154974 320671 154974 320671 0 mprj/c0_dbg_r0\[7\]
rlabel metal2 137494 287130 137494 287130 0 mprj/c0_dbg_r0\[8\]
rlabel metal2 154882 326417 154882 326417 0 mprj/c0_dbg_r0\[9\]
rlabel metal2 116610 231778 116610 231778 0 mprj/c0_disable
rlabel metal2 116702 240822 116702 240822 0 mprj/c0_i_core_int_sreg\[0\]
rlabel metal1 153778 328746 153778 328746 0 mprj/c0_i_core_int_sreg\[10\]
rlabel metal2 154790 331551 154790 331551 0 mprj/c0_i_core_int_sreg\[11\]
rlabel metal1 155066 311202 155066 311202 0 mprj/c0_i_core_int_sreg\[12\]
rlabel metal2 139150 311236 139150 311236 0 mprj/c0_i_core_int_sreg\[13\]
rlabel metal2 137310 316064 137310 316064 0 mprj/c0_i_core_int_sreg\[14\]
rlabel metal2 115874 320552 115874 320552 0 mprj/c0_i_core_int_sreg\[15\]
rlabel metal2 140254 247078 140254 247078 0 mprj/c0_i_core_int_sreg\[1\]
rlabel metal2 116794 253232 116794 253232 0 mprj/c0_i_core_int_sreg\[2\]
rlabel metal3 156362 308108 156362 308108 0 mprj/c0_i_core_int_sreg\[3\]
rlabel metal2 154882 311083 154882 311083 0 mprj/c0_i_core_int_sreg\[4\]
rlabel metal2 154790 313973 154790 313973 0 mprj/c0_i_core_int_sreg\[5\]
rlabel metal2 154882 317815 154882 317815 0 mprj/c0_i_core_int_sreg\[6\]
rlabel metal2 133446 281588 133446 281588 0 mprj/c0_i_core_int_sreg\[7\]
rlabel metal2 154974 324377 154974 324377 0 mprj/c0_i_core_int_sreg\[8\]
rlabel metal2 154790 327233 154790 327233 0 mprj/c0_i_core_int_sreg\[9\]
rlabel metal3 109940 171885 109940 171885 0 mprj/c0_i_irq
rlabel metal3 109940 172263 109940 172263 0 mprj/c0_i_mc_core_int
rlabel metal2 119370 233206 119370 233206 0 mprj/c0_i_mem_ack
rlabel metal2 115230 240754 115230 240754 0 mprj/c0_i_mem_data\[0\]
rlabel metal2 154974 330089 154974 330089 0 mprj/c0_i_mem_data\[10\]
rlabel via2 154606 332843 154606 332843 0 mprj/c0_i_mem_data\[11\]
rlabel metal2 154974 335461 154974 335461 0 mprj/c0_i_mem_data\[12\]
rlabel metal2 140622 310148 140622 310148 0 mprj/c0_i_mem_data\[13\]
rlabel metal2 119922 314908 119922 314908 0 mprj/c0_i_mem_data\[14\]
rlabel metal2 115230 321028 115230 321028 0 mprj/c0_i_mem_data\[15\]
rlabel metal2 119462 247656 119462 247656 0 mprj/c0_i_mem_data\[1\]
rlabel metal2 119554 253538 119554 253538 0 mprj/c0_i_mem_data\[2\]
rlabel metal2 154882 308091 154882 308091 0 mprj/c0_i_mem_data\[3\]
rlabel metal2 154790 311117 154790 311117 0 mprj/c0_i_mem_data\[4\]
rlabel metal2 155618 313021 155618 313021 0 mprj/c0_i_mem_data\[5\]
rlabel metal2 139058 277134 139058 277134 0 mprj/c0_i_mem_data\[6\]
rlabel metal2 155066 320807 155066 320807 0 mprj/c0_i_mem_data\[7\]
rlabel metal2 113206 260749 113206 260749 0 mprj/c0_i_mem_data\[8\]
rlabel metal2 154974 327335 154974 327335 0 mprj/c0_i_mem_data\[9\]
rlabel metal2 120750 233274 120750 233274 0 mprj/c0_i_mem_exception
rlabel metal3 109940 185485 109940 185485 0 mprj/c0_i_req_data\[0\]
rlabel metal2 154882 330191 154882 330191 0 mprj/c0_i_req_data\[10\]
rlabel metal3 156086 333132 156086 333132 0 mprj/c0_i_req_data\[11\]
rlabel metal2 133538 307768 133538 307768 0 mprj/c0_i_req_data\[12\]
rlabel metal2 154974 338453 154974 338453 0 mprj/c0_i_req_data\[13\]
rlabel metal2 117162 317390 117162 317390 0 mprj/c0_i_req_data\[14\]
rlabel metal2 154606 343927 154606 343927 0 mprj/c0_i_req_data\[15\]
rlabel metal3 154951 345508 154951 345508 0 mprj/c0_i_req_data\[16\]
rlabel metal2 154974 345559 154974 345559 0 mprj/c0_i_req_data\[17\]
rlabel metal2 155066 345661 155066 345661 0 mprj/c0_i_req_data\[18\]
rlabel metal2 154882 346069 154882 346069 0 mprj/c0_i_req_data\[19\]
rlabel metal2 120842 247724 120842 247724 0 mprj/c0_i_req_data\[1\]
rlabel metal2 154974 346647 154974 346647 0 mprj/c0_i_req_data\[20\]
rlabel metal2 154606 346715 154606 346715 0 mprj/c0_i_req_data\[21\]
rlabel metal2 154882 346953 154882 346953 0 mprj/c0_i_req_data\[22\]
rlabel metal2 155066 347021 155066 347021 0 mprj/c0_i_req_data\[23\]
rlabel metal2 154974 347429 154974 347429 0 mprj/c0_i_req_data\[24\]
rlabel metal2 154974 348007 154974 348007 0 mprj/c0_i_req_data\[25\]
rlabel metal2 154790 348109 154790 348109 0 mprj/c0_i_req_data\[26\]
rlabel metal2 154882 348313 154882 348313 0 mprj/c0_i_req_data\[27\]
rlabel metal2 155066 348347 155066 348347 0 mprj/c0_i_req_data\[28\]
rlabel metal3 156822 349180 156822 349180 0 mprj/c0_i_req_data\[29\]
rlabel metal2 114126 254524 114126 254524 0 mprj/c0_i_req_data\[2\]
rlabel metal2 154882 349299 154882 349299 0 mprj/c0_i_req_data\[30\]
rlabel metal2 154974 349469 154974 349469 0 mprj/c0_i_req_data\[31\]
rlabel metal2 154790 308295 154790 308295 0 mprj/c0_i_req_data\[3\]
rlabel metal1 153686 311882 153686 311882 0 mprj/c0_i_req_data\[4\]
rlabel metal2 154974 314925 154974 314925 0 mprj/c0_i_req_data\[5\]
rlabel metal2 122314 276726 122314 276726 0 mprj/c0_i_req_data\[6\]
rlabel metal2 122406 281146 122406 281146 0 mprj/c0_i_req_data\[7\]
rlabel metal2 122498 288490 122498 288490 0 mprj/c0_i_req_data\[8\]
rlabel metal2 154882 327437 154882 327437 0 mprj/c0_i_req_data\[9\]
rlabel metal3 109940 174605 109940 174605 0 mprj/c0_i_req_data_valid
rlabel metal2 122130 235348 122130 235348 0 mprj/c0_o_c_data_page
rlabel metal3 109940 176441 109940 176441 0 mprj/c0_o_c_instr_long
rlabel metal2 140162 239190 140162 239190 0 mprj/c0_o_c_instr_page
rlabel metal2 120934 250920 120934 250920 0 mprj/c0_o_icache_flush
rlabel metal1 131330 193834 131330 193834 0 mprj/c0_o_instr_long_addr\[0\]
rlabel metal2 137402 248438 137402 248438 0 mprj/c0_o_instr_long_addr\[1\]
rlabel metal3 156868 305660 156868 305660 0 mprj/c0_o_instr_long_addr\[2\]
rlabel metal2 155066 308397 155066 308397 0 mprj/c0_o_instr_long_addr\[3\]
rlabel via2 154974 312171 154974 312171 0 mprj/c0_o_instr_long_addr\[4\]
rlabel metal2 154790 315095 154790 315095 0 mprj/c0_o_instr_long_addr\[5\]
rlabel metal2 119738 279106 119738 279106 0 mprj/c0_o_instr_long_addr\[6\]
rlabel metal2 116978 283594 116978 283594 0 mprj/c0_o_instr_long_addr\[7\]
rlabel metal3 109940 186845 109940 186845 0 mprj/c0_o_mem_addr\[0\]
rlabel metal2 155158 330259 155158 330259 0 mprj/c0_o_mem_addr\[10\]
rlabel metal2 154790 333149 154790 333149 0 mprj/c0_o_mem_addr\[11\]
rlabel metal2 155066 335835 155066 335835 0 mprj/c0_o_mem_addr\[12\]
rlabel metal2 155066 338487 155066 338487 0 mprj/c0_o_mem_addr\[13\]
rlabel metal2 121210 317458 121210 317458 0 mprj/c0_o_mem_addr\[14\]
rlabel metal2 119370 322150 119370 322150 0 mprj/c0_o_mem_addr\[15\]
rlabel metal2 138782 249186 138782 249186 0 mprj/c0_o_mem_addr\[1\]
rlabel metal2 154790 305507 154790 305507 0 mprj/c0_o_mem_addr\[2\]
rlabel via2 154974 309179 154974 309179 0 mprj/c0_o_mem_addr\[3\]
rlabel metal2 154606 312273 154606 312273 0 mprj/c0_o_mem_addr\[4\]
rlabel metal2 154882 315265 154882 315265 0 mprj/c0_o_mem_addr\[5\]
rlabel metal2 136114 271490 136114 271490 0 mprj/c0_o_mem_addr\[6\]
rlabel metal2 154882 322031 154882 322031 0 mprj/c0_o_mem_addr\[7\]
rlabel metal2 121026 289068 121026 289068 0 mprj/c0_o_mem_addr\[8\]
rlabel metal3 156408 327964 156408 327964 0 mprj/c0_o_mem_addr\[9\]
rlabel metal3 109940 187389 109940 187389 0 mprj/c0_o_mem_addr_high\[0\]
rlabel metal2 154882 302617 154882 302617 0 mprj/c0_o_mem_addr_high\[1\]
rlabel via2 154974 306459 154974 306459 0 mprj/c0_o_mem_addr_high\[2\]
rlabel metal2 154606 309485 154606 309485 0 mprj/c0_o_mem_addr_high\[3\]
rlabel metal2 154882 312477 154882 312477 0 mprj/c0_o_mem_addr_high\[4\]
rlabel metal2 154974 316183 154974 316183 0 mprj/c0_o_mem_addr_high\[5\]
rlabel metal2 114310 278664 114310 278664 0 mprj/c0_o_mem_addr_high\[6\]
rlabel metal2 155066 322269 155066 322269 0 mprj/c0_o_mem_addr_high\[7\]
rlabel metal3 109940 188205 109940 188205 0 mprj/c0_o_mem_data\[0\]
rlabel metal2 155066 330429 155066 330429 0 mprj/c0_o_mem_data\[10\]
rlabel metal2 154974 333217 154974 333217 0 mprj/c0_o_mem_data\[11\]
rlabel metal2 154698 335903 154698 335903 0 mprj/c0_o_mem_data\[12\]
rlabel metal2 154882 338691 154882 338691 0 mprj/c0_o_mem_data\[13\]
rlabel metal2 154974 341479 154974 341479 0 mprj/c0_o_mem_data\[14\]
rlabel metal2 154974 344165 154974 344165 0 mprj/c0_o_mem_data\[15\]
rlabel metal3 155994 302668 155994 302668 0 mprj/c0_o_mem_data\[1\]
rlabel metal2 154882 305677 154882 305677 0 mprj/c0_o_mem_data\[2\]
rlabel metal2 154974 309383 154974 309383 0 mprj/c0_o_mem_data\[3\]
rlabel metal2 154790 312375 154790 312375 0 mprj/c0_o_mem_data\[4\]
rlabel metal2 155066 315435 155066 315435 0 mprj/c0_o_mem_data\[5\]
rlabel metal2 154974 319073 154974 319073 0 mprj/c0_o_mem_data\[6\]
rlabel metal2 115598 284274 115598 284274 0 mprj/c0_o_mem_data\[7\]
rlabel metal2 155066 325023 155066 325023 0 mprj/c0_o_mem_data\[8\]
rlabel metal2 155066 327675 155066 327675 0 mprj/c0_o_mem_data\[9\]
rlabel metal3 109940 178685 109940 178685 0 mprj/c0_o_mem_long
rlabel metal3 109940 179161 109940 179161 0 mprj/c0_o_mem_req
rlabel metal2 141542 244290 141542 244290 0 mprj/c0_o_mem_sel\[0\]
rlabel metal2 155158 302787 155158 302787 0 mprj/c0_o_mem_sel\[1\]
rlabel metal3 109940 180045 109940 180045 0 mprj/c0_o_mem_we
rlabel metal3 109940 180521 109940 180521 0 mprj/c0_o_req_active
rlabel metal3 109940 189565 109940 189565 0 mprj/c0_o_req_addr\[0\]
rlabel metal2 154974 331279 154974 331279 0 mprj/c0_o_req_addr\[10\]
rlabel metal2 154882 333319 154882 333319 0 mprj/c0_o_req_addr\[11\]
rlabel metal2 119830 308516 119830 308516 0 mprj/c0_o_req_addr\[12\]
rlabel metal2 154698 338793 154698 338793 0 mprj/c0_o_req_addr\[13\]
rlabel metal2 154790 341581 154790 341581 0 mprj/c0_o_req_addr\[14\]
rlabel metal2 120750 322898 120750 322898 0 mprj/c0_o_req_addr\[15\]
rlabel metal2 114034 250580 114034 250580 0 mprj/c0_o_req_addr\[1\]
rlabel metal2 154882 306629 154882 306629 0 mprj/c0_o_req_addr\[2\]
rlabel metal2 154790 309689 154790 309689 0 mprj/c0_o_req_addr\[3\]
rlabel metal2 154974 313361 154974 313361 0 mprj/c0_o_req_addr\[4\]
rlabel metal2 155066 316353 155066 316353 0 mprj/c0_o_req_addr\[5\]
rlabel metal2 154790 319379 154790 319379 0 mprj/c0_o_req_addr\[6\]
rlabel via2 154974 323085 154974 323085 0 mprj/c0_o_req_addr\[7\]
rlabel via2 154606 325805 154606 325805 0 mprj/c0_o_req_addr\[8\]
rlabel via2 154606 328525 154606 328525 0 mprj/c0_o_req_addr\[9\]
rlabel metal2 113850 238578 113850 238578 0 mprj/c0_o_req_ppl_submit
rlabel metal3 109940 175149 109940 175149 0 mprj/c0_rst
rlabel metal3 109940 190109 109940 190109 0 mprj/c0_sr_bus_addr\[0\]
rlabel metal2 154882 331449 154882 331449 0 mprj/c0_sr_bus_addr\[10\]
rlabel metal2 154974 334169 154974 334169 0 mprj/c0_sr_bus_addr\[11\]
rlabel metal2 133630 309842 133630 309842 0 mprj/c0_sr_bus_addr\[12\]
rlabel metal2 134734 314636 134734 314636 0 mprj/c0_sr_bus_addr\[13\]
rlabel metal2 139242 319464 139242 319464 0 mprj/c0_sr_bus_addr\[14\]
rlabel via2 154974 345083 154974 345083 0 mprj/c0_sr_bus_addr\[15\]
rlabel metal2 141634 251498 141634 251498 0 mprj/c0_sr_bus_addr\[1\]
rlabel metal2 154974 306799 154974 306799 0 mprj/c0_sr_bus_addr\[2\]
rlabel metal2 154882 309859 154882 309859 0 mprj/c0_sr_bus_addr\[3\]
rlabel via2 154974 313565 154974 313565 0 mprj/c0_sr_bus_addr\[4\]
rlabel metal1 153732 316370 153732 316370 0 mprj/c0_sr_bus_addr\[5\]
rlabel metal2 154882 319549 154882 319549 0 mprj/c0_sr_bus_addr\[6\]
rlabel metal2 114402 285668 114402 285668 0 mprj/c0_sr_bus_addr\[7\]
rlabel metal2 155066 325873 155066 325873 0 mprj/c0_sr_bus_addr\[8\]
rlabel metal2 154974 328729 154974 328729 0 mprj/c0_sr_bus_addr\[9\]
rlabel metal2 113942 245344 113942 245344 0 mprj/c0_sr_bus_data_o\[0\]
rlabel metal2 155066 331517 155066 331517 0 mprj/c0_sr_bus_data_o\[10\]
rlabel metal1 154100 333982 154100 333982 0 mprj/c0_sr_bus_data_o\[11\]
rlabel metal2 154606 337127 154606 337127 0 mprj/c0_sr_bus_data_o\[12\]
rlabel metal2 141818 314738 141818 314738 0 mprj/c0_sr_bus_data_o\[13\]
rlabel metal1 155480 335342 155480 335342 0 mprj/c0_sr_bus_data_o\[14\]
rlabel metal1 155112 306374 155112 306374 0 mprj/c0_sr_bus_data_o\[15\]
rlabel metal2 140346 251906 140346 251906 0 mprj/c0_sr_bus_data_o\[1\]
rlabel metal2 154790 306833 154790 306833 0 mprj/c0_sr_bus_data_o\[2\]
rlabel metal2 154882 310607 154882 310607 0 mprj/c0_sr_bus_data_o\[3\]
rlabel metal2 154606 313667 154606 313667 0 mprj/c0_sr_bus_data_o\[4\]
rlabel metal2 115506 274618 115506 274618 0 mprj/c0_sr_bus_data_o\[5\]
rlabel metal2 133354 280840 133354 280840 0 mprj/c0_sr_bus_data_o\[6\]
rlabel metal2 154974 323425 154974 323425 0 mprj/c0_sr_bus_data_o\[7\]
rlabel metal2 154790 326043 154790 326043 0 mprj/c0_sr_bus_data_o\[8\]
rlabel metal2 155066 328763 155066 328763 0 mprj/c0_sr_bus_data_o\[9\]
rlabel metal3 109940 181949 109940 181949 0 mprj/c0_sr_bus_we
rlabel metal2 154974 350217 154974 350217 0 mprj/c1_clk
rlabel metal3 156730 354892 156730 354892 0 mprj/c1_dbg_pc\[0\]
rlabel metal2 155066 387243 155066 387243 0 mprj/c1_dbg_pc\[10\]
rlabel metal2 154882 389997 154882 389997 0 mprj/c1_dbg_pc\[11\]
rlabel metal2 154882 392751 154882 392751 0 mprj/c1_dbg_pc\[12\]
rlabel metal2 154790 395573 154790 395573 0 mprj/c1_dbg_pc\[13\]
rlabel metal2 155066 398225 155066 398225 0 mprj/c1_dbg_pc\[14\]
rlabel metal1 153962 401574 153962 401574 0 mprj/c1_dbg_pc\[15\]
rlabel metal2 155112 364320 155112 364320 0 mprj/c1_dbg_pc\[1\]
rlabel metal2 114494 420240 114494 420240 0 mprj/c1_dbg_pc\[2\]
rlabel metal2 154974 365449 154974 365449 0 mprj/c1_dbg_pc\[3\]
rlabel metal2 154790 369019 154790 369019 0 mprj/c1_dbg_pc\[4\]
rlabel metal2 155158 372079 155158 372079 0 mprj/c1_dbg_pc\[5\]
rlabel metal2 141726 442918 141726 442918 0 mprj/c1_dbg_pc\[6\]
rlabel metal2 155066 378777 155066 378777 0 mprj/c1_dbg_pc\[7\]
rlabel metal2 139058 453968 139058 453968 0 mprj/c1_dbg_pc\[8\]
rlabel metal2 155158 384625 155158 384625 0 mprj/c1_dbg_pc\[9\]
rlabel metal2 137770 408476 137770 408476 0 mprj/c1_dbg_r0\[0\]
rlabel metal2 154882 387413 154882 387413 0 mprj/c1_dbg_r0\[10\]
rlabel metal2 154974 390099 154974 390099 0 mprj/c1_dbg_r0\[11\]
rlabel metal2 154974 392853 154974 392853 0 mprj/c1_dbg_r0\[12\]
rlabel metal2 154882 395675 154882 395675 0 mprj/c1_dbg_r0\[13\]
rlabel metal2 154882 398395 154882 398395 0 mprj/c1_dbg_r0\[14\]
rlabel metal2 154974 401115 154974 401115 0 mprj/c1_dbg_r0\[15\]
rlabel metal2 115138 413950 115138 413950 0 mprj/c1_dbg_r0\[1\]
rlabel metal2 154882 362491 154882 362491 0 mprj/c1_dbg_r0\[2\]
rlabel via2 154698 365483 154698 365483 0 mprj/c1_dbg_r0\[3\]
rlabel metal2 154698 369291 154698 369291 0 mprj/c1_dbg_r0\[4\]
rlabel metal2 154974 372181 154974 372181 0 mprj/c1_dbg_r0\[5\]
rlabel metal2 117162 442986 117162 442986 0 mprj/c1_dbg_r0\[6\]
rlabel metal3 156086 378556 156086 378556 0 mprj/c1_dbg_r0\[7\]
rlabel metal2 154606 381973 154606 381973 0 mprj/c1_dbg_r0\[8\]
rlabel metal2 155066 384727 155066 384727 0 mprj/c1_dbg_r0\[9\]
rlabel metal2 154606 350387 154606 350387 0 mprj/c1_disable
rlabel metal2 154882 355657 154882 355657 0 mprj/c1_i_core_int_sreg\[0\]
rlabel metal2 154974 387617 154974 387617 0 mprj/c1_i_core_int_sreg\[10\]
rlabel metal3 156684 390252 156684 390252 0 mprj/c1_i_core_int_sreg\[11\]
rlabel metal2 155066 393125 155066 393125 0 mprj/c1_i_core_int_sreg\[12\]
rlabel via2 154698 395709 154698 395709 0 mprj/c1_i_core_int_sreg\[13\]
rlabel metal1 153686 398786 153686 398786 0 mprj/c1_i_core_int_sreg\[14\]
rlabel metal2 141542 488512 141542 488512 0 mprj/c1_i_core_int_sreg\[15\]
rlabel metal2 154974 359431 154974 359431 0 mprj/c1_i_core_int_sreg\[1\]
rlabel metal2 118542 423368 118542 423368 0 mprj/c1_i_core_int_sreg\[2\]
rlabel metal3 156868 365772 156868 365772 0 mprj/c1_i_core_int_sreg\[3\]
rlabel metal2 155158 369393 155158 369393 0 mprj/c1_i_core_int_sreg\[4\]
rlabel metal2 154790 372419 154790 372419 0 mprj/c1_i_core_int_sreg\[5\]
rlabel metal2 139150 445400 139150 445400 0 mprj/c1_i_core_int_sreg\[6\]
rlabel metal2 118358 449412 118358 449412 0 mprj/c1_i_core_int_sreg\[7\]
rlabel metal2 154974 382143 154974 382143 0 mprj/c1_i_core_int_sreg\[8\]
rlabel via2 154974 384829 154974 384829 0 mprj/c1_i_core_int_sreg\[9\]
rlabel metal2 155066 351135 155066 351135 0 mprj/c1_i_irq
rlabel metal3 156638 350812 156638 350812 0 mprj/c1_i_mc_core_int
rlabel metal2 154882 351475 154882 351475 0 mprj/c1_i_mem_ack
rlabel metal2 119922 409122 119922 409122 0 mprj/c1_i_mem_data\[0\]
rlabel metal2 155250 388807 155250 388807 0 mprj/c1_i_mem_data\[10\]
rlabel metal2 154974 390439 154974 390439 0 mprj/c1_i_mem_data\[11\]
rlabel via2 154974 393227 154974 393227 0 mprj/c1_i_mem_data\[12\]
rlabel metal2 140162 479468 140162 479468 0 mprj/c1_i_mem_data\[13\]
rlabel metal2 137310 483582 137310 483582 0 mprj/c1_i_mem_data\[14\]
rlabel metal1 155204 405586 155204 405586 0 mprj/c1_i_mem_data\[15\]
rlabel metal2 142002 415310 142002 415310 0 mprj/c1_i_mem_data\[1\]
rlabel metal2 154974 362729 154974 362729 0 mprj/c1_i_mem_data\[2\]
rlabel metal2 154882 366435 154882 366435 0 mprj/c1_i_mem_data\[3\]
rlabel metal2 154882 369461 154882 369461 0 mprj/c1_i_mem_data\[4\]
rlabel metal2 154974 372521 154974 372521 0 mprj/c1_i_mem_data\[5\]
rlabel metal2 121026 443258 121026 443258 0 mprj/c1_i_mem_data\[6\]
rlabel metal2 120842 449888 120842 449888 0 mprj/c1_i_mem_data\[7\]
rlabel metal2 154698 382891 154698 382891 0 mprj/c1_i_mem_data\[8\]
rlabel metal2 155066 385713 155066 385713 0 mprj/c1_i_mem_data\[9\]
rlabel metal2 154790 351509 154790 351509 0 mprj/c1_i_mem_exception
rlabel metal1 153824 356014 153824 356014 0 mprj/c1_i_req_data\[0\]
rlabel metal2 154882 388603 154882 388603 0 mprj/c1_i_req_data\[10\]
rlabel metal3 155994 390796 155994 390796 0 mprj/c1_i_req_data\[11\]
rlabel metal2 154882 393975 154882 393975 0 mprj/c1_i_req_data\[12\]
rlabel metal2 122682 452948 122682 452948 0 mprj/c1_i_req_data\[13\]
rlabel metal2 122314 485452 122314 485452 0 mprj/c1_i_req_data\[14\]
rlabel metal2 122406 483174 122406 483174 0 mprj/c1_i_req_data\[15\]
rlabel metal2 154882 403733 154882 403733 0 mprj/c1_i_req_data\[16\]
rlabel metal2 154974 403903 154974 403903 0 mprj/c1_i_req_data\[17\]
rlabel metal2 154790 403971 154790 403971 0 mprj/c1_i_req_data\[18\]
rlabel metal2 154698 404209 154698 404209 0 mprj/c1_i_req_data\[19\]
rlabel metal2 122590 416126 122590 416126 0 mprj/c1_i_req_data\[1\]
rlabel metal2 155802 406079 155802 406079 0 mprj/c1_i_req_data\[20\]
rlabel metal2 154882 405127 154882 405127 0 mprj/c1_i_req_data\[21\]
rlabel metal2 154974 405229 154974 405229 0 mprj/c1_i_req_data\[22\]
rlabel metal2 154790 405433 154790 405433 0 mprj/c1_i_req_data\[23\]
rlabel via2 154606 405467 154606 405467 0 mprj/c1_i_req_data\[24\]
rlabel metal2 154698 407439 154698 407439 0 mprj/c1_i_req_data\[25\]
rlabel metal2 154790 406521 154790 406521 0 mprj/c1_i_req_data\[26\]
rlabel metal2 154882 406691 154882 406691 0 mprj/c1_i_req_data\[27\]
rlabel metal2 154974 406759 154974 406759 0 mprj/c1_i_req_data\[28\]
rlabel via2 154606 406861 154606 406861 0 mprj/c1_i_req_data\[29\]
rlabel metal3 156684 363052 156684 363052 0 mprj/c1_i_req_data\[2\]
rlabel metal3 156914 407116 156914 407116 0 mprj/c1_i_req_data\[30\]
rlabel metal2 154974 407915 154974 407915 0 mprj/c1_i_req_data\[31\]
rlabel metal2 154698 366605 154698 366605 0 mprj/c1_i_req_data\[3\]
rlabel metal2 154974 369631 154974 369631 0 mprj/c1_i_req_data\[4\]
rlabel metal2 154698 373405 154698 373405 0 mprj/c1_i_req_data\[5\]
rlabel metal2 154882 376329 154882 376329 0 mprj/c1_i_req_data\[6\]
rlabel via2 154974 379355 154974 379355 0 mprj/c1_i_req_data\[7\]
rlabel metal2 154974 382993 154974 382993 0 mprj/c1_i_req_data\[8\]
rlabel metal2 154882 385781 154882 385781 0 mprj/c1_i_req_data\[9\]
rlabel metal2 154974 351713 154974 351713 0 mprj/c1_i_req_data_valid
rlabel metal3 156776 351900 156776 351900 0 mprj/c1_o_c_data_page
rlabel metal2 154882 352563 154882 352563 0 mprj/c1_o_c_instr_long
rlabel metal2 154790 352835 154790 352835 0 mprj/c1_o_c_instr_page
rlabel metal2 155066 352869 155066 352869 0 mprj/c1_o_icache_flush
rlabel metal2 154790 356779 154790 356779 0 mprj/c1_o_instr_long_addr\[0\]
rlabel metal2 155066 359941 155066 359941 0 mprj/c1_o_instr_long_addr\[1\]
rlabel metal2 155066 363783 155066 363783 0 mprj/c1_o_instr_long_addr\[2\]
rlabel metal2 155158 366809 155158 366809 0 mprj/c1_o_instr_long_addr\[3\]
rlabel metal3 156730 369852 156730 369852 0 mprj/c1_o_instr_long_addr\[4\]
rlabel metal2 154790 373507 154790 373507 0 mprj/c1_o_instr_long_addr\[5\]
rlabel metal2 154974 376431 154974 376431 0 mprj/c1_o_instr_long_addr\[6\]
rlabel metal2 155066 380171 155066 380171 0 mprj/c1_o_instr_long_addr\[7\]
rlabel metal2 154882 356847 154882 356847 0 mprj/c1_o_mem_addr\[0\]
rlabel metal2 154974 388637 154974 388637 0 mprj/c1_o_mem_addr\[10\]
rlabel metal2 154974 391357 154974 391357 0 mprj/c1_o_mem_addr\[11\]
rlabel metal2 154974 394553 154974 394553 0 mprj/c1_o_mem_addr\[12\]
rlabel metal2 154790 397307 154790 397307 0 mprj/c1_o_mem_addr\[13\]
rlabel metal2 154790 399687 154790 399687 0 mprj/c1_o_mem_addr\[14\]
rlabel metal1 153916 402458 153916 402458 0 mprj/c1_o_mem_addr\[15\]
rlabel via2 154974 360043 154974 360043 0 mprj/c1_o_mem_addr\[1\]
rlabel metal2 154882 363885 154882 363885 0 mprj/c1_o_mem_addr\[2\]
rlabel metal2 154974 366911 154974 366911 0 mprj/c1_o_mem_addr\[3\]
rlabel metal2 154698 370617 154698 370617 0 mprj/c1_o_mem_addr\[4\]
rlabel metal2 154882 373541 154882 373541 0 mprj/c1_o_mem_addr\[5\]
rlabel metal2 114218 445774 114218 445774 0 mprj/c1_o_mem_addr\[6\]
rlabel metal2 118266 451248 118266 451248 0 mprj/c1_o_mem_addr\[7\]
rlabel metal3 156040 382908 156040 382908 0 mprj/c1_o_mem_addr\[8\]
rlabel metal2 155250 389980 155250 389980 0 mprj/c1_o_mem_addr\[9\]
rlabel metal2 155066 357221 155066 357221 0 mprj/c1_o_mem_addr_high\[0\]
rlabel metal2 154790 361029 154790 361029 0 mprj/c1_o_mem_addr_high\[1\]
rlabel via2 154974 364123 154974 364123 0 mprj/c1_o_mem_addr_high\[2\]
rlabel metal2 154790 367897 154790 367897 0 mprj/c1_o_mem_addr_high\[3\]
rlabel metal2 154882 370821 154882 370821 0 mprj/c1_o_mem_addr_high\[4\]
rlabel metal2 154606 373881 154606 373881 0 mprj/c1_o_mem_addr_high\[5\]
rlabel metal2 120934 446386 120934 446386 0 mprj/c1_o_mem_addr_high\[6\]
rlabel metal2 154974 380511 154974 380511 0 mprj/c1_o_mem_addr_high\[7\]
rlabel metal2 154974 356949 154974 356949 0 mprj/c1_o_mem_data\[0\]
rlabel metal2 113206 520999 113206 520999 0 mprj/c1_o_mem_data\[10\]
rlabel metal2 154790 391561 154790 391561 0 mprj/c1_o_mem_data\[11\]
rlabel metal2 154790 394281 154790 394281 0 mprj/c1_o_mem_data\[12\]
rlabel metal2 154882 397035 154882 397035 0 mprj/c1_o_mem_data\[13\]
rlabel metal2 155066 399789 155066 399789 0 mprj/c1_o_mem_data\[14\]
rlabel metal2 154790 402543 154790 402543 0 mprj/c1_o_mem_data\[15\]
rlabel metal2 115874 417792 115874 417792 0 mprj/c1_o_mem_data\[1\]
rlabel metal2 154790 364089 154790 364089 0 mprj/c1_o_mem_data\[2\]
rlabel metal2 154882 367693 154882 367693 0 mprj/c1_o_mem_data\[3\]
rlabel metal2 154790 370787 154790 370787 0 mprj/c1_o_mem_data\[4\]
rlabel metal2 154974 373711 154974 373711 0 mprj/c1_o_mem_data\[5\]
rlabel metal2 140346 447032 140346 447032 0 mprj/c1_o_mem_data\[6\]
rlabel metal2 154882 380409 154882 380409 0 mprj/c1_o_mem_data\[7\]
rlabel metal2 154882 383367 154882 383367 0 mprj/c1_o_mem_data\[8\]
rlabel metal2 154698 386087 154698 386087 0 mprj/c1_o_mem_data\[9\]
rlabel metal2 154974 353073 154974 353073 0 mprj/c1_o_mem_long
rlabel metal2 154882 353175 154882 353175 0 mprj/c1_o_mem_req
rlabel metal2 154974 357289 154974 357289 0 mprj/c1_o_mem_sel\[0\]
rlabel metal2 154882 361131 154882 361131 0 mprj/c1_o_mem_sel\[1\]
rlabel metal2 154882 354093 154882 354093 0 mprj/c1_o_mem_we
rlabel metal3 156868 353804 156868 353804 0 mprj/c1_o_req_active
rlabel metal2 137678 412522 137678 412522 0 mprj/c1_o_req_addr\[0\]
rlabel metal2 154698 388943 154698 388943 0 mprj/c1_o_req_addr\[10\]
rlabel metal2 154698 391663 154698 391663 0 mprj/c1_o_req_addr\[11\]
rlabel metal2 154606 394485 154606 394485 0 mprj/c1_o_req_addr\[12\]
rlabel metal2 155066 397239 155066 397239 0 mprj/c1_o_req_addr\[13\]
rlabel metal2 133262 485690 133262 485690 0 mprj/c1_o_req_addr\[14\]
rlabel metal2 133170 490518 133170 490518 0 mprj/c1_o_req_addr\[15\]
rlabel metal2 133538 418030 133538 418030 0 mprj/c1_o_req_addr\[1\]
rlabel metal2 155158 365007 155158 365007 0 mprj/c1_o_req_addr\[2\]
rlabel metal3 156822 367676 156822 367676 0 mprj/c1_o_req_addr\[3\]
rlabel metal2 154974 370991 154974 370991 0 mprj/c1_o_req_addr\[4\]
rlabel metal3 156776 374204 156776 374204 0 mprj/c1_o_req_addr\[5\]
rlabel metal2 119738 447134 119738 447134 0 mprj/c1_o_req_addr\[6\]
rlabel metal2 154974 380783 154974 380783 0 mprj/c1_o_req_addr\[7\]
rlabel metal2 138966 457436 138966 457436 0 mprj/c1_o_req_addr\[8\]
rlabel via2 154974 386155 154974 386155 0 mprj/c1_o_req_addr\[9\]
rlabel metal2 154790 354263 154790 354263 0 mprj/c1_o_req_ppl_submit
rlabel metal2 154974 354433 154974 354433 0 mprj/c1_rst
rlabel metal2 117254 413304 117254 413304 0 mprj/c1_sr_bus_addr\[0\]
rlabel metal2 155066 389793 155066 389793 0 mprj/c1_sr_bus_addr\[10\]
rlabel via2 154974 391867 154974 391867 0 mprj/c1_sr_bus_addr\[11\]
rlabel via2 154698 394587 154698 394587 0 mprj/c1_sr_bus_addr\[12\]
rlabel metal2 134734 481542 134734 481542 0 mprj/c1_sr_bus_addr\[13\]
rlabel metal2 134642 486370 134642 486370 0 mprj/c1_sr_bus_addr\[14\]
rlabel metal2 134550 491198 134550 491198 0 mprj/c1_sr_bus_addr\[15\]
rlabel metal2 136114 418676 136114 418676 0 mprj/c1_sr_bus_addr\[1\]
rlabel metal2 154882 365109 154882 365109 0 mprj/c1_sr_bus_addr\[2\]
rlabel metal2 154974 368135 154974 368135 0 mprj/c1_sr_bus_addr\[3\]
rlabel metal2 155158 371059 155158 371059 0 mprj/c1_sr_bus_addr\[4\]
rlabel metal2 155158 375241 155158 375241 0 mprj/c1_sr_bus_addr\[5\]
rlabel metal2 154974 377791 154974 377791 0 mprj/c1_sr_bus_addr\[6\]
rlabel metal3 156822 381004 156822 381004 0 mprj/c1_sr_bus_addr\[7\]
rlabel metal2 154698 384217 154698 384217 0 mprj/c1_sr_bus_addr\[8\]
rlabel metal2 155158 387107 155158 387107 0 mprj/c1_sr_bus_addr\[9\]
rlabel metal1 154284 358734 154284 358734 0 mprj/c1_sr_bus_data_o\[0\]
rlabel metal1 153732 390490 153732 390490 0 mprj/c1_sr_bus_data_o\[10\]
rlabel metal2 154790 392649 154790 392649 0 mprj/c1_sr_bus_data_o\[11\]
rlabel metal2 140254 478040 140254 478040 0 mprj/c1_sr_bus_data_o\[12\]
rlabel metal2 141634 482970 141634 482970 0 mprj/c1_sr_bus_data_o\[13\]
rlabel metal2 155066 400877 155066 400877 0 mprj/c1_sr_bus_data_o\[14\]
rlabel metal3 156684 403036 156684 403036 0 mprj/c1_sr_bus_data_o\[15\]
rlabel metal2 154606 362287 154606 362287 0 mprj/c1_sr_bus_data_o\[1\]
rlabel metal2 154790 365177 154790 365177 0 mprj/c1_sr_bus_data_o\[2\]
rlabel metal2 154606 368339 154606 368339 0 mprj/c1_sr_bus_data_o\[3\]
rlabel metal2 154882 371875 154882 371875 0 mprj/c1_sr_bus_data_o\[4\]
rlabel metal1 154054 375360 154054 375360 0 mprj/c1_sr_bus_data_o\[5\]
rlabel metal2 154974 378063 154974 378063 0 mprj/c1_sr_bus_data_o\[6\]
rlabel metal2 154974 381633 154974 381633 0 mprj/c1_sr_bus_data_o\[7\]
rlabel metal2 154882 384387 154882 384387 0 mprj/c1_sr_bus_data_o\[8\]
rlabel metal2 154790 387175 154790 387175 0 mprj/c1_sr_bus_data_o\[9\]
rlabel via2 154606 354603 154606 354603 0 mprj/c1_sr_bus_we
rlabel metal1 256358 51034 256358 51034 0 mprj/dcache_clk
rlabel metal2 232806 259828 232806 259828 0 mprj/dcache_mem_ack
rlabel metal2 256726 76585 256726 76585 0 mprj/dcache_mem_addr\[0\]
rlabel metal1 255806 206958 255806 206958 0 mprj/dcache_mem_addr\[10\]
rlabel metal2 256726 219079 256726 219079 0 mprj/dcache_mem_addr\[11\]
rlabel metal2 256358 276301 256358 276301 0 mprj/dcache_mem_addr\[12\]
rlabel metal2 235566 284308 235566 284308 0 mprj/dcache_mem_addr\[13\]
rlabel metal2 256726 256071 256726 256071 0 mprj/dcache_mem_addr\[14\]
rlabel metal1 256910 289782 256910 289782 0 mprj/dcache_mem_addr\[15\]
rlabel metal1 255852 280126 255852 280126 0 mprj/dcache_mem_addr\[16\]
rlabel metal2 257646 294831 257646 294831 0 mprj/dcache_mem_addr\[17\]
rlabel metal2 256726 288235 256726 288235 0 mprj/dcache_mem_addr\[18\]
rlabel metal1 253184 292502 253184 292502 0 mprj/dcache_mem_addr\[19\]
rlabel metal1 255714 92446 255714 92446 0 mprj/dcache_mem_addr\[1\]
rlabel metal2 256726 296463 256726 296463 0 mprj/dcache_mem_addr\[20\]
rlabel metal2 256726 300577 256726 300577 0 mprj/dcache_mem_addr\[21\]
rlabel metal2 257738 308499 257738 308499 0 mprj/dcache_mem_addr\[22\]
rlabel metal2 256726 308805 256726 308805 0 mprj/dcache_mem_addr\[23\]
rlabel metal2 256726 108783 256726 108783 0 mprj/dcache_mem_addr\[2\]
rlabel metal2 256726 121125 256726 121125 0 mprj/dcache_mem_addr\[3\]
rlabel metal2 256726 133467 256726 133467 0 mprj/dcache_mem_addr\[4\]
rlabel metal2 256726 145775 256726 145775 0 mprj/dcache_mem_addr\[5\]
rlabel metal2 232898 286756 232898 286756 0 mprj/dcache_mem_addr\[6\]
rlabel metal2 234278 240142 234278 240142 0 mprj/dcache_mem_addr\[7\]
rlabel metal2 235474 247010 235474 247010 0 mprj/dcache_mem_addr\[8\]
rlabel metal2 256726 194395 256726 194395 0 mprj/dcache_mem_addr\[9\]
rlabel metal2 256726 56049 256726 56049 0 mprj/dcache_mem_cache_enable
rlabel metal2 256726 57749 256726 57749 0 mprj/dcache_mem_exception
rlabel metal1 253644 78642 253644 78642 0 mprj/dcache_mem_i_data\[0\]
rlabel metal2 256266 263007 256266 263007 0 mprj/dcache_mem_i_data\[10\]
rlabel via2 256726 220779 256726 220779 0 mprj/dcache_mem_i_data\[11\]
rlabel metal2 256726 233121 256726 233121 0 mprj/dcache_mem_i_data\[12\]
rlabel metal2 256726 245429 256726 245429 0 mprj/dcache_mem_i_data\[13\]
rlabel metal2 256726 257771 256726 257771 0 mprj/dcache_mem_i_data\[14\]
rlabel metal2 256726 270113 256726 270113 0 mprj/dcache_mem_i_data\[15\]
rlabel metal2 256726 94741 256726 94741 0 mprj/dcache_mem_i_data\[1\]
rlabel metal2 256726 111197 256726 111197 0 mprj/dcache_mem_i_data\[2\]
rlabel metal3 217948 300409 217948 300409 0 mprj/dcache_mem_i_data\[3\]
rlabel metal2 256726 135167 256726 135167 0 mprj/dcache_mem_i_data\[4\]
rlabel metal2 256726 147475 256726 147475 0 mprj/dcache_mem_i_data\[5\]
rlabel metal2 256726 159817 256726 159817 0 mprj/dcache_mem_i_data\[6\]
rlabel metal2 256726 172159 256726 172159 0 mprj/dcache_mem_i_data\[7\]
rlabel metal2 256726 184467 256726 184467 0 mprj/dcache_mem_i_data\[8\]
rlabel metal2 256726 196809 256726 196809 0 mprj/dcache_mem_i_data\[9\]
rlabel metal1 252954 80002 252954 80002 0 mprj/dcache_mem_o_data\[0\]
rlabel metal2 256726 210851 256726 210851 0 mprj/dcache_mem_o_data\[10\]
rlabel metal2 256726 223193 256726 223193 0 mprj/dcache_mem_o_data\[11\]
rlabel metal2 257370 259335 257370 259335 0 mprj/dcache_mem_o_data\[12\]
rlabel metal2 256726 247843 256726 247843 0 mprj/dcache_mem_o_data\[13\]
rlabel metal2 256726 260185 256726 260185 0 mprj/dcache_mem_o_data\[14\]
rlabel metal1 253966 292774 253966 292774 0 mprj/dcache_mem_o_data\[15\]
rlabel metal2 256726 96475 256726 96475 0 mprj/dcache_mem_o_data\[1\]
rlabel metal1 255760 112914 255760 112914 0 mprj/dcache_mem_o_data\[2\]
rlabel metal2 234002 213282 234002 213282 0 mprj/dcache_mem_o_data\[3\]
rlabel metal2 257554 147577 257554 147577 0 mprj/dcache_mem_o_data\[4\]
rlabel metal2 256726 149889 256726 149889 0 mprj/dcache_mem_o_data\[5\]
rlabel metal2 238234 235348 238234 235348 0 mprj/dcache_mem_o_data\[6\]
rlabel metal2 257830 205955 257830 205955 0 mprj/dcache_mem_o_data\[7\]
rlabel metal2 256726 186201 256726 186201 0 mprj/dcache_mem_o_data\[8\]
rlabel metal2 256726 198509 256726 198509 0 mprj/dcache_mem_o_data\[9\]
rlabel metal2 256726 60163 256726 60163 0 mprj/dcache_mem_req
rlabel metal2 256726 82433 256726 82433 0 mprj/dcache_mem_sel\[0\]
rlabel metal2 256082 196877 256082 196877 0 mprj/dcache_mem_sel\[1\]
rlabel metal2 256726 61863 256726 61863 0 mprj/dcache_mem_we
rlabel metal2 256726 52989 256726 52989 0 mprj/dcache_rst
rlabel metal1 253598 64430 253598 64430 0 mprj/dcache_wb_4_burst
rlabel metal2 236762 214268 236762 214268 0 mprj/dcache_wb_ack
rlabel via2 256726 84133 256726 84133 0 mprj/dcache_wb_adr\[0\]
rlabel metal2 256726 213265 256726 213265 0 mprj/dcache_wb_adr\[10\]
rlabel metal1 253138 224910 253138 224910 0 mprj/dcache_wb_adr\[11\]
rlabel metal2 256726 237235 256726 237235 0 mprj/dcache_wb_adr\[12\]
rlabel metal2 256726 249543 256726 249543 0 mprj/dcache_wb_adr\[13\]
rlabel metal2 256726 261885 256726 261885 0 mprj/dcache_wb_adr\[14\]
rlabel metal2 256726 274227 256726 274227 0 mprj/dcache_wb_adr\[15\]
rlabel metal2 256726 282421 256726 282421 0 mprj/dcache_wb_adr\[16\]
rlabel metal2 257370 306901 257370 306901 0 mprj/dcache_wb_adr\[17\]
rlabel metal2 256726 290649 256726 290649 0 mprj/dcache_wb_adr\[18\]
rlabel metal2 256726 294763 256726 294763 0 mprj/dcache_wb_adr\[19\]
rlabel metal2 256726 100555 256726 100555 0 mprj/dcache_wb_adr\[1\]
rlabel metal2 256726 298877 256726 298877 0 mprj/dcache_wb_adr\[20\]
rlabel metal2 256726 302991 256726 302991 0 mprj/dcache_wb_adr\[21\]
rlabel metal2 256818 308125 256818 308125 0 mprj/dcache_wb_adr\[22\]
rlabel metal2 256726 311185 256726 311185 0 mprj/dcache_wb_adr\[23\]
rlabel metal2 256726 115311 256726 115311 0 mprj/dcache_wb_adr\[2\]
rlabel metal2 232622 213996 232622 213996 0 mprj/dcache_wb_adr\[3\]
rlabel metal2 256726 139281 256726 139281 0 mprj/dcache_wb_adr\[4\]
rlabel metal2 256726 151589 256726 151589 0 mprj/dcache_wb_adr\[5\]
rlabel metal2 256726 163931 256726 163931 0 mprj/dcache_wb_adr\[6\]
rlabel metal2 256726 176273 256726 176273 0 mprj/dcache_wb_adr\[7\]
rlabel metal2 230138 251226 230138 251226 0 mprj/dcache_wb_adr\[8\]
rlabel metal2 230230 258094 230230 258094 0 mprj/dcache_wb_adr\[9\]
rlabel metal2 229862 178772 229862 178772 0 mprj/dcache_wb_cyc
rlabel metal2 256726 70091 256726 70091 0 mprj/dcache_wb_err
rlabel metal2 256726 86547 256726 86547 0 mprj/dcache_wb_i_dat\[0\]
rlabel metal1 254380 215254 254380 215254 0 mprj/dcache_wb_i_dat\[10\]
rlabel metal2 256726 227307 256726 227307 0 mprj/dcache_wb_i_dat\[11\]
rlabel metal2 231518 281520 231518 281520 0 mprj/dcache_wb_i_dat\[12\]
rlabel metal2 256726 251957 256726 251957 0 mprj/dcache_wb_i_dat\[13\]
rlabel metal2 231610 296718 231610 296718 0 mprj/dcache_wb_i_dat\[14\]
rlabel metal2 256726 275927 256726 275927 0 mprj/dcache_wb_i_dat\[15\]
rlabel metal2 256726 102969 256726 102969 0 mprj/dcache_wb_i_dat\[1\]
rlabel metal2 256726 117011 256726 117011 0 mprj/dcache_wb_i_dat\[2\]
rlabel metal2 234186 215322 234186 215322 0 mprj/dcache_wb_i_dat\[3\]
rlabel metal2 256726 141661 256726 141661 0 mprj/dcache_wb_i_dat\[4\]
rlabel metal2 256726 154003 256726 154003 0 mprj/dcache_wb_i_dat\[5\]
rlabel metal2 256726 166345 256726 166345 0 mprj/dcache_wb_i_dat\[6\]
rlabel via2 256726 177973 256726 177973 0 mprj/dcache_wb_i_dat\[7\]
rlabel metal2 256726 190315 256726 190315 0 mprj/dcache_wb_i_dat\[8\]
rlabel metal2 256726 202623 256726 202623 0 mprj/dcache_wb_i_dat\[9\]
rlabel metal1 253046 88298 253046 88298 0 mprj/dcache_wb_o_dat\[0\]
rlabel metal2 256726 217345 256726 217345 0 mprj/dcache_wb_o_dat\[10\]
rlabel metal1 253736 228990 253736 228990 0 mprj/dcache_wb_o_dat\[11\]
rlabel metal2 256726 241315 256726 241315 0 mprj/dcache_wb_o_dat\[12\]
rlabel metal2 256726 253657 256726 253657 0 mprj/dcache_wb_o_dat\[13\]
rlabel metal2 256726 265999 256726 265999 0 mprj/dcache_wb_o_dat\[14\]
rlabel metal2 256726 278307 256726 278307 0 mprj/dcache_wb_o_dat\[15\]
rlabel metal2 256726 104669 256726 104669 0 mprj/dcache_wb_o_dat\[1\]
rlabel metal1 254334 120054 254334 120054 0 mprj/dcache_wb_o_dat\[2\]
rlabel metal2 256174 215951 256174 215951 0 mprj/dcache_wb_o_dat\[3\]
rlabel metal1 253690 143514 253690 143514 0 mprj/dcache_wb_o_dat\[4\]
rlabel metal2 256726 155703 256726 155703 0 mprj/dcache_wb_o_dat\[5\]
rlabel metal2 256726 168045 256726 168045 0 mprj/dcache_wb_o_dat\[6\]
rlabel metal2 256726 180387 256726 180387 0 mprj/dcache_wb_o_dat\[7\]
rlabel metal1 253092 193154 253092 193154 0 mprj/dcache_wb_o_dat\[8\]
rlabel metal2 256726 205037 256726 205037 0 mprj/dcache_wb_o_dat\[9\]
rlabel metal2 256726 90627 256726 90627 0 mprj/dcache_wb_sel\[0\]
rlabel metal2 256726 107083 256726 107083 0 mprj/dcache_wb_sel\[1\]
rlabel metal2 256726 72505 256726 72505 0 mprj/dcache_wb_stb
rlabel metal2 256726 74205 256726 74205 0 mprj/dcache_wb_we
rlabel metal2 234278 360774 234278 360774 0 mprj/ic0_clk
rlabel metal3 252548 386036 252548 386036 0 mprj/ic0_mem_ack
rlabel metal2 251206 396559 251206 396559 0 mprj/ic0_mem_addr\[0\]
rlabel metal3 253008 448460 253008 448460 0 mprj/ic0_mem_addr\[10\]
rlabel metal1 252034 446454 252034 446454 0 mprj/ic0_mem_addr\[11\]
rlabel metal3 252870 458252 252870 458252 0 mprj/ic0_mem_addr\[12\]
rlabel metal2 251206 462757 251206 462757 0 mprj/ic0_mem_addr\[13\]
rlabel metal3 252916 468044 252916 468044 0 mprj/ic0_mem_addr\[14\]
rlabel metal2 251206 472481 251206 472481 0 mprj/ic0_mem_addr\[15\]
rlabel metal3 252364 403172 252364 403172 0 mprj/ic0_mem_addr\[1\]
rlabel metal2 251206 408901 251206 408901 0 mprj/ic0_mem_addr\[2\]
rlabel metal2 251206 414103 251206 414103 0 mprj/ic0_mem_addr\[3\]
rlabel metal2 251206 418625 251206 418625 0 mprj/ic0_mem_addr\[4\]
rlabel metal1 250102 423674 250102 423674 0 mprj/ic0_mem_addr\[5\]
rlabel metal2 251206 428349 251206 428349 0 mprj/ic0_mem_addr\[6\]
rlabel metal2 238602 395692 238602 395692 0 mprj/ic0_mem_addr\[7\]
rlabel metal2 251206 438073 251206 438073 0 mprj/ic0_mem_addr\[8\]
rlabel metal3 252272 443564 252272 443564 0 mprj/ic0_mem_addr\[9\]
rlabel metal3 252686 387260 252686 387260 0 mprj/ic0_mem_cache_flush
rlabel metal2 251206 397885 251206 397885 0 mprj/ic0_mem_data\[0\]
rlabel metal2 251206 449123 251206 449123 0 mprj/ic0_mem_data\[10\]
rlabel metal2 251206 454325 251206 454325 0 mprj/ic0_mem_data\[11\]
rlabel metal2 251206 458847 251206 458847 0 mprj/ic0_mem_data\[12\]
rlabel metal2 251206 464049 251206 464049 0 mprj/ic0_mem_data\[13\]
rlabel via2 251206 469285 251206 469285 0 mprj/ic0_mem_data\[14\]
rlabel metal2 251206 473773 251206 473773 0 mprj/ic0_mem_data\[15\]
rlabel metal2 251206 477683 251206 477683 0 mprj/ic0_mem_data\[16\]
rlabel metal1 250424 478890 250424 478890 0 mprj/ic0_mem_data\[17\]
rlabel metal3 253008 480284 253008 480284 0 mprj/ic0_mem_data\[18\]
rlabel metal2 251206 480879 251206 480879 0 mprj/ic0_mem_data\[19\]
rlabel metal3 252686 404396 252686 404396 0 mprj/ic0_mem_data\[1\]
rlabel metal2 251206 482205 251206 482205 0 mprj/ic0_mem_data\[20\]
rlabel metal2 251206 483497 251206 483497 0 mprj/ic0_mem_data\[21\]
rlabel metal2 251206 484789 251206 484789 0 mprj/ic0_mem_data\[22\]
rlabel metal2 251206 486115 251206 486115 0 mprj/ic0_mem_data\[23\]
rlabel metal2 251206 487407 251206 487407 0 mprj/ic0_mem_data\[24\]
rlabel metal2 251206 488699 251206 488699 0 mprj/ic0_mem_data\[25\]
rlabel metal2 251206 489991 251206 489991 0 mprj/ic0_mem_data\[26\]
rlabel metal3 252226 491300 252226 491300 0 mprj/ic0_mem_data\[27\]
rlabel metal2 251206 491929 251206 491929 0 mprj/ic0_mem_data\[28\]
rlabel metal2 251206 493221 251206 493221 0 mprj/ic0_mem_data\[29\]
rlabel metal2 251206 410193 251206 410193 0 mprj/ic0_mem_data\[2\]
rlabel metal2 251206 494513 251206 494513 0 mprj/ic0_mem_data\[30\]
rlabel metal2 251206 495839 251206 495839 0 mprj/ic0_mem_data\[31\]
rlabel via2 251206 415429 251206 415429 0 mprj/ic0_mem_data\[3\]
rlabel metal2 251206 419917 251206 419917 0 mprj/ic0_mem_data\[4\]
rlabel metal2 251206 425153 251206 425153 0 mprj/ic0_mem_data\[5\]
rlabel metal2 251206 429641 251206 429641 0 mprj/ic0_mem_data\[6\]
rlabel metal2 251206 434877 251206 434877 0 mprj/ic0_mem_data\[7\]
rlabel metal2 251206 439399 251206 439399 0 mprj/ic0_mem_data\[8\]
rlabel metal2 251206 444601 251206 444601 0 mprj/ic0_mem_data\[9\]
rlabel metal1 250332 387838 250332 387838 0 mprj/ic0_mem_ppl_submit
rlabel metal2 251206 389453 251206 389453 0 mprj/ic0_mem_req
rlabel metal2 251206 384251 251206 384251 0 mprj/ic0_rst
rlabel metal2 251206 390745 251206 390745 0 mprj/ic0_wb_ack
rlabel metal2 251206 399177 251206 399177 0 mprj/ic0_wb_adr\[0\]
rlabel metal2 251206 450415 251206 450415 0 mprj/ic0_wb_adr\[10\]
rlabel metal2 251206 455617 251206 455617 0 mprj/ic0_wb_adr\[11\]
rlabel metal2 251206 460139 251206 460139 0 mprj/ic0_wb_adr\[12\]
rlabel metal1 250700 465086 250700 465086 0 mprj/ic0_wb_adr\[13\]
rlabel metal2 251298 469863 251298 469863 0 mprj/ic0_wb_adr\[14\]
rlabel metal2 251206 475065 251206 475065 0 mprj/ic0_wb_adr\[15\]
rlabel metal2 251206 404991 251206 404991 0 mprj/ic0_wb_adr\[1\]
rlabel metal2 251206 411519 251206 411519 0 mprj/ic0_wb_adr\[2\]
rlabel metal2 251298 416075 251298 416075 0 mprj/ic0_wb_adr\[3\]
rlabel metal2 251206 421243 251206 421243 0 mprj/ic0_wb_adr\[4\]
rlabel via2 251206 426445 251206 426445 0 mprj/ic0_wb_adr\[5\]
rlabel metal2 251206 430967 251206 430967 0 mprj/ic0_wb_adr\[6\]
rlabel via2 251206 436203 251206 436203 0 mprj/ic0_wb_adr\[7\]
rlabel metal2 251206 440691 251206 440691 0 mprj/ic0_wb_adr\[8\]
rlabel metal2 251206 445893 251206 445893 0 mprj/ic0_wb_adr\[9\]
rlabel metal2 251206 392071 251206 392071 0 mprj/ic0_wb_cyc
rlabel via2 251206 393363 251206 393363 0 mprj/ic0_wb_err
rlabel metal1 251206 393890 251206 393890 0 mprj/ic0_wb_i_dat\[0\]
rlabel metal2 251206 451707 251206 451707 0 mprj/ic0_wb_i_dat\[10\]
rlabel metal2 238510 409768 238510 409768 0 mprj/ic0_wb_i_dat\[11\]
rlabel metal1 252126 446318 252126 446318 0 mprj/ic0_wb_i_dat\[12\]
rlabel metal2 251206 466633 251206 466633 0 mprj/ic0_wb_i_dat\[13\]
rlabel metal2 230138 419526 230138 419526 0 mprj/ic0_wb_i_dat\[14\]
rlabel metal2 251206 476357 251206 476357 0 mprj/ic0_wb_i_dat\[15\]
rlabel metal3 252640 406844 252640 406844 0 mprj/ic0_wb_i_dat\[1\]
rlabel metal2 251206 412811 251206 412811 0 mprj/ic0_wb_i_dat\[2\]
rlabel metal2 251206 417333 251206 417333 0 mprj/ic0_wb_i_dat\[3\]
rlabel metal3 252318 422756 252318 422756 0 mprj/ic0_wb_i_dat\[4\]
rlabel metal2 251298 427091 251298 427091 0 mprj/ic0_wb_i_dat\[5\]
rlabel metal2 251206 432259 251206 432259 0 mprj/ic0_wb_i_dat\[6\]
rlabel metal2 231794 396746 231794 396746 0 mprj/ic0_wb_i_dat\[7\]
rlabel metal2 251206 441983 251206 441983 0 mprj/ic0_wb_i_dat\[8\]
rlabel metal2 251206 447185 251206 447185 0 mprj/ic0_wb_i_dat\[9\]
rlabel metal2 231242 373286 231242 373286 0 mprj/ic0_wb_sel\[0\]
rlabel metal2 251206 407609 251206 407609 0 mprj/ic0_wb_sel\[1\]
rlabel metal1 251804 388450 251804 388450 0 mprj/ic0_wb_stb
rlabel metal2 251206 395267 251206 395267 0 mprj/ic0_wb_we
rlabel metal3 252824 533188 252824 533188 0 mprj/ic1_clk
rlabel metal2 251206 535551 251206 535551 0 mprj/ic1_mem_ack
rlabel metal2 251206 546567 251206 546567 0 mprj/ic1_mem_addr\[0\]
rlabel metal2 251206 597805 251206 597805 0 mprj/ic1_mem_addr\[10\]
rlabel metal3 252778 602956 252778 602956 0 mprj/ic1_mem_addr\[11\]
rlabel metal2 251206 607529 251206 607529 0 mprj/ic1_mem_addr\[12\]
rlabel via2 251206 612765 251206 612765 0 mprj/ic1_mem_addr\[13\]
rlabel metal2 251206 617253 251206 617253 0 mprj/ic1_mem_addr\[14\]
rlabel metal2 251206 622489 251206 622489 0 mprj/ic1_mem_addr\[15\]
rlabel metal2 251206 552415 251206 552415 0 mprj/ic1_mem_addr\[1\]
rlabel metal2 251298 558229 251298 558229 0 mprj/ic1_mem_addr\[2\]
rlabel metal2 251206 563431 251206 563431 0 mprj/ic1_mem_addr\[3\]
rlabel metal2 251206 568633 251206 568633 0 mprj/ic1_mem_addr\[4\]
rlabel metal2 251206 573155 251206 573155 0 mprj/ic1_mem_addr\[5\]
rlabel metal2 251206 578357 251206 578357 0 mprj/ic1_mem_addr\[6\]
rlabel metal2 251206 582879 251206 582879 0 mprj/ic1_mem_addr\[7\]
rlabel metal2 229954 491878 229954 491878 0 mprj/ic1_mem_addr\[8\]
rlabel metal2 251206 592603 251206 592603 0 mprj/ic1_mem_addr\[9\]
rlabel metal2 233082 437716 233082 437716 0 mprj/ic1_mem_cache_flush
rlabel metal2 232990 464984 232990 464984 0 mprj/ic1_mem_data\[0\]
rlabel metal2 251206 599131 251206 599131 0 mprj/ic1_mem_data\[10\]
rlabel metal2 251206 603653 251206 603653 0 mprj/ic1_mem_data\[11\]
rlabel metal2 229862 505750 229862 505750 0 mprj/ic1_mem_data\[12\]
rlabel metal2 251298 613411 251298 613411 0 mprj/ic1_mem_data\[13\]
rlabel metal2 251206 618579 251206 618579 0 mprj/ic1_mem_data\[14\]
rlabel via2 251206 623781 251206 623781 0 mprj/ic1_mem_data\[15\]
rlabel metal2 231334 517480 231334 517480 0 mprj/ic1_mem_data\[16\]
rlabel metal2 231242 518126 231242 518126 0 mprj/ic1_mem_data\[17\]
rlabel metal2 251206 629595 251206 629595 0 mprj/ic1_mem_data\[18\]
rlabel metal2 232622 520234 232622 520234 0 mprj/ic1_mem_data\[19\]
rlabel metal2 232898 468520 232898 468520 0 mprj/ic1_mem_data\[1\]
rlabel metal2 251206 632213 251206 632213 0 mprj/ic1_mem_data\[20\]
rlabel metal2 251206 633131 251206 633131 0 mprj/ic1_mem_data\[21\]
rlabel metal2 251298 634117 251298 634117 0 mprj/ic1_mem_data\[22\]
rlabel metal2 251206 635409 251206 635409 0 mprj/ic1_mem_data\[23\]
rlabel metal3 252042 637228 252042 637228 0 mprj/ic1_mem_data\[24\]
rlabel metal2 251206 638027 251206 638027 0 mprj/ic1_mem_data\[25\]
rlabel metal2 251206 639319 251206 639319 0 mprj/ic1_mem_data\[26\]
rlabel metal2 251206 640611 251206 640611 0 mprj/ic1_mem_data\[27\]
rlabel metal2 251206 641937 251206 641937 0 mprj/ic1_mem_data\[28\]
rlabel metal2 251206 643229 251206 643229 0 mprj/ic1_mem_data\[29\]
rlabel metal2 251206 559521 251206 559521 0 mprj/ic1_mem_data\[2\]
rlabel metal2 234002 529176 234002 529176 0 mprj/ic1_mem_data\[30\]
rlabel metal2 234186 529176 234186 529176 0 mprj/ic1_mem_data\[31\]
rlabel metal2 251206 564723 251206 564723 0 mprj/ic1_mem_data\[3\]
rlabel metal2 234370 478856 234370 478856 0 mprj/ic1_mem_data\[4\]
rlabel metal2 231426 482290 231426 482290 0 mprj/ic1_mem_data\[5\]
rlabel metal1 250332 579734 250332 579734 0 mprj/ic1_mem_data\[6\]
rlabel metal2 251206 584171 251206 584171 0 mprj/ic1_mem_data\[7\]
rlabel metal2 251206 589407 251206 589407 0 mprj/ic1_mem_data\[8\]
rlabel metal2 251206 593895 251206 593895 0 mprj/ic1_mem_data\[9\]
rlabel metal2 235750 457470 235750 457470 0 mprj/ic1_mem_ppl_submit
rlabel metal2 251206 538781 251206 538781 0 mprj/ic1_mem_req
rlabel metal2 235842 456756 235842 456756 0 mprj/ic1_rst
rlabel metal2 251206 540073 251206 540073 0 mprj/ic1_wb_ack
rlabel metal2 235474 465052 235474 465052 0 mprj/ic1_wb_adr\[0\]
rlabel metal2 251206 600423 251206 600423 0 mprj/ic1_wb_adr\[10\]
rlabel metal2 251206 604945 251206 604945 0 mprj/ic1_wb_adr\[11\]
rlabel metal2 229770 506396 229770 506396 0 mprj/ic1_wb_adr\[12\]
rlabel metal2 235290 509150 235290 509150 0 mprj/ic1_wb_adr\[13\]
rlabel metal2 251206 619871 251206 619871 0 mprj/ic1_wb_adr\[14\]
rlabel metal2 251298 624427 251298 624427 0 mprj/ic1_wb_adr\[15\]
rlabel metal2 236946 469812 236946 469812 0 mprj/ic1_wb_adr\[1\]
rlabel metal2 251206 560813 251206 560813 0 mprj/ic1_wb_adr\[2\]
rlabel metal2 251206 566049 251206 566049 0 mprj/ic1_wb_adr\[3\]
rlabel metal2 238326 479536 238326 479536 0 mprj/ic1_wb_adr\[4\]
rlabel metal2 251206 575773 251206 575773 0 mprj/ic1_wb_adr\[5\]
rlabel metal2 251206 580295 251206 580295 0 mprj/ic1_wb_adr\[6\]
rlabel metal2 251206 585497 251206 585497 0 mprj/ic1_wb_adr\[7\]
rlabel via2 251206 590733 251206 590733 0 mprj/ic1_wb_adr\[8\]
rlabel metal2 251206 595221 251206 595221 0 mprj/ic1_wb_adr\[9\]
rlabel metal1 250378 540974 250378 540974 0 mprj/ic1_wb_cyc
rlabel metal3 252180 542980 252180 542980 0 mprj/ic1_wb_err
rlabel metal2 251206 549797 251206 549797 0 mprj/ic1_wb_i_dat\[0\]
rlabel metal1 250240 601698 250240 601698 0 mprj/ic1_wb_i_dat\[10\]
rlabel metal3 252088 606628 252088 606628 0 mprj/ic1_wb_i_dat\[11\]
rlabel metal2 238142 507144 238142 507144 0 mprj/ic1_wb_i_dat\[12\]
rlabel metal2 251206 615961 251206 615961 0 mprj/ic1_wb_i_dat\[13\]
rlabel metal2 251206 621163 251206 621163 0 mprj/ic1_wb_i_dat\[14\]
rlabel metal2 251206 625685 251206 625685 0 mprj/ic1_wb_i_dat\[15\]
rlabel metal2 251206 556325 251206 556325 0 mprj/ic1_wb_i_dat\[1\]
rlabel metal2 251206 562139 251206 562139 0 mprj/ic1_wb_i_dat\[2\]
rlabel metal2 251206 567341 251206 567341 0 mprj/ic1_wb_i_dat\[3\]
rlabel metal2 251206 571863 251206 571863 0 mprj/ic1_wb_i_dat\[4\]
rlabel metal1 250378 577014 250378 577014 0 mprj/ic1_wb_i_dat\[5\]
rlabel metal2 251206 581587 251206 581587 0 mprj/ic1_wb_i_dat\[6\]
rlabel metal3 252134 587044 252134 587044 0 mprj/ic1_wb_i_dat\[7\]
rlabel metal2 251298 591311 251298 591311 0 mprj/ic1_wb_i_dat\[8\]
rlabel metal3 252870 596836 252870 596836 0 mprj/ic1_wb_i_dat\[9\]
rlabel metal2 251206 551089 251206 551089 0 mprj/ic1_wb_sel\[0\]
rlabel via2 251206 557651 251206 557651 0 mprj/ic1_wb_sel\[1\]
rlabel metal2 251206 543983 251206 543983 0 mprj/ic1_wb_stb
rlabel metal2 251206 545275 251206 545275 0 mprj/ic1_wb_we
rlabel metal2 159084 270028 159084 270028 0 mprj/inner_clock
rlabel metal2 160786 270028 160786 270028 0 mprj/inner_disable
rlabel metal2 161260 131852 161260 131852 0 mprj/inner_embed_mode
rlabel metal2 162580 270028 162580 270028 0 mprj/inner_ext_irq
rlabel metal2 160340 270028 160340 270028 0 mprj/inner_reset
rlabel metal2 163224 270028 163224 270028 0 mprj/inner_wb_4_burst
rlabel metal2 164328 270028 164328 270028 0 mprj/inner_wb_8_burst
rlabel metal2 164880 270028 164880 270028 0 mprj/inner_wb_ack
rlabel metal1 168728 137326 168728 137326 0 mprj/inner_wb_adr\[0\]
rlabel metal1 195086 140726 195086 140726 0 mprj/inner_wb_adr\[10\]
rlabel metal2 198000 270028 198000 270028 0 mprj/inner_wb_adr\[11\]
rlabel metal2 200484 270028 200484 270028 0 mprj/inner_wb_adr\[12\]
rlabel metal2 203152 270028 203152 270028 0 mprj/inner_wb_adr\[13\]
rlabel metal2 205728 270028 205728 270028 0 mprj/inner_wb_adr\[14\]
rlabel metal2 208120 270028 208120 270028 0 mprj/inner_wb_adr\[15\]
rlabel metal2 210420 270028 210420 270028 0 mprj/inner_wb_adr\[16\]
rlabel metal2 211386 270028 211386 270028 0 mprj/inner_wb_adr\[17\]
rlabel metal2 212076 270028 212076 270028 0 mprj/inner_wb_adr\[18\]
rlabel metal2 212904 270028 212904 270028 0 mprj/inner_wb_adr\[19\]
rlabel metal2 172608 270028 172608 270028 0 mprj/inner_wb_adr\[1\]
rlabel metal2 214008 270028 214008 270028 0 mprj/inner_wb_adr\[20\]
rlabel metal2 214560 270028 214560 270028 0 mprj/inner_wb_adr\[21\]
rlabel metal2 215572 270028 215572 270028 0 mprj/inner_wb_adr\[22\]
rlabel metal1 215786 139910 215786 139910 0 mprj/inner_wb_adr\[23\]
rlabel metal2 175644 270028 175644 270028 0 mprj/inner_wb_adr\[2\]
rlabel metal2 178312 270028 178312 270028 0 mprj/inner_wb_adr\[3\]
rlabel metal2 180888 270028 180888 270028 0 mprj/inner_wb_adr\[4\]
rlabel metal2 183280 270028 183280 270028 0 mprj/inner_wb_adr\[5\]
rlabel metal2 185580 270028 185580 270028 0 mprj/inner_wb_adr\[6\]
rlabel metal2 188064 270028 188064 270028 0 mprj/inner_wb_adr\[7\]
rlabel metal2 190732 270028 190732 270028 0 mprj/inner_wb_adr\[8\]
rlabel metal2 193308 270028 193308 270028 0 mprj/inner_wb_adr\[9\]
rlabel metal2 165846 270028 165846 270028 0 mprj/inner_wb_cyc
rlabel metal2 166720 270028 166720 270028 0 mprj/inner_wb_err
rlabel metal2 170032 270028 170032 270028 0 mprj/inner_wb_i_dat\[0\]
rlabel metal2 196344 270028 196344 270028 0 mprj/inner_wb_i_dat\[10\]
rlabel metal2 198966 270028 198966 270028 0 mprj/inner_wb_i_dat\[11\]
rlabel metal2 201588 270028 201588 270028 0 mprj/inner_wb_i_dat\[12\]
rlabel metal1 203366 137326 203366 137326 0 mprj/inner_wb_i_dat\[13\]
rlabel metal2 206280 270028 206280 270028 0 mprj/inner_wb_i_dat\[14\]
rlabel metal2 208764 270028 208764 270028 0 mprj/inner_wb_i_dat\[15\]
rlabel metal2 173160 270028 173160 270028 0 mprj/inner_wb_i_dat\[1\]
rlabel metal2 176794 270028 176794 270028 0 mprj/inner_wb_i_dat\[2\]
rlabel metal1 178526 140454 178526 140454 0 mprj/inner_wb_i_dat\[3\]
rlabel metal2 181440 270028 181440 270028 0 mprj/inner_wb_i_dat\[4\]
rlabel metal2 183924 270028 183924 270028 0 mprj/inner_wb_i_dat\[5\]
rlabel metal2 186592 270028 186592 270028 0 mprj/inner_wb_i_dat\[6\]
rlabel metal2 189168 270028 189168 270028 0 mprj/inner_wb_i_dat\[7\]
rlabel metal1 190946 137326 190946 137326 0 mprj/inner_wb_i_dat\[8\]
rlabel metal2 193860 270028 193860 270028 0 mprj/inner_wb_i_dat\[9\]
rlabel metal1 170246 137326 170246 137326 0 mprj/inner_wb_o_dat\[0\]
rlabel metal2 197448 270028 197448 270028 0 mprj/inner_wb_o_dat\[10\]
rlabel metal2 199840 270028 199840 270028 0 mprj/inner_wb_o_dat\[11\]
rlabel metal2 202140 270028 202140 270028 0 mprj/inner_wb_o_dat\[12\]
rlabel metal2 204624 270028 204624 270028 0 mprj/inner_wb_o_dat\[13\]
rlabel metal2 207246 270028 207246 270028 0 mprj/inner_wb_o_dat\[14\]
rlabel metal2 209868 270028 209868 270028 0 mprj/inner_wb_o_dat\[15\]
rlabel metal2 174172 270028 174172 270028 0 mprj/inner_wb_o_dat\[1\]
rlabel metal1 177008 137326 177008 137326 0 mprj/inner_wb_o_dat\[2\]
rlabel metal2 179784 270028 179784 270028 0 mprj/inner_wb_o_dat\[3\]
rlabel metal2 182406 270028 182406 270028 0 mprj/inner_wb_o_dat\[4\]
rlabel metal2 185028 270028 185028 270028 0 mprj/inner_wb_o_dat\[5\]
rlabel metal1 186806 140658 186806 140658 0 mprj/inner_wb_o_dat\[6\]
rlabel metal2 189720 270028 189720 270028 0 mprj/inner_wb_o_dat\[7\]
rlabel metal2 192204 270028 192204 270028 0 mprj/inner_wb_o_dat\[8\]
rlabel metal2 194872 270028 194872 270028 0 mprj/inner_wb_o_dat\[9\]
rlabel metal2 171504 270028 171504 270028 0 mprj/inner_wb_sel\[0\]
rlabel metal1 174386 139434 174386 139434 0 mprj/inner_wb_sel\[1\]
rlabel metal2 167364 270028 167364 270028 0 mprj/inner_wb_stb
rlabel metal2 168514 270028 168514 270028 0 mprj/inner_wb_we
rlabel metal2 154974 57103 154974 57103 0 mprj/iram_addr\[0\]
rlabel metal3 133860 40577 133860 40577 0 mprj/iram_addr\[1\]
rlabel metal3 133860 47823 133860 47823 0 mprj/iram_addr\[2\]
rlabel metal3 133860 56081 133860 56081 0 mprj/iram_addr\[3\]
rlabel metal3 133860 63833 133860 63833 0 mprj/iram_addr\[4\]
rlabel metal3 133860 71449 133860 71449 0 mprj/iram_addr\[5\]
rlabel metal3 133860 79337 133860 79337 0 mprj/iram_addr\[6\]
rlabel metal3 133860 27453 133860 27453 0 mprj/iram_clk
rlabel metal2 154974 59449 154974 59449 0 mprj/iram_i_data\[0\]
rlabel metal3 133860 102593 133860 102593 0 mprj/iram_i_data\[10\]
rlabel metal3 133860 107489 133860 107489 0 mprj/iram_i_data\[11\]
rlabel metal3 156776 116620 156776 116620 0 mprj/iram_i_data\[12\]
rlabel metal3 133860 118029 133860 118029 0 mprj/iram_i_data\[13\]
rlabel metal3 133860 123265 133860 123265 0 mprj/iram_i_data\[14\]
rlabel metal3 133860 127995 133860 127995 0 mprj/iram_i_data\[15\]
rlabel metal3 133860 43161 133860 43161 0 mprj/iram_i_data\[1\]
rlabel metal3 133860 50777 133860 50777 0 mprj/iram_i_data\[2\]
rlabel metal3 133860 58665 133860 58665 0 mprj/iram_i_data\[3\]
rlabel metal2 154974 81889 154974 81889 0 mprj/iram_i_data\[4\]
rlabel metal3 133860 73799 133860 73799 0 mprj/iram_i_data\[5\]
rlabel metal3 133860 81921 133860 81921 0 mprj/iram_i_data\[6\]
rlabel metal2 154882 96033 154882 96033 0 mprj/iram_i_data\[7\]
rlabel metal2 154974 101065 154974 101065 0 mprj/iram_i_data\[8\]
rlabel metal3 133860 97425 133860 97425 0 mprj/iram_i_data\[9\]
rlabel metal3 133860 37789 133860 37789 0 mprj/iram_o_data\[0\]
rlabel metal3 133860 104807 133860 104807 0 mprj/iram_o_data\[10\]
rlabel metal3 156454 114716 156454 114716 0 mprj/iram_o_data\[11\]
rlabel metal3 133860 115377 133860 115377 0 mprj/iram_o_data\[12\]
rlabel metal3 133860 120613 133860 120613 0 mprj/iram_o_data\[13\]
rlabel metal3 133860 125479 133860 125479 0 mprj/iram_o_data\[14\]
rlabel metal3 133860 130579 133860 130579 0 mprj/iram_o_data\[15\]
rlabel metal3 133860 45473 133860 45473 0 mprj/iram_o_data\[1\]
rlabel metal3 133860 53361 133860 53361 0 mprj/iram_o_data\[2\]
rlabel metal3 133860 61249 133860 61249 0 mprj/iram_o_data\[3\]
rlabel metal3 133860 68797 133860 68797 0 mprj/iram_o_data\[4\]
rlabel metal3 133860 76753 133860 76753 0 mprj/iram_o_data\[5\]
rlabel metal2 154974 95455 154974 95455 0 mprj/iram_o_data\[6\]
rlabel metal2 154974 99433 154974 99433 0 mprj/iram_o_data\[7\]
rlabel metal3 133860 94841 133860 94841 0 mprj/iram_o_data\[8\]
rlabel metal3 133860 99941 133860 99941 0 mprj/iram_o_data\[9\]
rlabel metal2 154974 55471 154974 55471 0 mprj/iram_we
rlabel metal2 579731 340 579731 340 0 user_clock2
rlabel metal2 581026 12927 581026 12927 0 user_irq[0]
rlabel metal2 581985 340 581985 340 0 user_irq[1]
rlabel metal2 583418 1894 583418 1894 0 user_irq[2]
rlabel metal2 598 1894 598 1894 0 wb_clk_i
rlabel metal2 1557 340 1557 340 0 wb_rst_i
rlabel metal2 2898 8116 2898 8116 0 wbs_ack_o
rlabel metal1 83720 18598 83720 18598 0 wbs_adr_i[0]
rlabel metal2 47649 340 47649 340 0 wbs_adr_i[10]
rlabel metal2 51237 340 51237 340 0 wbs_adr_i[11]
rlabel metal1 108376 21590 108376 21590 0 wbs_adr_i[12]
rlabel metal2 58006 20469 58006 20469 0 wbs_adr_i[13]
rlabel metal2 61863 340 61863 340 0 wbs_adr_i[14]
rlabel metal2 65313 340 65313 340 0 wbs_adr_i[15]
rlabel metal1 116886 18802 116886 18802 0 wbs_adr_i[16]
rlabel metal1 114724 24582 114724 24582 0 wbs_adr_i[17]
rlabel metal2 76077 340 76077 340 0 wbs_adr_i[18]
rlabel metal2 79481 340 79481 340 0 wbs_adr_i[19]
rlabel metal2 12137 340 12137 340 0 wbs_adr_i[1]
rlabel metal2 82846 18327 82846 18327 0 wbs_adr_i[20]
rlabel metal2 86657 340 86657 340 0 wbs_adr_i[21]
rlabel metal2 90153 340 90153 340 0 wbs_adr_i[22]
rlabel metal2 93886 18990 93886 18990 0 wbs_adr_i[23]
rlabel metal2 97474 5362 97474 5362 0 wbs_adr_i[24]
rlabel metal2 100917 340 100917 340 0 wbs_adr_i[25]
rlabel metal2 104321 340 104321 340 0 wbs_adr_i[26]
rlabel metal1 133124 24038 133124 24038 0 wbs_adr_i[27]
rlabel metal2 111642 2727 111642 2727 0 wbs_adr_i[28]
rlabel metal2 114993 340 114993 340 0 wbs_adr_i[29]
rlabel metal2 17066 1928 17066 1928 0 wbs_adr_i[2]
rlabel metal2 118818 5430 118818 5430 0 wbs_adr_i[30]
rlabel metal2 121486 19143 121486 19143 0 wbs_adr_i[31]
rlabel metal2 20746 17562 20746 17562 0 wbs_adr_i[3]
rlabel metal2 26397 340 26397 340 0 wbs_adr_i[4]
rlabel metal2 30130 6756 30130 6756 0 wbs_adr_i[5]
rlabel metal1 97566 17238 97566 17238 0 wbs_adr_i[6]
rlabel metal2 36977 340 36977 340 0 wbs_adr_i[7]
rlabel metal2 40710 3339 40710 3339 0 wbs_adr_i[8]
rlabel metal2 44298 2642 44298 2642 0 wbs_adr_i[9]
rlabel metal2 3857 340 3857 340 0 wbs_cyc_i
rlabel metal2 8786 6042 8786 6042 0 wbs_dat_i[0]
rlabel metal2 48990 4002 48990 4002 0 wbs_dat_i[10]
rlabel metal2 52578 3254 52578 3254 0 wbs_dat_i[11]
rlabel metal2 56074 2591 56074 2591 0 wbs_dat_i[12]
rlabel metal2 59662 4036 59662 4036 0 wbs_dat_i[13]
rlabel metal2 63250 6790 63250 6790 0 wbs_dat_i[14]
rlabel metal2 66746 3288 66746 3288 0 wbs_dat_i[15]
rlabel metal2 70097 340 70097 340 0 wbs_dat_i[16]
rlabel metal2 73830 2659 73830 2659 0 wbs_dat_i[17]
rlabel metal2 77418 6110 77418 6110 0 wbs_dat_i[18]
rlabel metal2 80914 7436 80914 7436 0 wbs_dat_i[19]
rlabel metal2 13570 7402 13570 7402 0 wbs_dat_i[1]
rlabel metal2 84502 4104 84502 4104 0 wbs_dat_i[20]
rlabel metal2 87761 340 87761 340 0 wbs_dat_i[21]
rlabel metal2 91586 7487 91586 7487 0 wbs_dat_i[22]
rlabel metal2 94937 340 94937 340 0 wbs_dat_i[23]
rlabel metal2 98433 340 98433 340 0 wbs_dat_i[24]
rlabel metal2 102258 8218 102258 8218 0 wbs_dat_i[25]
rlabel metal2 105754 3322 105754 3322 0 wbs_dat_i[26]
rlabel metal2 109342 4699 109342 4699 0 wbs_dat_i[27]
rlabel metal2 112838 4767 112838 4767 0 wbs_dat_i[28]
rlabel metal2 116426 8286 116426 8286 0 wbs_dat_i[29]
rlabel metal2 18262 2676 18262 2676 0 wbs_dat_i[2]
rlabel metal2 119922 4716 119922 4716 0 wbs_dat_i[30]
rlabel metal2 123273 340 123273 340 0 wbs_dat_i[31]
rlabel metal2 23046 4631 23046 4631 0 wbs_dat_i[3]
rlabel metal2 27738 3968 27738 3968 0 wbs_dat_i[4]
rlabel metal2 31326 2608 31326 2608 0 wbs_dat_i[5]
rlabel metal2 34677 340 34677 340 0 wbs_dat_i[6]
rlabel metal2 38410 3271 38410 3271 0 wbs_dat_i[7]
rlabel metal2 41906 8099 41906 8099 0 wbs_dat_i[8]
rlabel metal2 45494 4648 45494 4648 0 wbs_dat_i[9]
rlabel metal2 9837 340 9837 340 0 wbs_dat_o[0]
rlabel metal1 106582 21522 106582 21522 0 wbs_dat_o[10]
rlabel metal2 53537 340 53537 340 0 wbs_dat_o[11]
rlabel metal2 57270 2132 57270 2132 0 wbs_dat_o[12]
rlabel metal2 60858 8864 60858 8864 0 wbs_dat_o[13]
rlabel metal2 64354 4070 64354 4070 0 wbs_dat_o[14]
rlabel metal2 67797 340 67797 340 0 wbs_dat_o[15]
rlabel metal2 71530 4682 71530 4682 0 wbs_dat_o[16]
rlabel metal2 75026 6671 75026 6671 0 wbs_dat_o[17]
rlabel metal2 78423 340 78423 340 0 wbs_dat_o[18]
rlabel metal2 81873 340 81873 340 0 wbs_dat_o[19]
rlabel metal2 14529 340 14529 340 0 wbs_dat_o[1]
rlabel metal1 125948 22950 125948 22950 0 wbs_dat_o[20]
rlabel metal2 133170 25772 133170 25772 0 wbs_dat_o[21]
rlabel metal2 134826 25109 134826 25109 0 wbs_dat_o[22]
rlabel metal2 96041 340 96041 340 0 wbs_dat_o[23]
rlabel metal2 99866 6144 99866 6144 0 wbs_dat_o[24]
rlabel metal2 103362 1860 103362 1860 0 wbs_dat_o[25]
rlabel metal2 134642 25500 134642 25500 0 wbs_dat_o[26]
rlabel metal1 134090 23902 134090 23902 0 wbs_dat_o[27]
rlabel metal2 114034 7504 114034 7504 0 wbs_dat_o[28]
rlabel metal2 117622 1826 117622 1826 0 wbs_dat_o[29]
rlabel metal2 19458 1928 19458 1928 0 wbs_dat_o[2]
rlabel metal2 120881 340 120881 340 0 wbs_dat_o[30]
rlabel metal2 124706 2234 124706 2234 0 wbs_dat_o[31]
rlabel metal2 24242 1962 24242 1962 0 wbs_dat_o[3]
rlabel metal2 28697 340 28697 340 0 wbs_dat_o[4]
rlabel metal2 32193 340 32193 340 0 wbs_dat_o[5]
rlabel metal2 35926 20333 35926 20333 0 wbs_dat_o[6]
rlabel metal2 39369 340 39369 340 0 wbs_dat_o[7]
rlabel metal2 43102 2064 43102 2064 0 wbs_dat_o[8]
rlabel metal1 102626 24242 102626 24242 0 wbs_dat_o[9]
rlabel metal2 134550 25704 134550 25704 0 wbs_sel_i[0]
rlabel metal1 86848 21454 86848 21454 0 wbs_sel_i[1]
rlabel metal2 20417 340 20417 340 0 wbs_sel_i[2]
rlabel metal2 25346 2098 25346 2098 0 wbs_sel_i[3]
rlabel metal2 4186 18973 4186 18973 0 wbs_stb_i
rlabel metal2 6486 1996 6486 1996 0 wbs_we_i
<< properties >>
string FIXED_BBOX 0 0 584000 704000
<< end >>
