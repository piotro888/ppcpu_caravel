// This is the unpowered netlist.
module core1 (i_clk,
    i_disable,
    i_irq,
    i_mc_core_int,
    i_mem_ack,
    i_mem_exception,
    i_req_data_valid,
    i_rst,
    o_c_data_page,
    o_c_instr_long,
    o_c_instr_page,
    o_icache_flush,
    o_mem_long,
    o_mem_req,
    o_mem_we,
    o_req_active,
    o_req_ppl_submit,
    sr_bus_we,
    dbg_pc,
    dbg_r0,
    i_core_int_sreg,
    i_mem_data,
    i_req_data,
    o_instr_long_addr,
    o_mem_addr,
    o_mem_addr_high,
    o_mem_data,
    o_mem_sel,
    o_req_addr,
    sr_bus_addr,
    sr_bus_data_o);
 input i_clk;
 input i_disable;
 input i_irq;
 input i_mc_core_int;
 input i_mem_ack;
 input i_mem_exception;
 input i_req_data_valid;
 input i_rst;
 output o_c_data_page;
 output o_c_instr_long;
 output o_c_instr_page;
 output o_icache_flush;
 output o_mem_long;
 output o_mem_req;
 output o_mem_we;
 output o_req_active;
 output o_req_ppl_submit;
 output sr_bus_we;
 output [15:0] dbg_pc;
 output [15:0] dbg_r0;
 input [15:0] i_core_int_sreg;
 input [15:0] i_mem_data;
 input [31:0] i_req_data;
 output [7:0] o_instr_long_addr;
 output [15:0] o_mem_addr;
 output [7:0] o_mem_addr_high;
 output [15:0] o_mem_data;
 output [1:0] o_mem_sel;
 output [15:0] o_req_addr;
 output [15:0] sr_bus_addr;
 output [15:0] sr_bus_data_o;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1074_;
 wire _1075_;
 wire _1076_;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire _1080_;
 wire _1081_;
 wire _1082_;
 wire _1083_;
 wire _1084_;
 wire _1085_;
 wire _1086_;
 wire _1087_;
 wire _1088_;
 wire _1089_;
 wire _1090_;
 wire _1091_;
 wire _1092_;
 wire _1093_;
 wire _1094_;
 wire _1095_;
 wire _1096_;
 wire _1097_;
 wire _1098_;
 wire _1099_;
 wire _1100_;
 wire _1101_;
 wire _1102_;
 wire _1103_;
 wire _1104_;
 wire _1105_;
 wire _1106_;
 wire _1107_;
 wire _1108_;
 wire _1109_;
 wire _1110_;
 wire _1111_;
 wire _1112_;
 wire _1113_;
 wire _1114_;
 wire _1115_;
 wire _1116_;
 wire _1117_;
 wire _1118_;
 wire _1119_;
 wire _1120_;
 wire _1121_;
 wire _1122_;
 wire _1123_;
 wire _1124_;
 wire _1125_;
 wire _1126_;
 wire _1127_;
 wire _1128_;
 wire _1129_;
 wire _1130_;
 wire _1131_;
 wire _1132_;
 wire _1133_;
 wire _1134_;
 wire _1135_;
 wire _1136_;
 wire _1137_;
 wire _1138_;
 wire _1139_;
 wire _1140_;
 wire _1141_;
 wire _1142_;
 wire _1143_;
 wire _1144_;
 wire _1145_;
 wire _1146_;
 wire _1147_;
 wire _1148_;
 wire _1149_;
 wire _1150_;
 wire _1151_;
 wire _1152_;
 wire _1153_;
 wire _1154_;
 wire _1155_;
 wire _1156_;
 wire _1157_;
 wire _1158_;
 wire _1159_;
 wire _1160_;
 wire _1161_;
 wire _1162_;
 wire _1163_;
 wire _1164_;
 wire _1165_;
 wire _1166_;
 wire _1167_;
 wire _1168_;
 wire _1169_;
 wire _1170_;
 wire _1171_;
 wire _1172_;
 wire _1173_;
 wire _1174_;
 wire _1175_;
 wire _1176_;
 wire _1177_;
 wire _1178_;
 wire _1179_;
 wire _1180_;
 wire _1181_;
 wire _1182_;
 wire _1183_;
 wire _1184_;
 wire _1185_;
 wire _1186_;
 wire _1187_;
 wire _1188_;
 wire _1189_;
 wire _1190_;
 wire _1191_;
 wire _1192_;
 wire _1193_;
 wire _1194_;
 wire _1195_;
 wire _1196_;
 wire _1197_;
 wire _1198_;
 wire _1199_;
 wire _1200_;
 wire _1201_;
 wire _1202_;
 wire _1203_;
 wire _1204_;
 wire _1205_;
 wire _1206_;
 wire _1207_;
 wire _1208_;
 wire _1209_;
 wire _1210_;
 wire _1211_;
 wire _1212_;
 wire _1213_;
 wire _1214_;
 wire _1215_;
 wire _1216_;
 wire _1217_;
 wire _1218_;
 wire _1219_;
 wire _1220_;
 wire _1221_;
 wire _1222_;
 wire _1223_;
 wire _1224_;
 wire _1225_;
 wire _1226_;
 wire _1227_;
 wire _1228_;
 wire _1229_;
 wire _1230_;
 wire _1231_;
 wire _1232_;
 wire _1233_;
 wire _1234_;
 wire _1235_;
 wire _1236_;
 wire _1237_;
 wire _1238_;
 wire _1239_;
 wire _1240_;
 wire _1241_;
 wire _1242_;
 wire _1243_;
 wire _1244_;
 wire _1245_;
 wire _1246_;
 wire _1247_;
 wire _1248_;
 wire _1249_;
 wire _1250_;
 wire _1251_;
 wire _1252_;
 wire _1253_;
 wire _1254_;
 wire _1255_;
 wire _1256_;
 wire _1257_;
 wire _1258_;
 wire _1259_;
 wire _1260_;
 wire _1261_;
 wire _1262_;
 wire _1263_;
 wire _1264_;
 wire _1265_;
 wire _1266_;
 wire _1267_;
 wire _1268_;
 wire _1269_;
 wire _1270_;
 wire _1271_;
 wire _1272_;
 wire _1273_;
 wire _1274_;
 wire _1275_;
 wire _1276_;
 wire _1277_;
 wire _1278_;
 wire _1279_;
 wire _1280_;
 wire _1281_;
 wire _1282_;
 wire _1283_;
 wire _1284_;
 wire _1285_;
 wire _1286_;
 wire _1287_;
 wire _1288_;
 wire _1289_;
 wire _1290_;
 wire _1291_;
 wire _1292_;
 wire _1293_;
 wire _1294_;
 wire _1295_;
 wire _1296_;
 wire _1297_;
 wire _1298_;
 wire _1299_;
 wire _1300_;
 wire _1301_;
 wire _1302_;
 wire _1303_;
 wire _1304_;
 wire _1305_;
 wire _1306_;
 wire _1307_;
 wire _1308_;
 wire _1309_;
 wire _1310_;
 wire _1311_;
 wire _1312_;
 wire _1313_;
 wire _1314_;
 wire _1315_;
 wire _1316_;
 wire _1317_;
 wire _1318_;
 wire _1319_;
 wire _1320_;
 wire _1321_;
 wire _1322_;
 wire _1323_;
 wire _1324_;
 wire _1325_;
 wire _1326_;
 wire _1327_;
 wire _1328_;
 wire _1329_;
 wire _1330_;
 wire _1331_;
 wire _1332_;
 wire _1333_;
 wire _1334_;
 wire _1335_;
 wire _1336_;
 wire _1337_;
 wire _1338_;
 wire _1339_;
 wire _1340_;
 wire _1341_;
 wire _1342_;
 wire _1343_;
 wire _1344_;
 wire _1345_;
 wire _1346_;
 wire _1347_;
 wire _1348_;
 wire _1349_;
 wire _1350_;
 wire _1351_;
 wire _1352_;
 wire _1353_;
 wire _1354_;
 wire _1355_;
 wire _1356_;
 wire _1357_;
 wire _1358_;
 wire _1359_;
 wire _1360_;
 wire _1361_;
 wire _1362_;
 wire _1363_;
 wire _1364_;
 wire _1365_;
 wire _1366_;
 wire _1367_;
 wire _1368_;
 wire _1369_;
 wire _1370_;
 wire _1371_;
 wire _1372_;
 wire _1373_;
 wire _1374_;
 wire _1375_;
 wire _1376_;
 wire _1377_;
 wire _1378_;
 wire _1379_;
 wire _1380_;
 wire _1381_;
 wire _1382_;
 wire _1383_;
 wire _1384_;
 wire _1385_;
 wire _1386_;
 wire _1387_;
 wire _1388_;
 wire _1389_;
 wire _1390_;
 wire _1391_;
 wire _1392_;
 wire _1393_;
 wire _1394_;
 wire _1395_;
 wire _1396_;
 wire _1397_;
 wire _1398_;
 wire _1399_;
 wire _1400_;
 wire _1401_;
 wire _1402_;
 wire _1403_;
 wire _1404_;
 wire _1405_;
 wire _1406_;
 wire _1407_;
 wire _1408_;
 wire _1409_;
 wire _1410_;
 wire _1411_;
 wire _1412_;
 wire _1413_;
 wire _1414_;
 wire _1415_;
 wire _1416_;
 wire _1417_;
 wire _1418_;
 wire _1419_;
 wire _1420_;
 wire _1421_;
 wire _1422_;
 wire _1423_;
 wire _1424_;
 wire _1425_;
 wire _1426_;
 wire _1427_;
 wire _1428_;
 wire _1429_;
 wire _1430_;
 wire _1431_;
 wire _1432_;
 wire _1433_;
 wire _1434_;
 wire _1435_;
 wire _1436_;
 wire _1437_;
 wire _1438_;
 wire _1439_;
 wire _1440_;
 wire _1441_;
 wire _1442_;
 wire _1443_;
 wire _1444_;
 wire _1445_;
 wire _1446_;
 wire _1447_;
 wire _1448_;
 wire _1449_;
 wire _1450_;
 wire _1451_;
 wire _1452_;
 wire _1453_;
 wire _1454_;
 wire _1455_;
 wire _1456_;
 wire _1457_;
 wire _1458_;
 wire _1459_;
 wire _1460_;
 wire _1461_;
 wire _1462_;
 wire _1463_;
 wire _1464_;
 wire _1465_;
 wire _1466_;
 wire _1467_;
 wire _1468_;
 wire _1469_;
 wire _1470_;
 wire _1471_;
 wire _1472_;
 wire _1473_;
 wire _1474_;
 wire _1475_;
 wire _1476_;
 wire _1477_;
 wire _1478_;
 wire _1479_;
 wire _1480_;
 wire _1481_;
 wire _1482_;
 wire _1483_;
 wire _1484_;
 wire _1485_;
 wire _1486_;
 wire _1487_;
 wire _1488_;
 wire _1489_;
 wire _1490_;
 wire _1491_;
 wire _1492_;
 wire _1493_;
 wire _1494_;
 wire _1495_;
 wire _1496_;
 wire _1497_;
 wire _1498_;
 wire _1499_;
 wire _1500_;
 wire _1501_;
 wire _1502_;
 wire _1503_;
 wire _1504_;
 wire _1505_;
 wire _1506_;
 wire _1507_;
 wire _1508_;
 wire _1509_;
 wire _1510_;
 wire _1511_;
 wire _1512_;
 wire _1513_;
 wire _1514_;
 wire _1515_;
 wire _1516_;
 wire _1517_;
 wire _1518_;
 wire _1519_;
 wire _1520_;
 wire _1521_;
 wire _1522_;
 wire _1523_;
 wire _1524_;
 wire _1525_;
 wire _1526_;
 wire _1527_;
 wire _1528_;
 wire _1529_;
 wire _1530_;
 wire _1531_;
 wire _1532_;
 wire _1533_;
 wire _1534_;
 wire _1535_;
 wire _1536_;
 wire _1537_;
 wire _1538_;
 wire _1539_;
 wire _1540_;
 wire _1541_;
 wire _1542_;
 wire _1543_;
 wire _1544_;
 wire _1545_;
 wire _1546_;
 wire _1547_;
 wire _1548_;
 wire _1549_;
 wire _1550_;
 wire _1551_;
 wire _1552_;
 wire _1553_;
 wire _1554_;
 wire _1555_;
 wire _1556_;
 wire _1557_;
 wire _1558_;
 wire _1559_;
 wire _1560_;
 wire _1561_;
 wire _1562_;
 wire _1563_;
 wire _1564_;
 wire _1565_;
 wire _1566_;
 wire _1567_;
 wire _1568_;
 wire _1569_;
 wire _1570_;
 wire _1571_;
 wire _1572_;
 wire _1573_;
 wire _1574_;
 wire _1575_;
 wire _1576_;
 wire _1577_;
 wire _1578_;
 wire _1579_;
 wire _1580_;
 wire _1581_;
 wire _1582_;
 wire _1583_;
 wire _1584_;
 wire _1585_;
 wire _1586_;
 wire _1587_;
 wire _1588_;
 wire _1589_;
 wire _1590_;
 wire _1591_;
 wire _1592_;
 wire _1593_;
 wire _1594_;
 wire _1595_;
 wire _1596_;
 wire _1597_;
 wire _1598_;
 wire _1599_;
 wire _1600_;
 wire _1601_;
 wire _1602_;
 wire _1603_;
 wire _1604_;
 wire _1605_;
 wire _1606_;
 wire _1607_;
 wire _1608_;
 wire _1609_;
 wire _1610_;
 wire _1611_;
 wire _1612_;
 wire _1613_;
 wire _1614_;
 wire _1615_;
 wire _1616_;
 wire _1617_;
 wire _1618_;
 wire _1619_;
 wire _1620_;
 wire _1621_;
 wire _1622_;
 wire _1623_;
 wire _1624_;
 wire _1625_;
 wire _1626_;
 wire _1627_;
 wire _1628_;
 wire _1629_;
 wire _1630_;
 wire _1631_;
 wire _1632_;
 wire _1633_;
 wire _1634_;
 wire _1635_;
 wire _1636_;
 wire _1637_;
 wire _1638_;
 wire _1639_;
 wire _1640_;
 wire _1641_;
 wire _1642_;
 wire _1643_;
 wire _1644_;
 wire _1645_;
 wire _1646_;
 wire _1647_;
 wire _1648_;
 wire _1649_;
 wire _1650_;
 wire _1651_;
 wire _1652_;
 wire _1653_;
 wire _1654_;
 wire _1655_;
 wire _1656_;
 wire _1657_;
 wire _1658_;
 wire _1659_;
 wire _1660_;
 wire _1661_;
 wire _1662_;
 wire _1663_;
 wire _1664_;
 wire _1665_;
 wire _1666_;
 wire _1667_;
 wire _1668_;
 wire _1669_;
 wire _1670_;
 wire _1671_;
 wire _1672_;
 wire _1673_;
 wire _1674_;
 wire _1675_;
 wire _1676_;
 wire _1677_;
 wire _1678_;
 wire _1679_;
 wire _1680_;
 wire _1681_;
 wire _1682_;
 wire _1683_;
 wire _1684_;
 wire _1685_;
 wire _1686_;
 wire _1687_;
 wire _1688_;
 wire _1689_;
 wire _1690_;
 wire _1691_;
 wire _1692_;
 wire _1693_;
 wire _1694_;
 wire _1695_;
 wire _1696_;
 wire _1697_;
 wire _1698_;
 wire _1699_;
 wire _1700_;
 wire _1701_;
 wire _1702_;
 wire _1703_;
 wire _1704_;
 wire _1705_;
 wire _1706_;
 wire _1707_;
 wire _1708_;
 wire _1709_;
 wire _1710_;
 wire _1711_;
 wire _1712_;
 wire _1713_;
 wire _1714_;
 wire _1715_;
 wire _1716_;
 wire _1717_;
 wire _1718_;
 wire _1719_;
 wire _1720_;
 wire _1721_;
 wire _1722_;
 wire _1723_;
 wire _1724_;
 wire _1725_;
 wire _1726_;
 wire _1727_;
 wire _1728_;
 wire _1729_;
 wire _1730_;
 wire _1731_;
 wire _1732_;
 wire _1733_;
 wire _1734_;
 wire _1735_;
 wire _1736_;
 wire _1737_;
 wire _1738_;
 wire _1739_;
 wire _1740_;
 wire _1741_;
 wire _1742_;
 wire _1743_;
 wire _1744_;
 wire _1745_;
 wire _1746_;
 wire _1747_;
 wire _1748_;
 wire _1749_;
 wire _1750_;
 wire _1751_;
 wire _1752_;
 wire _1753_;
 wire _1754_;
 wire _1755_;
 wire _1756_;
 wire _1757_;
 wire _1758_;
 wire _1759_;
 wire _1760_;
 wire _1761_;
 wire _1762_;
 wire _1763_;
 wire _1764_;
 wire _1765_;
 wire _1766_;
 wire _1767_;
 wire _1768_;
 wire _1769_;
 wire _1770_;
 wire _1771_;
 wire _1772_;
 wire _1773_;
 wire _1774_;
 wire _1775_;
 wire _1776_;
 wire _1777_;
 wire _1778_;
 wire _1779_;
 wire _1780_;
 wire _1781_;
 wire _1782_;
 wire _1783_;
 wire _1784_;
 wire _1785_;
 wire _1786_;
 wire _1787_;
 wire _1788_;
 wire _1789_;
 wire _1790_;
 wire _1791_;
 wire _1792_;
 wire _1793_;
 wire _1794_;
 wire _1795_;
 wire _1796_;
 wire _1797_;
 wire _1798_;
 wire _1799_;
 wire _1800_;
 wire _1801_;
 wire _1802_;
 wire _1803_;
 wire _1804_;
 wire _1805_;
 wire _1806_;
 wire _1807_;
 wire _1808_;
 wire _1809_;
 wire _1810_;
 wire _1811_;
 wire _1812_;
 wire _1813_;
 wire _1814_;
 wire _1815_;
 wire _1816_;
 wire _1817_;
 wire _1818_;
 wire _1819_;
 wire _1820_;
 wire _1821_;
 wire _1822_;
 wire _1823_;
 wire _1824_;
 wire _1825_;
 wire _1826_;
 wire _1827_;
 wire _1828_;
 wire _1829_;
 wire _1830_;
 wire _1831_;
 wire _1832_;
 wire _1833_;
 wire _1834_;
 wire _1835_;
 wire _1836_;
 wire _1837_;
 wire _1838_;
 wire _1839_;
 wire _1840_;
 wire _1841_;
 wire _1842_;
 wire _1843_;
 wire _1844_;
 wire _1845_;
 wire _1846_;
 wire _1847_;
 wire _1848_;
 wire _1849_;
 wire _1850_;
 wire _1851_;
 wire _1852_;
 wire _1853_;
 wire _1854_;
 wire _1855_;
 wire _1856_;
 wire _1857_;
 wire _1858_;
 wire _1859_;
 wire _1860_;
 wire _1861_;
 wire _1862_;
 wire _1863_;
 wire _1864_;
 wire _1865_;
 wire _1866_;
 wire _1867_;
 wire _1868_;
 wire _1869_;
 wire _1870_;
 wire _1871_;
 wire _1872_;
 wire _1873_;
 wire _1874_;
 wire _1875_;
 wire _1876_;
 wire _1877_;
 wire _1878_;
 wire _1879_;
 wire _1880_;
 wire _1881_;
 wire _1882_;
 wire _1883_;
 wire _1884_;
 wire _1885_;
 wire _1886_;
 wire _1887_;
 wire _1888_;
 wire _1889_;
 wire _1890_;
 wire _1891_;
 wire _1892_;
 wire _1893_;
 wire _1894_;
 wire _1895_;
 wire _1896_;
 wire _1897_;
 wire _1898_;
 wire _1899_;
 wire _1900_;
 wire _1901_;
 wire _1902_;
 wire _1903_;
 wire _1904_;
 wire _1905_;
 wire _1906_;
 wire _1907_;
 wire _1908_;
 wire _1909_;
 wire _1910_;
 wire _1911_;
 wire _1912_;
 wire _1913_;
 wire _1914_;
 wire _1915_;
 wire _1916_;
 wire _1917_;
 wire _1918_;
 wire _1919_;
 wire _1920_;
 wire _1921_;
 wire _1922_;
 wire _1923_;
 wire _1924_;
 wire _1925_;
 wire _1926_;
 wire _1927_;
 wire _1928_;
 wire _1929_;
 wire _1930_;
 wire _1931_;
 wire _1932_;
 wire _1933_;
 wire _1934_;
 wire _1935_;
 wire _1936_;
 wire _1937_;
 wire _1938_;
 wire _1939_;
 wire _1940_;
 wire _1941_;
 wire _1942_;
 wire _1943_;
 wire _1944_;
 wire _1945_;
 wire _1946_;
 wire _1947_;
 wire _1948_;
 wire _1949_;
 wire _1950_;
 wire _1951_;
 wire _1952_;
 wire _1953_;
 wire _1954_;
 wire _1955_;
 wire _1956_;
 wire _1957_;
 wire _1958_;
 wire _1959_;
 wire _1960_;
 wire _1961_;
 wire _1962_;
 wire _1963_;
 wire _1964_;
 wire _1965_;
 wire _1966_;
 wire _1967_;
 wire _1968_;
 wire _1969_;
 wire _1970_;
 wire _1971_;
 wire _1972_;
 wire _1973_;
 wire _1974_;
 wire _1975_;
 wire _1976_;
 wire _1977_;
 wire _1978_;
 wire _1979_;
 wire _1980_;
 wire _1981_;
 wire _1982_;
 wire _1983_;
 wire _1984_;
 wire _1985_;
 wire _1986_;
 wire _1987_;
 wire _1988_;
 wire _1989_;
 wire _1990_;
 wire _1991_;
 wire _1992_;
 wire _1993_;
 wire _1994_;
 wire _1995_;
 wire _1996_;
 wire _1997_;
 wire _1998_;
 wire _1999_;
 wire _2000_;
 wire _2001_;
 wire _2002_;
 wire _2003_;
 wire _2004_;
 wire _2005_;
 wire _2006_;
 wire _2007_;
 wire _2008_;
 wire _2009_;
 wire _2010_;
 wire _2011_;
 wire _2012_;
 wire _2013_;
 wire _2014_;
 wire _2015_;
 wire _2016_;
 wire _2017_;
 wire _2018_;
 wire _2019_;
 wire _2020_;
 wire _2021_;
 wire _2022_;
 wire _2023_;
 wire _2024_;
 wire _2025_;
 wire _2026_;
 wire _2027_;
 wire _2028_;
 wire _2029_;
 wire _2030_;
 wire _2031_;
 wire _2032_;
 wire _2033_;
 wire _2034_;
 wire _2035_;
 wire _2036_;
 wire _2037_;
 wire _2038_;
 wire _2039_;
 wire _2040_;
 wire _2041_;
 wire _2042_;
 wire _2043_;
 wire _2044_;
 wire _2045_;
 wire _2046_;
 wire _2047_;
 wire _2048_;
 wire _2049_;
 wire _2050_;
 wire _2051_;
 wire _2052_;
 wire _2053_;
 wire _2054_;
 wire _2055_;
 wire _2056_;
 wire _2057_;
 wire _2058_;
 wire _2059_;
 wire _2060_;
 wire _2061_;
 wire _2062_;
 wire _2063_;
 wire _2064_;
 wire _2065_;
 wire _2066_;
 wire _2067_;
 wire _2068_;
 wire _2069_;
 wire _2070_;
 wire _2071_;
 wire _2072_;
 wire _2073_;
 wire _2074_;
 wire _2075_;
 wire _2076_;
 wire _2077_;
 wire _2078_;
 wire _2079_;
 wire _2080_;
 wire _2081_;
 wire _2082_;
 wire _2083_;
 wire _2084_;
 wire _2085_;
 wire _2086_;
 wire _2087_;
 wire _2088_;
 wire _2089_;
 wire _2090_;
 wire _2091_;
 wire _2092_;
 wire _2093_;
 wire _2094_;
 wire _2095_;
 wire _2096_;
 wire _2097_;
 wire _2098_;
 wire _2099_;
 wire _2100_;
 wire _2101_;
 wire _2102_;
 wire _2103_;
 wire _2104_;
 wire _2105_;
 wire _2106_;
 wire _2107_;
 wire _2108_;
 wire _2109_;
 wire _2110_;
 wire _2111_;
 wire _2112_;
 wire _2113_;
 wire _2114_;
 wire _2115_;
 wire _2116_;
 wire _2117_;
 wire _2118_;
 wire _2119_;
 wire _2120_;
 wire _2121_;
 wire _2122_;
 wire _2123_;
 wire _2124_;
 wire _2125_;
 wire _2126_;
 wire _2127_;
 wire _2128_;
 wire _2129_;
 wire _2130_;
 wire _2131_;
 wire _2132_;
 wire _2133_;
 wire _2134_;
 wire _2135_;
 wire _2136_;
 wire _2137_;
 wire _2138_;
 wire _2139_;
 wire _2140_;
 wire _2141_;
 wire _2142_;
 wire _2143_;
 wire _2144_;
 wire _2145_;
 wire _2146_;
 wire _2147_;
 wire _2148_;
 wire _2149_;
 wire _2150_;
 wire _2151_;
 wire _2152_;
 wire _2153_;
 wire _2154_;
 wire _2155_;
 wire _2156_;
 wire _2157_;
 wire _2158_;
 wire _2159_;
 wire _2160_;
 wire _2161_;
 wire _2162_;
 wire _2163_;
 wire _2164_;
 wire _2165_;
 wire _2166_;
 wire _2167_;
 wire _2168_;
 wire _2169_;
 wire _2170_;
 wire _2171_;
 wire _2172_;
 wire _2173_;
 wire _2174_;
 wire _2175_;
 wire _2176_;
 wire _2177_;
 wire _2178_;
 wire _2179_;
 wire _2180_;
 wire _2181_;
 wire _2182_;
 wire _2183_;
 wire _2184_;
 wire _2185_;
 wire _2186_;
 wire _2187_;
 wire _2188_;
 wire _2189_;
 wire _2190_;
 wire _2191_;
 wire _2192_;
 wire _2193_;
 wire _2194_;
 wire _2195_;
 wire _2196_;
 wire _2197_;
 wire _2198_;
 wire _2199_;
 wire _2200_;
 wire _2201_;
 wire _2202_;
 wire _2203_;
 wire _2204_;
 wire _2205_;
 wire _2206_;
 wire _2207_;
 wire _2208_;
 wire _2209_;
 wire _2210_;
 wire _2211_;
 wire _2212_;
 wire _2213_;
 wire _2214_;
 wire _2215_;
 wire _2216_;
 wire _2217_;
 wire _2218_;
 wire _2219_;
 wire _2220_;
 wire _2221_;
 wire _2222_;
 wire _2223_;
 wire _2224_;
 wire _2225_;
 wire _2226_;
 wire _2227_;
 wire _2228_;
 wire _2229_;
 wire _2230_;
 wire _2231_;
 wire _2232_;
 wire _2233_;
 wire _2234_;
 wire _2235_;
 wire _2236_;
 wire _2237_;
 wire _2238_;
 wire _2239_;
 wire _2240_;
 wire _2241_;
 wire _2242_;
 wire _2243_;
 wire _2244_;
 wire _2245_;
 wire _2246_;
 wire _2247_;
 wire _2248_;
 wire _2249_;
 wire _2250_;
 wire _2251_;
 wire _2252_;
 wire _2253_;
 wire _2254_;
 wire _2255_;
 wire _2256_;
 wire _2257_;
 wire _2258_;
 wire _2259_;
 wire _2260_;
 wire _2261_;
 wire _2262_;
 wire _2263_;
 wire _2264_;
 wire _2265_;
 wire _2266_;
 wire _2267_;
 wire _2268_;
 wire _2269_;
 wire _2270_;
 wire _2271_;
 wire _2272_;
 wire _2273_;
 wire _2274_;
 wire _2275_;
 wire _2276_;
 wire _2277_;
 wire _2278_;
 wire _2279_;
 wire _2280_;
 wire _2281_;
 wire _2282_;
 wire _2283_;
 wire _2284_;
 wire _2285_;
 wire _2286_;
 wire _2287_;
 wire _2288_;
 wire _2289_;
 wire _2290_;
 wire _2291_;
 wire _2292_;
 wire _2293_;
 wire _2294_;
 wire _2295_;
 wire _2296_;
 wire _2297_;
 wire _2298_;
 wire _2299_;
 wire _2300_;
 wire _2301_;
 wire _2302_;
 wire _2303_;
 wire _2304_;
 wire _2305_;
 wire _2306_;
 wire _2307_;
 wire _2308_;
 wire _2309_;
 wire _2310_;
 wire _2311_;
 wire _2312_;
 wire _2313_;
 wire _2314_;
 wire _2315_;
 wire _2316_;
 wire _2317_;
 wire _2318_;
 wire _2319_;
 wire _2320_;
 wire _2321_;
 wire _2322_;
 wire _2323_;
 wire _2324_;
 wire _2325_;
 wire _2326_;
 wire _2327_;
 wire _2328_;
 wire _2329_;
 wire _2330_;
 wire _2331_;
 wire _2332_;
 wire _2333_;
 wire _2334_;
 wire _2335_;
 wire _2336_;
 wire _2337_;
 wire _2338_;
 wire _2339_;
 wire _2340_;
 wire _2341_;
 wire _2342_;
 wire _2343_;
 wire _2344_;
 wire _2345_;
 wire _2346_;
 wire _2347_;
 wire _2348_;
 wire _2349_;
 wire _2350_;
 wire _2351_;
 wire _2352_;
 wire _2353_;
 wire _2354_;
 wire _2355_;
 wire _2356_;
 wire _2357_;
 wire _2358_;
 wire _2359_;
 wire _2360_;
 wire _2361_;
 wire _2362_;
 wire _2363_;
 wire _2364_;
 wire _2365_;
 wire _2366_;
 wire _2367_;
 wire _2368_;
 wire _2369_;
 wire _2370_;
 wire _2371_;
 wire _2372_;
 wire _2373_;
 wire _2374_;
 wire _2375_;
 wire _2376_;
 wire _2377_;
 wire _2378_;
 wire _2379_;
 wire _2380_;
 wire _2381_;
 wire _2382_;
 wire _2383_;
 wire _2384_;
 wire _2385_;
 wire _2386_;
 wire _2387_;
 wire _2388_;
 wire _2389_;
 wire _2390_;
 wire _2391_;
 wire _2392_;
 wire _2393_;
 wire _2394_;
 wire _2395_;
 wire _2396_;
 wire _2397_;
 wire _2398_;
 wire _2399_;
 wire _2400_;
 wire _2401_;
 wire _2402_;
 wire _2403_;
 wire _2404_;
 wire _2405_;
 wire _2406_;
 wire _2407_;
 wire _2408_;
 wire _2409_;
 wire _2410_;
 wire _2411_;
 wire _2412_;
 wire _2413_;
 wire _2414_;
 wire _2415_;
 wire _2416_;
 wire _2417_;
 wire _2418_;
 wire _2419_;
 wire _2420_;
 wire _2421_;
 wire _2422_;
 wire _2423_;
 wire _2424_;
 wire _2425_;
 wire _2426_;
 wire _2427_;
 wire _2428_;
 wire _2429_;
 wire _2430_;
 wire _2431_;
 wire _2432_;
 wire _2433_;
 wire _2434_;
 wire _2435_;
 wire _2436_;
 wire _2437_;
 wire _2438_;
 wire _2439_;
 wire _2440_;
 wire _2441_;
 wire _2442_;
 wire _2443_;
 wire _2444_;
 wire _2445_;
 wire _2446_;
 wire _2447_;
 wire _2448_;
 wire _2449_;
 wire _2450_;
 wire _2451_;
 wire _2452_;
 wire _2453_;
 wire _2454_;
 wire _2455_;
 wire _2456_;
 wire _2457_;
 wire _2458_;
 wire _2459_;
 wire _2460_;
 wire _2461_;
 wire _2462_;
 wire _2463_;
 wire _2464_;
 wire _2465_;
 wire _2466_;
 wire _2467_;
 wire _2468_;
 wire _2469_;
 wire _2470_;
 wire _2471_;
 wire _2472_;
 wire _2473_;
 wire _2474_;
 wire _2475_;
 wire _2476_;
 wire _2477_;
 wire _2478_;
 wire _2479_;
 wire _2480_;
 wire _2481_;
 wire _2482_;
 wire _2483_;
 wire _2484_;
 wire _2485_;
 wire _2486_;
 wire _2487_;
 wire _2488_;
 wire _2489_;
 wire _2490_;
 wire _2491_;
 wire _2492_;
 wire _2493_;
 wire _2494_;
 wire _2495_;
 wire _2496_;
 wire _2497_;
 wire _2498_;
 wire _2499_;
 wire _2500_;
 wire _2501_;
 wire _2502_;
 wire _2503_;
 wire _2504_;
 wire _2505_;
 wire _2506_;
 wire _2507_;
 wire _2508_;
 wire _2509_;
 wire _2510_;
 wire _2511_;
 wire _2512_;
 wire _2513_;
 wire _2514_;
 wire _2515_;
 wire _2516_;
 wire _2517_;
 wire _2518_;
 wire _2519_;
 wire _2520_;
 wire _2521_;
 wire _2522_;
 wire _2523_;
 wire _2524_;
 wire _2525_;
 wire _2526_;
 wire _2527_;
 wire _2528_;
 wire _2529_;
 wire _2530_;
 wire _2531_;
 wire _2532_;
 wire _2533_;
 wire _2534_;
 wire _2535_;
 wire _2536_;
 wire _2537_;
 wire _2538_;
 wire _2539_;
 wire _2540_;
 wire _2541_;
 wire _2542_;
 wire _2543_;
 wire _2544_;
 wire _2545_;
 wire _2546_;
 wire _2547_;
 wire _2548_;
 wire _2549_;
 wire _2550_;
 wire _2551_;
 wire _2552_;
 wire _2553_;
 wire _2554_;
 wire _2555_;
 wire _2556_;
 wire _2557_;
 wire _2558_;
 wire _2559_;
 wire _2560_;
 wire _2561_;
 wire _2562_;
 wire _2563_;
 wire _2564_;
 wire _2565_;
 wire _2566_;
 wire _2567_;
 wire _2568_;
 wire _2569_;
 wire _2570_;
 wire _2571_;
 wire _2572_;
 wire _2573_;
 wire _2574_;
 wire _2575_;
 wire _2576_;
 wire _2577_;
 wire _2578_;
 wire _2579_;
 wire _2580_;
 wire _2581_;
 wire _2582_;
 wire _2583_;
 wire _2584_;
 wire _2585_;
 wire _2586_;
 wire _2587_;
 wire _2588_;
 wire _2589_;
 wire _2590_;
 wire _2591_;
 wire _2592_;
 wire _2593_;
 wire _2594_;
 wire _2595_;
 wire _2596_;
 wire _2597_;
 wire _2598_;
 wire _2599_;
 wire _2600_;
 wire _2601_;
 wire _2602_;
 wire _2603_;
 wire _2604_;
 wire _2605_;
 wire _2606_;
 wire _2607_;
 wire _2608_;
 wire _2609_;
 wire _2610_;
 wire _2611_;
 wire _2612_;
 wire _2613_;
 wire _2614_;
 wire _2615_;
 wire _2616_;
 wire _2617_;
 wire _2618_;
 wire _2619_;
 wire _2620_;
 wire _2621_;
 wire _2622_;
 wire _2623_;
 wire _2624_;
 wire _2625_;
 wire _2626_;
 wire _2627_;
 wire _2628_;
 wire _2629_;
 wire _2630_;
 wire _2631_;
 wire _2632_;
 wire _2633_;
 wire _2634_;
 wire _2635_;
 wire _2636_;
 wire _2637_;
 wire _2638_;
 wire _2639_;
 wire _2640_;
 wire _2641_;
 wire _2642_;
 wire _2643_;
 wire _2644_;
 wire _2645_;
 wire _2646_;
 wire _2647_;
 wire _2648_;
 wire _2649_;
 wire _2650_;
 wire _2651_;
 wire _2652_;
 wire _2653_;
 wire _2654_;
 wire _2655_;
 wire _2656_;
 wire _2657_;
 wire _2658_;
 wire _2659_;
 wire _2660_;
 wire _2661_;
 wire _2662_;
 wire _2663_;
 wire _2664_;
 wire _2665_;
 wire _2666_;
 wire _2667_;
 wire _2668_;
 wire _2669_;
 wire _2670_;
 wire _2671_;
 wire _2672_;
 wire _2673_;
 wire _2674_;
 wire _2675_;
 wire _2676_;
 wire _2677_;
 wire _2678_;
 wire _2679_;
 wire _2680_;
 wire _2681_;
 wire _2682_;
 wire _2683_;
 wire _2684_;
 wire _2685_;
 wire _2686_;
 wire _2687_;
 wire _2688_;
 wire _2689_;
 wire _2690_;
 wire _2691_;
 wire _2692_;
 wire _2693_;
 wire _2694_;
 wire _2695_;
 wire _2696_;
 wire _2697_;
 wire _2698_;
 wire _2699_;
 wire _2700_;
 wire _2701_;
 wire _2702_;
 wire _2703_;
 wire _2704_;
 wire _2705_;
 wire _2706_;
 wire _2707_;
 wire _2708_;
 wire _2709_;
 wire _2710_;
 wire _2711_;
 wire _2712_;
 wire _2713_;
 wire _2714_;
 wire _2715_;
 wire _2716_;
 wire _2717_;
 wire _2718_;
 wire _2719_;
 wire _2720_;
 wire _2721_;
 wire _2722_;
 wire _2723_;
 wire _2724_;
 wire _2725_;
 wire _2726_;
 wire _2727_;
 wire _2728_;
 wire _2729_;
 wire _2730_;
 wire _2731_;
 wire _2732_;
 wire _2733_;
 wire _2734_;
 wire _2735_;
 wire _2736_;
 wire _2737_;
 wire _2738_;
 wire _2739_;
 wire _2740_;
 wire _2741_;
 wire _2742_;
 wire _2743_;
 wire _2744_;
 wire _2745_;
 wire _2746_;
 wire _2747_;
 wire _2748_;
 wire _2749_;
 wire _2750_;
 wire _2751_;
 wire _2752_;
 wire _2753_;
 wire _2754_;
 wire _2755_;
 wire _2756_;
 wire _2757_;
 wire _2758_;
 wire _2759_;
 wire _2760_;
 wire _2761_;
 wire _2762_;
 wire _2763_;
 wire _2764_;
 wire _2765_;
 wire _2766_;
 wire _2767_;
 wire _2768_;
 wire _2769_;
 wire _2770_;
 wire _2771_;
 wire _2772_;
 wire _2773_;
 wire _2774_;
 wire _2775_;
 wire _2776_;
 wire _2777_;
 wire _2778_;
 wire _2779_;
 wire _2780_;
 wire _2781_;
 wire _2782_;
 wire _2783_;
 wire _2784_;
 wire _2785_;
 wire _2786_;
 wire _2787_;
 wire _2788_;
 wire _2789_;
 wire _2790_;
 wire _2791_;
 wire _2792_;
 wire _2793_;
 wire _2794_;
 wire _2795_;
 wire _2796_;
 wire _2797_;
 wire _2798_;
 wire _2799_;
 wire _2800_;
 wire _2801_;
 wire _2802_;
 wire _2803_;
 wire _2804_;
 wire _2805_;
 wire _2806_;
 wire _2807_;
 wire _2808_;
 wire _2809_;
 wire _2810_;
 wire _2811_;
 wire _2812_;
 wire _2813_;
 wire _2814_;
 wire _2815_;
 wire _2816_;
 wire _2817_;
 wire _2818_;
 wire _2819_;
 wire _2820_;
 wire _2821_;
 wire _2822_;
 wire _2823_;
 wire _2824_;
 wire _2825_;
 wire _2826_;
 wire _2827_;
 wire _2828_;
 wire _2829_;
 wire _2830_;
 wire _2831_;
 wire _2832_;
 wire _2833_;
 wire _2834_;
 wire _2835_;
 wire _2836_;
 wire _2837_;
 wire _2838_;
 wire _2839_;
 wire _2840_;
 wire _2841_;
 wire _2842_;
 wire _2843_;
 wire _2844_;
 wire _2845_;
 wire _2846_;
 wire _2847_;
 wire _2848_;
 wire _2849_;
 wire _2850_;
 wire _2851_;
 wire _2852_;
 wire _2853_;
 wire _2854_;
 wire _2855_;
 wire _2856_;
 wire _2857_;
 wire _2858_;
 wire _2859_;
 wire _2860_;
 wire _2861_;
 wire _2862_;
 wire _2863_;
 wire _2864_;
 wire _2865_;
 wire _2866_;
 wire _2867_;
 wire _2868_;
 wire _2869_;
 wire _2870_;
 wire _2871_;
 wire _2872_;
 wire _2873_;
 wire _2874_;
 wire _2875_;
 wire _2876_;
 wire _2877_;
 wire _2878_;
 wire _2879_;
 wire _2880_;
 wire _2881_;
 wire _2882_;
 wire _2883_;
 wire _2884_;
 wire _2885_;
 wire _2886_;
 wire _2887_;
 wire _2888_;
 wire _2889_;
 wire _2890_;
 wire _2891_;
 wire _2892_;
 wire _2893_;
 wire _2894_;
 wire _2895_;
 wire _2896_;
 wire _2897_;
 wire _2898_;
 wire _2899_;
 wire _2900_;
 wire _2901_;
 wire _2902_;
 wire _2903_;
 wire _2904_;
 wire _2905_;
 wire _2906_;
 wire _2907_;
 wire _2908_;
 wire _2909_;
 wire _2910_;
 wire _2911_;
 wire _2912_;
 wire _2913_;
 wire _2914_;
 wire _2915_;
 wire _2916_;
 wire _2917_;
 wire _2918_;
 wire _2919_;
 wire _2920_;
 wire _2921_;
 wire _2922_;
 wire _2923_;
 wire _2924_;
 wire _2925_;
 wire _2926_;
 wire _2927_;
 wire _2928_;
 wire _2929_;
 wire _2930_;
 wire _2931_;
 wire _2932_;
 wire _2933_;
 wire _2934_;
 wire _2935_;
 wire _2936_;
 wire _2937_;
 wire _2938_;
 wire _2939_;
 wire _2940_;
 wire _2941_;
 wire _2942_;
 wire _2943_;
 wire _2944_;
 wire _2945_;
 wire _2946_;
 wire _2947_;
 wire _2948_;
 wire _2949_;
 wire _2950_;
 wire _2951_;
 wire _2952_;
 wire _2953_;
 wire _2954_;
 wire _2955_;
 wire _2956_;
 wire _2957_;
 wire _2958_;
 wire _2959_;
 wire _2960_;
 wire _2961_;
 wire _2962_;
 wire _2963_;
 wire _2964_;
 wire _2965_;
 wire _2966_;
 wire _2967_;
 wire _2968_;
 wire _2969_;
 wire _2970_;
 wire _2971_;
 wire _2972_;
 wire _2973_;
 wire _2974_;
 wire _2975_;
 wire _2976_;
 wire _2977_;
 wire _2978_;
 wire _2979_;
 wire _2980_;
 wire _2981_;
 wire _2982_;
 wire _2983_;
 wire _2984_;
 wire _2985_;
 wire _2986_;
 wire _2987_;
 wire _2988_;
 wire _2989_;
 wire _2990_;
 wire _2991_;
 wire _2992_;
 wire _2993_;
 wire _2994_;
 wire _2995_;
 wire _2996_;
 wire _2997_;
 wire _2998_;
 wire _2999_;
 wire _3000_;
 wire _3001_;
 wire _3002_;
 wire _3003_;
 wire _3004_;
 wire _3005_;
 wire _3006_;
 wire _3007_;
 wire _3008_;
 wire _3009_;
 wire _3010_;
 wire _3011_;
 wire _3012_;
 wire _3013_;
 wire _3014_;
 wire _3015_;
 wire _3016_;
 wire _3017_;
 wire _3018_;
 wire _3019_;
 wire _3020_;
 wire _3021_;
 wire _3022_;
 wire _3023_;
 wire _3024_;
 wire _3025_;
 wire _3026_;
 wire _3027_;
 wire _3028_;
 wire _3029_;
 wire _3030_;
 wire _3031_;
 wire _3032_;
 wire _3033_;
 wire _3034_;
 wire _3035_;
 wire _3036_;
 wire _3037_;
 wire _3038_;
 wire _3039_;
 wire _3040_;
 wire _3041_;
 wire _3042_;
 wire _3043_;
 wire _3044_;
 wire _3045_;
 wire _3046_;
 wire _3047_;
 wire _3048_;
 wire _3049_;
 wire _3050_;
 wire _3051_;
 wire _3052_;
 wire _3053_;
 wire _3054_;
 wire _3055_;
 wire _3056_;
 wire _3057_;
 wire _3058_;
 wire _3059_;
 wire _3060_;
 wire _3061_;
 wire _3062_;
 wire _3063_;
 wire _3064_;
 wire _3065_;
 wire _3066_;
 wire _3067_;
 wire _3068_;
 wire _3069_;
 wire _3070_;
 wire _3071_;
 wire _3072_;
 wire _3073_;
 wire _3074_;
 wire _3075_;
 wire _3076_;
 wire _3077_;
 wire _3078_;
 wire _3079_;
 wire _3080_;
 wire _3081_;
 wire _3082_;
 wire _3083_;
 wire _3084_;
 wire _3085_;
 wire _3086_;
 wire _3087_;
 wire _3088_;
 wire _3089_;
 wire _3090_;
 wire _3091_;
 wire _3092_;
 wire _3093_;
 wire _3094_;
 wire _3095_;
 wire _3096_;
 wire _3097_;
 wire _3098_;
 wire _3099_;
 wire _3100_;
 wire _3101_;
 wire _3102_;
 wire _3103_;
 wire _3104_;
 wire _3105_;
 wire _3106_;
 wire _3107_;
 wire _3108_;
 wire _3109_;
 wire _3110_;
 wire _3111_;
 wire _3112_;
 wire _3113_;
 wire _3114_;
 wire _3115_;
 wire _3116_;
 wire _3117_;
 wire _3118_;
 wire _3119_;
 wire _3120_;
 wire _3121_;
 wire _3122_;
 wire _3123_;
 wire _3124_;
 wire _3125_;
 wire _3126_;
 wire _3127_;
 wire _3128_;
 wire _3129_;
 wire _3130_;
 wire _3131_;
 wire _3132_;
 wire _3133_;
 wire _3134_;
 wire _3135_;
 wire _3136_;
 wire _3137_;
 wire _3138_;
 wire _3139_;
 wire _3140_;
 wire _3141_;
 wire _3142_;
 wire _3143_;
 wire _3144_;
 wire _3145_;
 wire _3146_;
 wire _3147_;
 wire _3148_;
 wire _3149_;
 wire _3150_;
 wire _3151_;
 wire _3152_;
 wire _3153_;
 wire _3154_;
 wire _3155_;
 wire _3156_;
 wire _3157_;
 wire _3158_;
 wire _3159_;
 wire _3160_;
 wire _3161_;
 wire _3162_;
 wire _3163_;
 wire _3164_;
 wire _3165_;
 wire _3166_;
 wire _3167_;
 wire _3168_;
 wire _3169_;
 wire _3170_;
 wire _3171_;
 wire _3172_;
 wire _3173_;
 wire _3174_;
 wire _3175_;
 wire _3176_;
 wire _3177_;
 wire _3178_;
 wire _3179_;
 wire _3180_;
 wire _3181_;
 wire _3182_;
 wire _3183_;
 wire _3184_;
 wire _3185_;
 wire _3186_;
 wire _3187_;
 wire _3188_;
 wire _3189_;
 wire _3190_;
 wire _3191_;
 wire _3192_;
 wire _3193_;
 wire _3194_;
 wire _3195_;
 wire _3196_;
 wire _3197_;
 wire _3198_;
 wire _3199_;
 wire _3200_;
 wire _3201_;
 wire _3202_;
 wire _3203_;
 wire _3204_;
 wire _3205_;
 wire _3206_;
 wire _3207_;
 wire _3208_;
 wire _3209_;
 wire _3210_;
 wire _3211_;
 wire _3212_;
 wire _3213_;
 wire _3214_;
 wire _3215_;
 wire _3216_;
 wire _3217_;
 wire _3218_;
 wire _3219_;
 wire _3220_;
 wire _3221_;
 wire _3222_;
 wire _3223_;
 wire _3224_;
 wire _3225_;
 wire _3226_;
 wire _3227_;
 wire _3228_;
 wire _3229_;
 wire _3230_;
 wire _3231_;
 wire _3232_;
 wire _3233_;
 wire _3234_;
 wire _3235_;
 wire _3236_;
 wire _3237_;
 wire _3238_;
 wire _3239_;
 wire _3240_;
 wire _3241_;
 wire _3242_;
 wire _3243_;
 wire _3244_;
 wire _3245_;
 wire _3246_;
 wire _3247_;
 wire _3248_;
 wire _3249_;
 wire _3250_;
 wire _3251_;
 wire _3252_;
 wire _3253_;
 wire _3254_;
 wire _3255_;
 wire _3256_;
 wire _3257_;
 wire _3258_;
 wire _3259_;
 wire _3260_;
 wire _3261_;
 wire _3262_;
 wire _3263_;
 wire _3264_;
 wire _3265_;
 wire _3266_;
 wire _3267_;
 wire _3268_;
 wire _3269_;
 wire _3270_;
 wire _3271_;
 wire _3272_;
 wire _3273_;
 wire _3274_;
 wire _3275_;
 wire _3276_;
 wire _3277_;
 wire _3278_;
 wire _3279_;
 wire _3280_;
 wire _3281_;
 wire _3282_;
 wire _3283_;
 wire _3284_;
 wire _3285_;
 wire _3286_;
 wire _3287_;
 wire _3288_;
 wire _3289_;
 wire _3290_;
 wire _3291_;
 wire _3292_;
 wire _3293_;
 wire _3294_;
 wire _3295_;
 wire _3296_;
 wire _3297_;
 wire _3298_;
 wire _3299_;
 wire _3300_;
 wire _3301_;
 wire _3302_;
 wire _3303_;
 wire _3304_;
 wire _3305_;
 wire _3306_;
 wire _3307_;
 wire _3308_;
 wire _3309_;
 wire _3310_;
 wire _3311_;
 wire _3312_;
 wire _3313_;
 wire _3314_;
 wire _3315_;
 wire _3316_;
 wire _3317_;
 wire _3318_;
 wire _3319_;
 wire _3320_;
 wire _3321_;
 wire _3322_;
 wire _3323_;
 wire _3324_;
 wire _3325_;
 wire _3326_;
 wire _3327_;
 wire _3328_;
 wire _3329_;
 wire _3330_;
 wire _3331_;
 wire _3332_;
 wire _3333_;
 wire _3334_;
 wire _3335_;
 wire _3336_;
 wire _3337_;
 wire _3338_;
 wire _3339_;
 wire _3340_;
 wire _3341_;
 wire _3342_;
 wire _3343_;
 wire _3344_;
 wire _3345_;
 wire _3346_;
 wire _3347_;
 wire _3348_;
 wire _3349_;
 wire _3350_;
 wire _3351_;
 wire _3352_;
 wire _3353_;
 wire _3354_;
 wire _3355_;
 wire _3356_;
 wire _3357_;
 wire _3358_;
 wire _3359_;
 wire \core_1.de_jmp_pred ;
 wire \core_1.dec_alu_carry_en ;
 wire \core_1.dec_alu_flags_ie ;
 wire \core_1.dec_jump_cond_code[0] ;
 wire \core_1.dec_jump_cond_code[1] ;
 wire \core_1.dec_jump_cond_code[2] ;
 wire \core_1.dec_jump_cond_code[3] ;
 wire \core_1.dec_jump_cond_code[4] ;
 wire \core_1.dec_l_reg_sel[0] ;
 wire \core_1.dec_l_reg_sel[1] ;
 wire \core_1.dec_l_reg_sel[2] ;
 wire \core_1.dec_mem_access ;
 wire \core_1.dec_mem_long ;
 wire \core_1.dec_mem_we ;
 wire \core_1.dec_mem_width ;
 wire \core_1.dec_pc_inc ;
 wire \core_1.dec_r_bus_imm ;
 wire \core_1.dec_r_reg_sel[0] ;
 wire \core_1.dec_r_reg_sel[1] ;
 wire \core_1.dec_r_reg_sel[2] ;
 wire \core_1.dec_rf_ie[0] ;
 wire \core_1.dec_rf_ie[1] ;
 wire \core_1.dec_rf_ie[2] ;
 wire \core_1.dec_rf_ie[3] ;
 wire \core_1.dec_rf_ie[4] ;
 wire \core_1.dec_rf_ie[5] ;
 wire \core_1.dec_rf_ie[6] ;
 wire \core_1.dec_rf_ie[7] ;
 wire \core_1.dec_sreg_irt ;
 wire \core_1.dec_sreg_jal_over ;
 wire \core_1.dec_sreg_load ;
 wire \core_1.dec_sreg_store ;
 wire \core_1.dec_sys ;
 wire \core_1.dec_used_operands[0] ;
 wire \core_1.dec_used_operands[1] ;
 wire \core_1.decode.i_flush ;
 wire \core_1.decode.i_imm_pass[0] ;
 wire \core_1.decode.i_imm_pass[10] ;
 wire \core_1.decode.i_imm_pass[11] ;
 wire \core_1.decode.i_imm_pass[12] ;
 wire \core_1.decode.i_imm_pass[13] ;
 wire \core_1.decode.i_imm_pass[14] ;
 wire \core_1.decode.i_imm_pass[15] ;
 wire \core_1.decode.i_imm_pass[1] ;
 wire \core_1.decode.i_imm_pass[2] ;
 wire \core_1.decode.i_imm_pass[3] ;
 wire \core_1.decode.i_imm_pass[4] ;
 wire \core_1.decode.i_imm_pass[5] ;
 wire \core_1.decode.i_imm_pass[6] ;
 wire \core_1.decode.i_imm_pass[7] ;
 wire \core_1.decode.i_imm_pass[8] ;
 wire \core_1.decode.i_imm_pass[9] ;
 wire \core_1.decode.i_instr_l[0] ;
 wire \core_1.decode.i_instr_l[10] ;
 wire \core_1.decode.i_instr_l[11] ;
 wire \core_1.decode.i_instr_l[12] ;
 wire \core_1.decode.i_instr_l[13] ;
 wire \core_1.decode.i_instr_l[14] ;
 wire \core_1.decode.i_instr_l[15] ;
 wire \core_1.decode.i_instr_l[1] ;
 wire \core_1.decode.i_instr_l[2] ;
 wire \core_1.decode.i_instr_l[3] ;
 wire \core_1.decode.i_instr_l[4] ;
 wire \core_1.decode.i_instr_l[5] ;
 wire \core_1.decode.i_instr_l[6] ;
 wire \core_1.decode.i_instr_l[7] ;
 wire \core_1.decode.i_instr_l[8] ;
 wire \core_1.decode.i_instr_l[9] ;
 wire \core_1.decode.i_jmp_pred_pass ;
 wire \core_1.decode.i_submit ;
 wire \core_1.decode.input_valid ;
 wire \core_1.decode.o_submit ;
 wire \core_1.decode.oc_alu_mode[11] ;
 wire \core_1.decode.oc_alu_mode[12] ;
 wire \core_1.decode.oc_alu_mode[13] ;
 wire \core_1.decode.oc_alu_mode[1] ;
 wire \core_1.decode.oc_alu_mode[2] ;
 wire \core_1.decode.oc_alu_mode[3] ;
 wire \core_1.decode.oc_alu_mode[4] ;
 wire \core_1.decode.oc_alu_mode[6] ;
 wire \core_1.decode.oc_alu_mode[7] ;
 wire \core_1.decode.oc_alu_mode[9] ;
 wire \core_1.ew_addr[0] ;
 wire \core_1.ew_addr_high[0] ;
 wire \core_1.ew_data[0] ;
 wire \core_1.ew_data[10] ;
 wire \core_1.ew_data[11] ;
 wire \core_1.ew_data[12] ;
 wire \core_1.ew_data[13] ;
 wire \core_1.ew_data[14] ;
 wire \core_1.ew_data[15] ;
 wire \core_1.ew_data[1] ;
 wire \core_1.ew_data[2] ;
 wire \core_1.ew_data[3] ;
 wire \core_1.ew_data[4] ;
 wire \core_1.ew_data[5] ;
 wire \core_1.ew_data[6] ;
 wire \core_1.ew_data[7] ;
 wire \core_1.ew_data[8] ;
 wire \core_1.ew_data[9] ;
 wire \core_1.ew_mem_access ;
 wire \core_1.ew_mem_width ;
 wire \core_1.ew_reg_ie[0] ;
 wire \core_1.ew_reg_ie[1] ;
 wire \core_1.ew_reg_ie[2] ;
 wire \core_1.ew_reg_ie[3] ;
 wire \core_1.ew_reg_ie[4] ;
 wire \core_1.ew_reg_ie[5] ;
 wire \core_1.ew_reg_ie[6] ;
 wire \core_1.ew_reg_ie[7] ;
 wire \core_1.ew_submit ;
 wire \core_1.execute.alu_flag_reg.o_d[0] ;
 wire \core_1.execute.alu_flag_reg.o_d[1] ;
 wire \core_1.execute.alu_flag_reg.o_d[2] ;
 wire \core_1.execute.alu_flag_reg.o_d[3] ;
 wire \core_1.execute.alu_flag_reg.o_d[4] ;
 wire \core_1.execute.alu_mul_div.cbit[0] ;
 wire \core_1.execute.alu_mul_div.cbit[1] ;
 wire \core_1.execute.alu_mul_div.cbit[2] ;
 wire \core_1.execute.alu_mul_div.cbit[3] ;
 wire \core_1.execute.alu_mul_div.comp ;
 wire \core_1.execute.alu_mul_div.div_cur[0] ;
 wire \core_1.execute.alu_mul_div.div_cur[10] ;
 wire \core_1.execute.alu_mul_div.div_cur[11] ;
 wire \core_1.execute.alu_mul_div.div_cur[12] ;
 wire \core_1.execute.alu_mul_div.div_cur[13] ;
 wire \core_1.execute.alu_mul_div.div_cur[14] ;
 wire \core_1.execute.alu_mul_div.div_cur[15] ;
 wire \core_1.execute.alu_mul_div.div_cur[1] ;
 wire \core_1.execute.alu_mul_div.div_cur[2] ;
 wire \core_1.execute.alu_mul_div.div_cur[3] ;
 wire \core_1.execute.alu_mul_div.div_cur[4] ;
 wire \core_1.execute.alu_mul_div.div_cur[5] ;
 wire \core_1.execute.alu_mul_div.div_cur[6] ;
 wire \core_1.execute.alu_mul_div.div_cur[7] ;
 wire \core_1.execute.alu_mul_div.div_cur[8] ;
 wire \core_1.execute.alu_mul_div.div_cur[9] ;
 wire \core_1.execute.alu_mul_div.div_res[0] ;
 wire \core_1.execute.alu_mul_div.div_res[10] ;
 wire \core_1.execute.alu_mul_div.div_res[11] ;
 wire \core_1.execute.alu_mul_div.div_res[12] ;
 wire \core_1.execute.alu_mul_div.div_res[13] ;
 wire \core_1.execute.alu_mul_div.div_res[14] ;
 wire \core_1.execute.alu_mul_div.div_res[15] ;
 wire \core_1.execute.alu_mul_div.div_res[1] ;
 wire \core_1.execute.alu_mul_div.div_res[2] ;
 wire \core_1.execute.alu_mul_div.div_res[3] ;
 wire \core_1.execute.alu_mul_div.div_res[4] ;
 wire \core_1.execute.alu_mul_div.div_res[5] ;
 wire \core_1.execute.alu_mul_div.div_res[6] ;
 wire \core_1.execute.alu_mul_div.div_res[7] ;
 wire \core_1.execute.alu_mul_div.div_res[8] ;
 wire \core_1.execute.alu_mul_div.div_res[9] ;
 wire \core_1.execute.alu_mul_div.i_div ;
 wire \core_1.execute.alu_mul_div.i_mod ;
 wire \core_1.execute.alu_mul_div.i_mul ;
 wire \core_1.execute.alu_mul_div.mul_res[0] ;
 wire \core_1.execute.alu_mul_div.mul_res[10] ;
 wire \core_1.execute.alu_mul_div.mul_res[11] ;
 wire \core_1.execute.alu_mul_div.mul_res[12] ;
 wire \core_1.execute.alu_mul_div.mul_res[13] ;
 wire \core_1.execute.alu_mul_div.mul_res[14] ;
 wire \core_1.execute.alu_mul_div.mul_res[15] ;
 wire \core_1.execute.alu_mul_div.mul_res[1] ;
 wire \core_1.execute.alu_mul_div.mul_res[2] ;
 wire \core_1.execute.alu_mul_div.mul_res[3] ;
 wire \core_1.execute.alu_mul_div.mul_res[4] ;
 wire \core_1.execute.alu_mul_div.mul_res[5] ;
 wire \core_1.execute.alu_mul_div.mul_res[6] ;
 wire \core_1.execute.alu_mul_div.mul_res[7] ;
 wire \core_1.execute.alu_mul_div.mul_res[8] ;
 wire \core_1.execute.alu_mul_div.mul_res[9] ;
 wire \core_1.execute.hold_valid ;
 wire \core_1.execute.irq_en ;
 wire \core_1.execute.mem_stage_pc[0] ;
 wire \core_1.execute.mem_stage_pc[10] ;
 wire \core_1.execute.mem_stage_pc[11] ;
 wire \core_1.execute.mem_stage_pc[12] ;
 wire \core_1.execute.mem_stage_pc[13] ;
 wire \core_1.execute.mem_stage_pc[14] ;
 wire \core_1.execute.mem_stage_pc[15] ;
 wire \core_1.execute.mem_stage_pc[1] ;
 wire \core_1.execute.mem_stage_pc[2] ;
 wire \core_1.execute.mem_stage_pc[3] ;
 wire \core_1.execute.mem_stage_pc[4] ;
 wire \core_1.execute.mem_stage_pc[5] ;
 wire \core_1.execute.mem_stage_pc[6] ;
 wire \core_1.execute.mem_stage_pc[7] ;
 wire \core_1.execute.mem_stage_pc[8] ;
 wire \core_1.execute.mem_stage_pc[9] ;
 wire \core_1.execute.next_ready_delayed ;
 wire \core_1.execute.pc_high_buff_out[0] ;
 wire \core_1.execute.pc_high_buff_out[1] ;
 wire \core_1.execute.pc_high_buff_out[2] ;
 wire \core_1.execute.pc_high_buff_out[3] ;
 wire \core_1.execute.pc_high_buff_out[4] ;
 wire \core_1.execute.pc_high_buff_out[5] ;
 wire \core_1.execute.pc_high_buff_out[6] ;
 wire \core_1.execute.pc_high_buff_out[7] ;
 wire \core_1.execute.pc_high_out[0] ;
 wire \core_1.execute.pc_high_out[1] ;
 wire \core_1.execute.pc_high_out[2] ;
 wire \core_1.execute.pc_high_out[3] ;
 wire \core_1.execute.pc_high_out[4] ;
 wire \core_1.execute.pc_high_out[5] ;
 wire \core_1.execute.pc_high_out[6] ;
 wire \core_1.execute.pc_high_out[7] ;
 wire \core_1.execute.prev_pc_high[0] ;
 wire \core_1.execute.prev_pc_high[1] ;
 wire \core_1.execute.prev_pc_high[2] ;
 wire \core_1.execute.prev_pc_high[3] ;
 wire \core_1.execute.prev_pc_high[4] ;
 wire \core_1.execute.prev_pc_high[5] ;
 wire \core_1.execute.prev_pc_high[6] ;
 wire \core_1.execute.prev_pc_high[7] ;
 wire \core_1.execute.prev_sys ;
 wire \core_1.execute.rf.reg_outputs[1][0] ;
 wire \core_1.execute.rf.reg_outputs[1][10] ;
 wire \core_1.execute.rf.reg_outputs[1][11] ;
 wire \core_1.execute.rf.reg_outputs[1][12] ;
 wire \core_1.execute.rf.reg_outputs[1][13] ;
 wire \core_1.execute.rf.reg_outputs[1][14] ;
 wire \core_1.execute.rf.reg_outputs[1][15] ;
 wire \core_1.execute.rf.reg_outputs[1][1] ;
 wire \core_1.execute.rf.reg_outputs[1][2] ;
 wire \core_1.execute.rf.reg_outputs[1][3] ;
 wire \core_1.execute.rf.reg_outputs[1][4] ;
 wire \core_1.execute.rf.reg_outputs[1][5] ;
 wire \core_1.execute.rf.reg_outputs[1][6] ;
 wire \core_1.execute.rf.reg_outputs[1][7] ;
 wire \core_1.execute.rf.reg_outputs[1][8] ;
 wire \core_1.execute.rf.reg_outputs[1][9] ;
 wire \core_1.execute.rf.reg_outputs[2][0] ;
 wire \core_1.execute.rf.reg_outputs[2][10] ;
 wire \core_1.execute.rf.reg_outputs[2][11] ;
 wire \core_1.execute.rf.reg_outputs[2][12] ;
 wire \core_1.execute.rf.reg_outputs[2][13] ;
 wire \core_1.execute.rf.reg_outputs[2][14] ;
 wire \core_1.execute.rf.reg_outputs[2][15] ;
 wire \core_1.execute.rf.reg_outputs[2][1] ;
 wire \core_1.execute.rf.reg_outputs[2][2] ;
 wire \core_1.execute.rf.reg_outputs[2][3] ;
 wire \core_1.execute.rf.reg_outputs[2][4] ;
 wire \core_1.execute.rf.reg_outputs[2][5] ;
 wire \core_1.execute.rf.reg_outputs[2][6] ;
 wire \core_1.execute.rf.reg_outputs[2][7] ;
 wire \core_1.execute.rf.reg_outputs[2][8] ;
 wire \core_1.execute.rf.reg_outputs[2][9] ;
 wire \core_1.execute.rf.reg_outputs[3][0] ;
 wire \core_1.execute.rf.reg_outputs[3][10] ;
 wire \core_1.execute.rf.reg_outputs[3][11] ;
 wire \core_1.execute.rf.reg_outputs[3][12] ;
 wire \core_1.execute.rf.reg_outputs[3][13] ;
 wire \core_1.execute.rf.reg_outputs[3][14] ;
 wire \core_1.execute.rf.reg_outputs[3][15] ;
 wire \core_1.execute.rf.reg_outputs[3][1] ;
 wire \core_1.execute.rf.reg_outputs[3][2] ;
 wire \core_1.execute.rf.reg_outputs[3][3] ;
 wire \core_1.execute.rf.reg_outputs[3][4] ;
 wire \core_1.execute.rf.reg_outputs[3][5] ;
 wire \core_1.execute.rf.reg_outputs[3][6] ;
 wire \core_1.execute.rf.reg_outputs[3][7] ;
 wire \core_1.execute.rf.reg_outputs[3][8] ;
 wire \core_1.execute.rf.reg_outputs[3][9] ;
 wire \core_1.execute.rf.reg_outputs[4][0] ;
 wire \core_1.execute.rf.reg_outputs[4][10] ;
 wire \core_1.execute.rf.reg_outputs[4][11] ;
 wire \core_1.execute.rf.reg_outputs[4][12] ;
 wire \core_1.execute.rf.reg_outputs[4][13] ;
 wire \core_1.execute.rf.reg_outputs[4][14] ;
 wire \core_1.execute.rf.reg_outputs[4][15] ;
 wire \core_1.execute.rf.reg_outputs[4][1] ;
 wire \core_1.execute.rf.reg_outputs[4][2] ;
 wire \core_1.execute.rf.reg_outputs[4][3] ;
 wire \core_1.execute.rf.reg_outputs[4][4] ;
 wire \core_1.execute.rf.reg_outputs[4][5] ;
 wire \core_1.execute.rf.reg_outputs[4][6] ;
 wire \core_1.execute.rf.reg_outputs[4][7] ;
 wire \core_1.execute.rf.reg_outputs[4][8] ;
 wire \core_1.execute.rf.reg_outputs[4][9] ;
 wire \core_1.execute.rf.reg_outputs[5][0] ;
 wire \core_1.execute.rf.reg_outputs[5][10] ;
 wire \core_1.execute.rf.reg_outputs[5][11] ;
 wire \core_1.execute.rf.reg_outputs[5][12] ;
 wire \core_1.execute.rf.reg_outputs[5][13] ;
 wire \core_1.execute.rf.reg_outputs[5][14] ;
 wire \core_1.execute.rf.reg_outputs[5][15] ;
 wire \core_1.execute.rf.reg_outputs[5][1] ;
 wire \core_1.execute.rf.reg_outputs[5][2] ;
 wire \core_1.execute.rf.reg_outputs[5][3] ;
 wire \core_1.execute.rf.reg_outputs[5][4] ;
 wire \core_1.execute.rf.reg_outputs[5][5] ;
 wire \core_1.execute.rf.reg_outputs[5][6] ;
 wire \core_1.execute.rf.reg_outputs[5][7] ;
 wire \core_1.execute.rf.reg_outputs[5][8] ;
 wire \core_1.execute.rf.reg_outputs[5][9] ;
 wire \core_1.execute.rf.reg_outputs[6][0] ;
 wire \core_1.execute.rf.reg_outputs[6][10] ;
 wire \core_1.execute.rf.reg_outputs[6][11] ;
 wire \core_1.execute.rf.reg_outputs[6][12] ;
 wire \core_1.execute.rf.reg_outputs[6][13] ;
 wire \core_1.execute.rf.reg_outputs[6][14] ;
 wire \core_1.execute.rf.reg_outputs[6][15] ;
 wire \core_1.execute.rf.reg_outputs[6][1] ;
 wire \core_1.execute.rf.reg_outputs[6][2] ;
 wire \core_1.execute.rf.reg_outputs[6][3] ;
 wire \core_1.execute.rf.reg_outputs[6][4] ;
 wire \core_1.execute.rf.reg_outputs[6][5] ;
 wire \core_1.execute.rf.reg_outputs[6][6] ;
 wire \core_1.execute.rf.reg_outputs[6][7] ;
 wire \core_1.execute.rf.reg_outputs[6][8] ;
 wire \core_1.execute.rf.reg_outputs[6][9] ;
 wire \core_1.execute.rf.reg_outputs[7][0] ;
 wire \core_1.execute.rf.reg_outputs[7][10] ;
 wire \core_1.execute.rf.reg_outputs[7][11] ;
 wire \core_1.execute.rf.reg_outputs[7][12] ;
 wire \core_1.execute.rf.reg_outputs[7][13] ;
 wire \core_1.execute.rf.reg_outputs[7][14] ;
 wire \core_1.execute.rf.reg_outputs[7][15] ;
 wire \core_1.execute.rf.reg_outputs[7][1] ;
 wire \core_1.execute.rf.reg_outputs[7][2] ;
 wire \core_1.execute.rf.reg_outputs[7][3] ;
 wire \core_1.execute.rf.reg_outputs[7][4] ;
 wire \core_1.execute.rf.reg_outputs[7][5] ;
 wire \core_1.execute.rf.reg_outputs[7][6] ;
 wire \core_1.execute.rf.reg_outputs[7][7] ;
 wire \core_1.execute.rf.reg_outputs[7][8] ;
 wire \core_1.execute.rf.reg_outputs[7][9] ;
 wire \core_1.execute.sreg_data_page ;
 wire \core_1.execute.sreg_irq_flags.i_d[2] ;
 wire \core_1.execute.sreg_irq_flags.o_d[0] ;
 wire \core_1.execute.sreg_irq_flags.o_d[1] ;
 wire \core_1.execute.sreg_irq_flags.o_d[2] ;
 wire \core_1.execute.sreg_irq_flags.o_d[3] ;
 wire \core_1.execute.sreg_irq_flags.o_d[4] ;
 wire \core_1.execute.sreg_irq_pc.o_d[0] ;
 wire \core_1.execute.sreg_irq_pc.o_d[10] ;
 wire \core_1.execute.sreg_irq_pc.o_d[11] ;
 wire \core_1.execute.sreg_irq_pc.o_d[12] ;
 wire \core_1.execute.sreg_irq_pc.o_d[13] ;
 wire \core_1.execute.sreg_irq_pc.o_d[14] ;
 wire \core_1.execute.sreg_irq_pc.o_d[15] ;
 wire \core_1.execute.sreg_irq_pc.o_d[1] ;
 wire \core_1.execute.sreg_irq_pc.o_d[2] ;
 wire \core_1.execute.sreg_irq_pc.o_d[3] ;
 wire \core_1.execute.sreg_irq_pc.o_d[4] ;
 wire \core_1.execute.sreg_irq_pc.o_d[5] ;
 wire \core_1.execute.sreg_irq_pc.o_d[6] ;
 wire \core_1.execute.sreg_irq_pc.o_d[7] ;
 wire \core_1.execute.sreg_irq_pc.o_d[8] ;
 wire \core_1.execute.sreg_irq_pc.o_d[9] ;
 wire \core_1.execute.sreg_jtr_buff.o_d[0] ;
 wire \core_1.execute.sreg_jtr_buff.o_d[1] ;
 wire \core_1.execute.sreg_jtr_buff.o_d[2] ;
 wire \core_1.execute.sreg_long_ptr_en ;
 wire \core_1.execute.sreg_priv_control.o_d[0] ;
 wire \core_1.execute.sreg_priv_control.o_d[10] ;
 wire \core_1.execute.sreg_priv_control.o_d[11] ;
 wire \core_1.execute.sreg_priv_control.o_d[12] ;
 wire \core_1.execute.sreg_priv_control.o_d[13] ;
 wire \core_1.execute.sreg_priv_control.o_d[14] ;
 wire \core_1.execute.sreg_priv_control.o_d[15] ;
 wire \core_1.execute.sreg_priv_control.o_d[4] ;
 wire \core_1.execute.sreg_priv_control.o_d[5] ;
 wire \core_1.execute.sreg_priv_control.o_d[6] ;
 wire \core_1.execute.sreg_priv_control.o_d[7] ;
 wire \core_1.execute.sreg_priv_control.o_d[8] ;
 wire \core_1.execute.sreg_priv_control.o_d[9] ;
 wire \core_1.execute.sreg_scratch.o_d[0] ;
 wire \core_1.execute.sreg_scratch.o_d[10] ;
 wire \core_1.execute.sreg_scratch.o_d[11] ;
 wire \core_1.execute.sreg_scratch.o_d[12] ;
 wire \core_1.execute.sreg_scratch.o_d[13] ;
 wire \core_1.execute.sreg_scratch.o_d[14] ;
 wire \core_1.execute.sreg_scratch.o_d[15] ;
 wire \core_1.execute.sreg_scratch.o_d[1] ;
 wire \core_1.execute.sreg_scratch.o_d[2] ;
 wire \core_1.execute.sreg_scratch.o_d[3] ;
 wire \core_1.execute.sreg_scratch.o_d[4] ;
 wire \core_1.execute.sreg_scratch.o_d[5] ;
 wire \core_1.execute.sreg_scratch.o_d[6] ;
 wire \core_1.execute.sreg_scratch.o_d[7] ;
 wire \core_1.execute.sreg_scratch.o_d[8] ;
 wire \core_1.execute.sreg_scratch.o_d[9] ;
 wire \core_1.execute.trap_flag ;
 wire \core_1.fetch.current_req_branch_pred ;
 wire \core_1.fetch.dbg_out ;
 wire \core_1.fetch.flush_event_invalidate ;
 wire \core_1.fetch.out_buffer_data_instr[0] ;
 wire \core_1.fetch.out_buffer_data_instr[10] ;
 wire \core_1.fetch.out_buffer_data_instr[11] ;
 wire \core_1.fetch.out_buffer_data_instr[12] ;
 wire \core_1.fetch.out_buffer_data_instr[13] ;
 wire \core_1.fetch.out_buffer_data_instr[14] ;
 wire \core_1.fetch.out_buffer_data_instr[15] ;
 wire \core_1.fetch.out_buffer_data_instr[16] ;
 wire \core_1.fetch.out_buffer_data_instr[17] ;
 wire \core_1.fetch.out_buffer_data_instr[18] ;
 wire \core_1.fetch.out_buffer_data_instr[19] ;
 wire \core_1.fetch.out_buffer_data_instr[1] ;
 wire \core_1.fetch.out_buffer_data_instr[20] ;
 wire \core_1.fetch.out_buffer_data_instr[21] ;
 wire \core_1.fetch.out_buffer_data_instr[22] ;
 wire \core_1.fetch.out_buffer_data_instr[23] ;
 wire \core_1.fetch.out_buffer_data_instr[24] ;
 wire \core_1.fetch.out_buffer_data_instr[25] ;
 wire \core_1.fetch.out_buffer_data_instr[26] ;
 wire \core_1.fetch.out_buffer_data_instr[27] ;
 wire \core_1.fetch.out_buffer_data_instr[28] ;
 wire \core_1.fetch.out_buffer_data_instr[29] ;
 wire \core_1.fetch.out_buffer_data_instr[2] ;
 wire \core_1.fetch.out_buffer_data_instr[30] ;
 wire \core_1.fetch.out_buffer_data_instr[31] ;
 wire \core_1.fetch.out_buffer_data_instr[3] ;
 wire \core_1.fetch.out_buffer_data_instr[4] ;
 wire \core_1.fetch.out_buffer_data_instr[5] ;
 wire \core_1.fetch.out_buffer_data_instr[6] ;
 wire \core_1.fetch.out_buffer_data_instr[7] ;
 wire \core_1.fetch.out_buffer_data_instr[8] ;
 wire \core_1.fetch.out_buffer_data_instr[9] ;
 wire \core_1.fetch.out_buffer_data_pred ;
 wire \core_1.fetch.out_buffer_valid ;
 wire \core_1.fetch.pc_flush_override ;
 wire \core_1.fetch.pc_reset_override ;
 wire \core_1.fetch.prev_req_branch_pred ;
 wire \core_1.fetch.prev_request_pc[0] ;
 wire \core_1.fetch.prev_request_pc[10] ;
 wire \core_1.fetch.prev_request_pc[11] ;
 wire \core_1.fetch.prev_request_pc[12] ;
 wire \core_1.fetch.prev_request_pc[13] ;
 wire \core_1.fetch.prev_request_pc[14] ;
 wire \core_1.fetch.prev_request_pc[15] ;
 wire \core_1.fetch.prev_request_pc[1] ;
 wire \core_1.fetch.prev_request_pc[2] ;
 wire \core_1.fetch.prev_request_pc[3] ;
 wire \core_1.fetch.prev_request_pc[4] ;
 wire \core_1.fetch.prev_request_pc[5] ;
 wire \core_1.fetch.prev_request_pc[6] ;
 wire \core_1.fetch.prev_request_pc[7] ;
 wire \core_1.fetch.prev_request_pc[8] ;
 wire \core_1.fetch.prev_request_pc[9] ;
 wire \core_1.fetch.submitable ;
 wire clknet_leaf_0_i_clk;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire clknet_leaf_1_i_clk;
 wire clknet_leaf_2_i_clk;
 wire clknet_leaf_3_i_clk;
 wire clknet_leaf_4_i_clk;
 wire clknet_leaf_5_i_clk;
 wire clknet_leaf_6_i_clk;
 wire clknet_leaf_7_i_clk;
 wire clknet_leaf_8_i_clk;
 wire clknet_leaf_9_i_clk;
 wire clknet_leaf_10_i_clk;
 wire clknet_leaf_11_i_clk;
 wire clknet_leaf_12_i_clk;
 wire clknet_leaf_13_i_clk;
 wire clknet_leaf_14_i_clk;
 wire clknet_leaf_15_i_clk;
 wire clknet_leaf_16_i_clk;
 wire clknet_leaf_17_i_clk;
 wire clknet_leaf_18_i_clk;
 wire clknet_leaf_19_i_clk;
 wire clknet_leaf_20_i_clk;
 wire clknet_leaf_21_i_clk;
 wire clknet_leaf_22_i_clk;
 wire clknet_leaf_23_i_clk;
 wire clknet_leaf_24_i_clk;
 wire clknet_leaf_25_i_clk;
 wire clknet_leaf_26_i_clk;
 wire clknet_leaf_27_i_clk;
 wire clknet_leaf_28_i_clk;
 wire clknet_leaf_29_i_clk;
 wire clknet_leaf_30_i_clk;
 wire clknet_leaf_31_i_clk;
 wire clknet_leaf_32_i_clk;
 wire clknet_leaf_33_i_clk;
 wire clknet_leaf_34_i_clk;
 wire clknet_leaf_35_i_clk;
 wire clknet_leaf_36_i_clk;
 wire clknet_leaf_37_i_clk;
 wire clknet_leaf_38_i_clk;
 wire clknet_leaf_39_i_clk;
 wire clknet_leaf_40_i_clk;
 wire clknet_leaf_41_i_clk;
 wire clknet_leaf_42_i_clk;
 wire clknet_leaf_43_i_clk;
 wire clknet_leaf_44_i_clk;
 wire clknet_leaf_45_i_clk;
 wire clknet_leaf_46_i_clk;
 wire clknet_leaf_47_i_clk;
 wire clknet_leaf_48_i_clk;
 wire clknet_leaf_49_i_clk;
 wire clknet_leaf_50_i_clk;
 wire clknet_0_i_clk;
 wire clknet_1_0_0_i_clk;
 wire clknet_1_0_1_i_clk;
 wire clknet_1_1_0_i_clk;
 wire clknet_1_1_1_i_clk;
 wire clknet_2_0_0_i_clk;
 wire clknet_2_1_0_i_clk;
 wire clknet_2_2_0_i_clk;
 wire clknet_2_3_0_i_clk;
 wire clknet_opt_1_0_i_clk;
 wire clknet_opt_1_1_i_clk;
 wire clknet_opt_2_0_i_clk;
 wire clknet_opt_2_1_i_clk;

 sky130_fd_sc_hd__buf_2 _3360_ (.A(\core_1.dec_r_reg_sel[2] ),
    .X(_0515_));
 sky130_fd_sc_hd__buf_2 _3361_ (.A(\core_1.dec_r_reg_sel[1] ),
    .X(_0516_));
 sky130_fd_sc_hd__buf_2 _3362_ (.A(\core_1.dec_r_reg_sel[0] ),
    .X(_0517_));
 sky130_fd_sc_hd__or3_2 _3363_ (.A(_0515_),
    .B(_0516_),
    .C(_0517_),
    .X(_0518_));
 sky130_fd_sc_hd__buf_6 _3364_ (.A(_0518_),
    .X(_0519_));
 sky130_fd_sc_hd__buf_6 _3365_ (.A(_0519_),
    .X(_0520_));
 sky130_fd_sc_hd__nor3b_4 _3366_ (.A(\core_1.dec_r_reg_sel[2] ),
    .B(_0517_),
    .C_N(_0516_),
    .Y(_0521_));
 sky130_fd_sc_hd__clkbuf_4 _3367_ (.A(_0521_),
    .X(_0522_));
 sky130_fd_sc_hd__buf_2 _3368_ (.A(_0515_),
    .X(_0523_));
 sky130_fd_sc_hd__clkbuf_2 _3369_ (.A(\core_1.dec_r_reg_sel[1] ),
    .X(_0524_));
 sky130_fd_sc_hd__clkbuf_2 _3370_ (.A(\core_1.dec_r_reg_sel[0] ),
    .X(_0525_));
 sky130_fd_sc_hd__and3b_4 _3371_ (.A_N(_0523_),
    .B(_0524_),
    .C(_0525_),
    .X(_0526_));
 sky130_fd_sc_hd__buf_2 _3372_ (.A(_0524_),
    .X(_0527_));
 sky130_fd_sc_hd__buf_2 _3373_ (.A(_0525_),
    .X(_0528_));
 sky130_fd_sc_hd__clkbuf_2 _3374_ (.A(_0523_),
    .X(_0529_));
 sky130_fd_sc_hd__and4b_1 _3375_ (.A_N(_0527_),
    .B(_0528_),
    .C(\core_1.execute.rf.reg_outputs[5][15] ),
    .D(_0529_),
    .X(_0530_));
 sky130_fd_sc_hd__a221o_2 _3376_ (.A1(\core_1.execute.rf.reg_outputs[2][15] ),
    .A2(_0522_),
    .B1(_0526_),
    .B2(\core_1.execute.rf.reg_outputs[3][15] ),
    .C1(_0530_),
    .X(_0531_));
 sky130_fd_sc_hd__buf_4 _3377_ (.A(_0524_),
    .X(_0532_));
 sky130_fd_sc_hd__buf_4 _3378_ (.A(_0525_),
    .X(_0533_));
 sky130_fd_sc_hd__nor2_2 _3379_ (.A(_0532_),
    .B(_0533_),
    .Y(_0534_));
 sky130_fd_sc_hd__or2b_1 _3380_ (.A(\core_1.execute.rf.reg_outputs[4][15] ),
    .B_N(_0529_),
    .X(_0535_));
 sky130_fd_sc_hd__buf_2 _3381_ (.A(_0515_),
    .X(_0536_));
 sky130_fd_sc_hd__buf_2 _3382_ (.A(_0524_),
    .X(_0537_));
 sky130_fd_sc_hd__buf_2 _3383_ (.A(_0525_),
    .X(_0538_));
 sky130_fd_sc_hd__and4_1 _3384_ (.A(\core_1.execute.rf.reg_outputs[7][15] ),
    .B(_0536_),
    .C(_0537_),
    .D(_0538_),
    .X(_0539_));
 sky130_fd_sc_hd__buf_2 _3385_ (.A(_0524_),
    .X(_0540_));
 sky130_fd_sc_hd__and4b_1 _3386_ (.A_N(_0528_),
    .B(_0540_),
    .C(_0536_),
    .D(\core_1.execute.rf.reg_outputs[6][15] ),
    .X(_0541_));
 sky130_fd_sc_hd__buf_2 _3387_ (.A(_0523_),
    .X(_0542_));
 sky130_fd_sc_hd__and4bb_1 _3388_ (.A_N(_0542_),
    .B_N(_0527_),
    .C(_0528_),
    .D(\core_1.execute.rf.reg_outputs[1][15] ),
    .X(_0543_));
 sky130_fd_sc_hd__a2111o_2 _3389_ (.A1(_0534_),
    .A2(_0535_),
    .B1(_0539_),
    .C1(_0541_),
    .D1(_0543_),
    .X(_0544_));
 sky130_fd_sc_hd__o22ai_4 _3390_ (.A1(net94),
    .A2(_0520_),
    .B1(_0531_),
    .B2(_0544_),
    .Y(_0545_));
 sky130_fd_sc_hd__inv_2 _3391_ (.A(_0545_),
    .Y(net200));
 sky130_fd_sc_hd__buf_4 _3392_ (.A(_0523_),
    .X(_0546_));
 sky130_fd_sc_hd__and4b_1 _3393_ (.A_N(_0532_),
    .B(_0533_),
    .C(\core_1.execute.rf.reg_outputs[5][14] ),
    .D(_0546_),
    .X(_0547_));
 sky130_fd_sc_hd__a221o_1 _3394_ (.A1(\core_1.execute.rf.reg_outputs[2][14] ),
    .A2(_0522_),
    .B1(_0526_),
    .B2(\core_1.execute.rf.reg_outputs[3][14] ),
    .C1(_0547_),
    .X(_0548_));
 sky130_fd_sc_hd__or2b_1 _3395_ (.A(\core_1.execute.rf.reg_outputs[4][14] ),
    .B_N(_0546_),
    .X(_0549_));
 sky130_fd_sc_hd__buf_2 _3396_ (.A(_0525_),
    .X(_0550_));
 sky130_fd_sc_hd__and4bb_1 _3397_ (.A_N(_0542_),
    .B_N(_0527_),
    .C(_0550_),
    .D(\core_1.execute.rf.reg_outputs[1][14] ),
    .X(_0551_));
 sky130_fd_sc_hd__and4b_1 _3398_ (.A_N(_0533_),
    .B(_0527_),
    .C(_0542_),
    .D(\core_1.execute.rf.reg_outputs[6][14] ),
    .X(_0552_));
 sky130_fd_sc_hd__and4_1 _3399_ (.A(\core_1.execute.rf.reg_outputs[7][14] ),
    .B(_0546_),
    .C(_0532_),
    .D(_0533_),
    .X(_0553_));
 sky130_fd_sc_hd__a2111o_1 _3400_ (.A1(_0534_),
    .A2(_0549_),
    .B1(_0551_),
    .C1(_0552_),
    .D1(_0553_),
    .X(_0554_));
 sky130_fd_sc_hd__or2_1 _3401_ (.A(_0548_),
    .B(_0554_),
    .X(_0555_));
 sky130_fd_sc_hd__o21ai_4 _3402_ (.A1(net93),
    .A2(_0520_),
    .B1(_0555_),
    .Y(_0556_));
 sky130_fd_sc_hd__clkinv_2 _3403_ (.A(_0556_),
    .Y(net199));
 sky130_fd_sc_hd__nor3b_2 _3404_ (.A(_0515_),
    .B(_0516_),
    .C_N(_0517_),
    .Y(_0557_));
 sky130_fd_sc_hd__buf_4 _3405_ (.A(_0557_),
    .X(_0558_));
 sky130_fd_sc_hd__and3b_4 _3406_ (.A_N(_0517_),
    .B(_0516_),
    .C(_0515_),
    .X(_0559_));
 sky130_fd_sc_hd__a22o_1 _3407_ (.A1(\core_1.execute.rf.reg_outputs[1][13] ),
    .A2(_0558_),
    .B1(_0559_),
    .B2(\core_1.execute.rf.reg_outputs[6][13] ),
    .X(_0560_));
 sky130_fd_sc_hd__and3b_1 _3408_ (.A_N(\core_1.dec_r_reg_sel[1] ),
    .B(\core_1.dec_r_reg_sel[0] ),
    .C(\core_1.dec_r_reg_sel[2] ),
    .X(_0561_));
 sky130_fd_sc_hd__buf_4 _3409_ (.A(_0561_),
    .X(_0562_));
 sky130_fd_sc_hd__nor3b_1 _3410_ (.A(_0516_),
    .B(_0517_),
    .C_N(\core_1.dec_r_reg_sel[2] ),
    .Y(_0563_));
 sky130_fd_sc_hd__buf_4 _3411_ (.A(_0563_),
    .X(_0564_));
 sky130_fd_sc_hd__a22o_1 _3412_ (.A1(\core_1.execute.rf.reg_outputs[5][13] ),
    .A2(_0562_),
    .B1(_0564_),
    .B2(\core_1.execute.rf.reg_outputs[4][13] ),
    .X(_0565_));
 sky130_fd_sc_hd__and4b_1 _3413_ (.A_N(_0523_),
    .B(_0524_),
    .C(_0525_),
    .D(\core_1.execute.rf.reg_outputs[3][13] ),
    .X(_0566_));
 sky130_fd_sc_hd__and4_1 _3414_ (.A(\core_1.execute.rf.reg_outputs[7][13] ),
    .B(_0523_),
    .C(_0524_),
    .D(_0525_),
    .X(_0567_));
 sky130_fd_sc_hd__nor3_2 _3415_ (.A(_0515_),
    .B(_0516_),
    .C(_0517_),
    .Y(_0568_));
 sky130_fd_sc_hd__buf_4 _3416_ (.A(_0568_),
    .X(_0569_));
 sky130_fd_sc_hd__a2111o_1 _3417_ (.A1(\core_1.execute.rf.reg_outputs[2][13] ),
    .A2(_0521_),
    .B1(_0566_),
    .C1(_0567_),
    .D1(_0569_),
    .X(_0570_));
 sky130_fd_sc_hd__o32ai_4 _3418_ (.A1(_0560_),
    .A2(_0565_),
    .A3(_0570_),
    .B1(_0519_),
    .B2(net92),
    .Y(_0571_));
 sky130_fd_sc_hd__clkinv_4 _3419_ (.A(_0571_),
    .Y(net198));
 sky130_fd_sc_hd__a22o_1 _3420_ (.A1(\core_1.execute.rf.reg_outputs[1][12] ),
    .A2(_0558_),
    .B1(_0559_),
    .B2(\core_1.execute.rf.reg_outputs[6][12] ),
    .X(_0572_));
 sky130_fd_sc_hd__a22o_1 _3421_ (.A1(\core_1.execute.rf.reg_outputs[5][12] ),
    .A2(_0562_),
    .B1(_0564_),
    .B2(\core_1.execute.rf.reg_outputs[4][12] ),
    .X(_0573_));
 sky130_fd_sc_hd__and4b_1 _3422_ (.A_N(_0542_),
    .B(_0527_),
    .C(_0550_),
    .D(\core_1.execute.rf.reg_outputs[3][12] ),
    .X(_0574_));
 sky130_fd_sc_hd__and4_1 _3423_ (.A(\core_1.execute.rf.reg_outputs[7][12] ),
    .B(_0542_),
    .C(_0527_),
    .D(_0550_),
    .X(_0575_));
 sky130_fd_sc_hd__a2111o_1 _3424_ (.A1(\core_1.execute.rf.reg_outputs[2][12] ),
    .A2(_0522_),
    .B1(_0574_),
    .C1(_0575_),
    .D1(_0569_),
    .X(_0576_));
 sky130_fd_sc_hd__o32ai_4 _3425_ (.A1(_0572_),
    .A2(_0573_),
    .A3(_0576_),
    .B1(_0520_),
    .B2(net91),
    .Y(_0577_));
 sky130_fd_sc_hd__inv_2 _3426_ (.A(_0577_),
    .Y(net197));
 sky130_fd_sc_hd__and4b_1 _3427_ (.A_N(_0540_),
    .B(_0528_),
    .C(\core_1.execute.rf.reg_outputs[5][11] ),
    .D(_0529_),
    .X(_0578_));
 sky130_fd_sc_hd__and4b_1 _3428_ (.A_N(_0550_),
    .B(_0540_),
    .C(_0529_),
    .D(\core_1.execute.rf.reg_outputs[6][11] ),
    .X(_0579_));
 sky130_fd_sc_hd__and4bb_1 _3429_ (.A_N(_0542_),
    .B_N(_0527_),
    .C(_0550_),
    .D(\core_1.execute.rf.reg_outputs[1][11] ),
    .X(_0580_));
 sky130_fd_sc_hd__a2111o_2 _3430_ (.A1(\core_1.execute.rf.reg_outputs[4][11] ),
    .A2(_0564_),
    .B1(_0578_),
    .C1(_0579_),
    .D1(_0580_),
    .X(_0581_));
 sky130_fd_sc_hd__and4b_1 _3431_ (.A_N(_0529_),
    .B(_0540_),
    .C(_0528_),
    .D(\core_1.execute.rf.reg_outputs[3][11] ),
    .X(_0582_));
 sky130_fd_sc_hd__and4_1 _3432_ (.A(\core_1.execute.rf.reg_outputs[7][11] ),
    .B(_0529_),
    .C(_0540_),
    .D(_0528_),
    .X(_0583_));
 sky130_fd_sc_hd__a2111o_1 _3433_ (.A1(\core_1.execute.rf.reg_outputs[2][11] ),
    .A2(_0522_),
    .B1(_0582_),
    .C1(_0583_),
    .D1(_0569_),
    .X(_0584_));
 sky130_fd_sc_hd__o22ai_4 _3434_ (.A1(net90),
    .A2(_0520_),
    .B1(_0581_),
    .B2(_0584_),
    .Y(_0585_));
 sky130_fd_sc_hd__clkinv_2 _3435_ (.A(_0585_),
    .Y(net196));
 sky130_fd_sc_hd__and4b_1 _3436_ (.A_N(_0550_),
    .B(_0527_),
    .C(_0542_),
    .D(\core_1.execute.rf.reg_outputs[6][10] ),
    .X(_0586_));
 sky130_fd_sc_hd__and4bb_1 _3437_ (.A_N(_0546_),
    .B_N(_0532_),
    .C(_0550_),
    .D(\core_1.execute.rf.reg_outputs[1][10] ),
    .X(_0587_));
 sky130_fd_sc_hd__and4b_1 _3438_ (.A_N(_0532_),
    .B(_0533_),
    .C(\core_1.execute.rf.reg_outputs[5][10] ),
    .D(_0546_),
    .X(_0588_));
 sky130_fd_sc_hd__a2111o_2 _3439_ (.A1(\core_1.execute.rf.reg_outputs[4][10] ),
    .A2(_0564_),
    .B1(_0586_),
    .C1(_0587_),
    .D1(_0588_),
    .X(_0589_));
 sky130_fd_sc_hd__and4_1 _3440_ (.A(\core_1.execute.rf.reg_outputs[7][10] ),
    .B(_0542_),
    .C(_0527_),
    .D(_0550_),
    .X(_0590_));
 sky130_fd_sc_hd__and4b_1 _3441_ (.A_N(_0546_),
    .B(_0527_),
    .C(_0550_),
    .D(\core_1.execute.rf.reg_outputs[3][10] ),
    .X(_0591_));
 sky130_fd_sc_hd__a2111o_1 _3442_ (.A1(\core_1.execute.rf.reg_outputs[2][10] ),
    .A2(_0522_),
    .B1(_0590_),
    .C1(_0591_),
    .D1(_0569_),
    .X(_0592_));
 sky130_fd_sc_hd__o22ai_4 _3443_ (.A1(net89),
    .A2(_0520_),
    .B1(_0589_),
    .B2(_0592_),
    .Y(_0593_));
 sky130_fd_sc_hd__clkinv_2 _3444_ (.A(_0593_),
    .Y(net195));
 sky130_fd_sc_hd__a22o_1 _3445_ (.A1(\core_1.execute.rf.reg_outputs[5][9] ),
    .A2(_0562_),
    .B1(_0564_),
    .B2(\core_1.execute.rf.reg_outputs[4][9] ),
    .X(_0594_));
 sky130_fd_sc_hd__a22o_1 _3446_ (.A1(\core_1.execute.rf.reg_outputs[1][9] ),
    .A2(_0558_),
    .B1(_0559_),
    .B2(\core_1.execute.rf.reg_outputs[6][9] ),
    .X(_0595_));
 sky130_fd_sc_hd__and4_1 _3447_ (.A(\core_1.execute.rf.reg_outputs[7][9] ),
    .B(_0536_),
    .C(_0537_),
    .D(_0538_),
    .X(_0596_));
 sky130_fd_sc_hd__and4b_1 _3448_ (.A_N(_0529_),
    .B(_0540_),
    .C(_0528_),
    .D(\core_1.execute.rf.reg_outputs[3][9] ),
    .X(_0597_));
 sky130_fd_sc_hd__a2111o_1 _3449_ (.A1(\core_1.execute.rf.reg_outputs[2][9] ),
    .A2(_0522_),
    .B1(_0596_),
    .C1(_0597_),
    .D1(_0569_),
    .X(_0598_));
 sky130_fd_sc_hd__or2_1 _3450_ (.A(net103),
    .B(_0519_),
    .X(_0599_));
 sky130_fd_sc_hd__o31ai_4 _3451_ (.A1(_0594_),
    .A2(_0595_),
    .A3(_0598_),
    .B1(_0599_),
    .Y(_0600_));
 sky130_fd_sc_hd__clkinv_2 _3452_ (.A(_0600_),
    .Y(net209));
 sky130_fd_sc_hd__a22o_1 _3453_ (.A1(\core_1.execute.rf.reg_outputs[1][8] ),
    .A2(_0557_),
    .B1(_0559_),
    .B2(\core_1.execute.rf.reg_outputs[6][8] ),
    .X(_0601_));
 sky130_fd_sc_hd__a22o_1 _3454_ (.A1(\core_1.execute.rf.reg_outputs[5][8] ),
    .A2(_0562_),
    .B1(_0564_),
    .B2(\core_1.execute.rf.reg_outputs[4][8] ),
    .X(_0602_));
 sky130_fd_sc_hd__and4_1 _3455_ (.A(\core_1.execute.rf.reg_outputs[7][8] ),
    .B(_0515_),
    .C(_0516_),
    .D(_0517_),
    .X(_0603_));
 sky130_fd_sc_hd__and4b_1 _3456_ (.A_N(_0515_),
    .B(_0516_),
    .C(_0517_),
    .D(\core_1.execute.rf.reg_outputs[3][8] ),
    .X(_0604_));
 sky130_fd_sc_hd__a2111o_1 _3457_ (.A1(\core_1.execute.rf.reg_outputs[2][8] ),
    .A2(_0521_),
    .B1(_0603_),
    .C1(_0604_),
    .D1(_0568_),
    .X(_0605_));
 sky130_fd_sc_hd__o32ai_4 _3458_ (.A1(_0601_),
    .A2(_0602_),
    .A3(_0605_),
    .B1(_0519_),
    .B2(net102),
    .Y(_0606_));
 sky130_fd_sc_hd__inv_2 _3459_ (.A(_0606_),
    .Y(net208));
 sky130_fd_sc_hd__and3_1 _3460_ (.A(_0523_),
    .B(_0524_),
    .C(_0525_),
    .X(_0607_));
 sky130_fd_sc_hd__a22o_1 _3461_ (.A1(\core_1.execute.rf.reg_outputs[5][7] ),
    .A2(_0562_),
    .B1(_0607_),
    .B2(\core_1.execute.rf.reg_outputs[7][7] ),
    .X(_0608_));
 sky130_fd_sc_hd__a22o_1 _3462_ (.A1(\core_1.execute.rf.reg_outputs[3][7] ),
    .A2(_0526_),
    .B1(_0558_),
    .B2(\core_1.execute.rf.reg_outputs[1][7] ),
    .X(_0609_));
 sky130_fd_sc_hd__and4bb_1 _3463_ (.A_N(_0532_),
    .B_N(_0533_),
    .C(\core_1.execute.rf.reg_outputs[4][7] ),
    .D(_0542_),
    .X(_0610_));
 sky130_fd_sc_hd__and4b_1 _3464_ (.A_N(_0533_),
    .B(_0532_),
    .C(_0546_),
    .D(\core_1.execute.rf.reg_outputs[6][7] ),
    .X(_0611_));
 sky130_fd_sc_hd__a2111o_1 _3465_ (.A1(\core_1.execute.rf.reg_outputs[2][7] ),
    .A2(_0522_),
    .B1(_0610_),
    .C1(_0611_),
    .D1(_0569_),
    .X(_0612_));
 sky130_fd_sc_hd__or2_1 _3466_ (.A(net101),
    .B(_0519_),
    .X(_0613_));
 sky130_fd_sc_hd__o31ai_4 _3467_ (.A1(_0608_),
    .A2(_0609_),
    .A3(_0612_),
    .B1(_0613_),
    .Y(_0614_));
 sky130_fd_sc_hd__clkinv_4 _3468_ (.A(_0614_),
    .Y(net207));
 sky130_fd_sc_hd__a22o_1 _3469_ (.A1(\core_1.execute.rf.reg_outputs[3][6] ),
    .A2(_0526_),
    .B1(_0558_),
    .B2(\core_1.execute.rf.reg_outputs[1][6] ),
    .X(_0615_));
 sky130_fd_sc_hd__a22o_1 _3470_ (.A1(\core_1.execute.rf.reg_outputs[5][6] ),
    .A2(_0562_),
    .B1(_0607_),
    .B2(\core_1.execute.rf.reg_outputs[7][6] ),
    .X(_0616_));
 sky130_fd_sc_hd__and4bb_1 _3471_ (.A_N(_0524_),
    .B_N(_0525_),
    .C(\core_1.execute.rf.reg_outputs[4][6] ),
    .D(_0515_),
    .X(_0617_));
 sky130_fd_sc_hd__and4b_1 _3472_ (.A_N(_0525_),
    .B(_0524_),
    .C(_0523_),
    .D(\core_1.execute.rf.reg_outputs[6][6] ),
    .X(_0618_));
 sky130_fd_sc_hd__a2111o_2 _3473_ (.A1(\core_1.execute.rf.reg_outputs[2][6] ),
    .A2(_0521_),
    .B1(_0617_),
    .C1(_0618_),
    .D1(_0568_),
    .X(_0619_));
 sky130_fd_sc_hd__or2_1 _3474_ (.A(net100),
    .B(_0519_),
    .X(_0620_));
 sky130_fd_sc_hd__o31ai_4 _3475_ (.A1(_0615_),
    .A2(_0616_),
    .A3(_0619_),
    .B1(_0620_),
    .Y(_0621_));
 sky130_fd_sc_hd__clkinv_4 _3476_ (.A(_0621_),
    .Y(net206));
 sky130_fd_sc_hd__a22o_1 _3477_ (.A1(\core_1.execute.rf.reg_outputs[5][5] ),
    .A2(_0562_),
    .B1(_0564_),
    .B2(\core_1.execute.rf.reg_outputs[4][5] ),
    .X(_0622_));
 sky130_fd_sc_hd__a22o_1 _3478_ (.A1(\core_1.execute.rf.reg_outputs[1][5] ),
    .A2(_0558_),
    .B1(_0559_),
    .B2(\core_1.execute.rf.reg_outputs[6][5] ),
    .X(_0623_));
 sky130_fd_sc_hd__and4b_1 _3479_ (.A_N(_0536_),
    .B(_0537_),
    .C(_0538_),
    .D(\core_1.execute.rf.reg_outputs[3][5] ),
    .X(_0624_));
 sky130_fd_sc_hd__and4_1 _3480_ (.A(\core_1.execute.rf.reg_outputs[7][5] ),
    .B(_0536_),
    .C(_0537_),
    .D(_0538_),
    .X(_0625_));
 sky130_fd_sc_hd__a2111o_1 _3481_ (.A1(\core_1.execute.rf.reg_outputs[2][5] ),
    .A2(_0521_),
    .B1(_0624_),
    .C1(_0625_),
    .D1(_0569_),
    .X(_0626_));
 sky130_fd_sc_hd__o32ai_4 _3482_ (.A1(_0622_),
    .A2(_0623_),
    .A3(_0626_),
    .B1(_0519_),
    .B2(net99),
    .Y(_0627_));
 sky130_fd_sc_hd__inv_2 _3483_ (.A(_0627_),
    .Y(net205));
 sky130_fd_sc_hd__a22o_1 _3484_ (.A1(\core_1.execute.rf.reg_outputs[5][4] ),
    .A2(_0562_),
    .B1(_0563_),
    .B2(\core_1.execute.rf.reg_outputs[4][4] ),
    .X(_0628_));
 sky130_fd_sc_hd__a22o_1 _3485_ (.A1(\core_1.execute.rf.reg_outputs[1][4] ),
    .A2(_0557_),
    .B1(_0559_),
    .B2(\core_1.execute.rf.reg_outputs[6][4] ),
    .X(_0629_));
 sky130_fd_sc_hd__and4b_1 _3486_ (.A_N(_0515_),
    .B(_0516_),
    .C(_0517_),
    .D(\core_1.execute.rf.reg_outputs[3][4] ),
    .X(_0630_));
 sky130_fd_sc_hd__and4_1 _3487_ (.A(\core_1.execute.rf.reg_outputs[7][4] ),
    .B(\core_1.dec_r_reg_sel[2] ),
    .C(_0516_),
    .D(_0517_),
    .X(_0631_));
 sky130_fd_sc_hd__a2111o_1 _3488_ (.A1(\core_1.execute.rf.reg_outputs[2][4] ),
    .A2(_0521_),
    .B1(_0630_),
    .C1(_0631_),
    .D1(_0568_),
    .X(_0632_));
 sky130_fd_sc_hd__o32ai_4 _3489_ (.A1(_0628_),
    .A2(_0629_),
    .A3(_0632_),
    .B1(_0518_),
    .B2(net98),
    .Y(_0633_));
 sky130_fd_sc_hd__inv_2 _3490_ (.A(_0633_),
    .Y(net204));
 sky130_fd_sc_hd__a22o_1 _3491_ (.A1(\core_1.execute.rf.reg_outputs[5][3] ),
    .A2(_0562_),
    .B1(_0564_),
    .B2(\core_1.execute.rf.reg_outputs[4][3] ),
    .X(_0634_));
 sky130_fd_sc_hd__a22o_1 _3492_ (.A1(\core_1.execute.rf.reg_outputs[3][3] ),
    .A2(_0526_),
    .B1(_0558_),
    .B2(\core_1.execute.rf.reg_outputs[1][3] ),
    .X(_0635_));
 sky130_fd_sc_hd__and4_1 _3493_ (.A(\core_1.execute.rf.reg_outputs[7][3] ),
    .B(_0536_),
    .C(_0537_),
    .D(_0538_),
    .X(_0636_));
 sky130_fd_sc_hd__and4b_1 _3494_ (.A_N(_0528_),
    .B(_0537_),
    .C(_0536_),
    .D(\core_1.execute.rf.reg_outputs[6][3] ),
    .X(_0637_));
 sky130_fd_sc_hd__a2111o_1 _3495_ (.A1(\core_1.execute.rf.reg_outputs[2][3] ),
    .A2(_0522_),
    .B1(_0636_),
    .C1(_0637_),
    .D1(_0569_),
    .X(_0638_));
 sky130_fd_sc_hd__o32a_4 _3496_ (.A1(_0634_),
    .A2(_0635_),
    .A3(_0638_),
    .B1(_0520_),
    .B2(net97),
    .X(_0639_));
 sky130_fd_sc_hd__clkbuf_8 _3497_ (.A(_0639_),
    .X(net203));
 sky130_fd_sc_hd__and4b_1 _3498_ (.A_N(_0542_),
    .B(_0540_),
    .C(_0528_),
    .D(\core_1.execute.rf.reg_outputs[3][2] ),
    .X(_0640_));
 sky130_fd_sc_hd__a221o_1 _3499_ (.A1(\core_1.execute.rf.reg_outputs[2][2] ),
    .A2(_0522_),
    .B1(_0558_),
    .B2(\core_1.execute.rf.reg_outputs[1][2] ),
    .C1(_0640_),
    .X(_0641_));
 sky130_fd_sc_hd__or2b_1 _3500_ (.A(\core_1.execute.rf.reg_outputs[4][2] ),
    .B_N(_0529_),
    .X(_0642_));
 sky130_fd_sc_hd__and4b_1 _3501_ (.A_N(_0540_),
    .B(_0538_),
    .C(\core_1.execute.rf.reg_outputs[5][2] ),
    .D(_0536_),
    .X(_0643_));
 sky130_fd_sc_hd__and4_1 _3502_ (.A(\core_1.execute.rf.reg_outputs[7][2] ),
    .B(_0529_),
    .C(_0540_),
    .D(_0528_),
    .X(_0644_));
 sky130_fd_sc_hd__and4b_1 _3503_ (.A_N(_0550_),
    .B(_0540_),
    .C(_0529_),
    .D(\core_1.execute.rf.reg_outputs[6][2] ),
    .X(_0645_));
 sky130_fd_sc_hd__a2111o_1 _3504_ (.A1(_0534_),
    .A2(_0642_),
    .B1(_0643_),
    .C1(_0644_),
    .D1(_0645_),
    .X(_0646_));
 sky130_fd_sc_hd__o22ai_4 _3505_ (.A1(net96),
    .A2(_0519_),
    .B1(_0641_),
    .B2(_0646_),
    .Y(_0647_));
 sky130_fd_sc_hd__inv_4 _3506_ (.A(_0647_),
    .Y(net202));
 sky130_fd_sc_hd__a22o_1 _3507_ (.A1(\core_1.execute.rf.reg_outputs[5][1] ),
    .A2(_0562_),
    .B1(_0564_),
    .B2(\core_1.execute.rf.reg_outputs[4][1] ),
    .X(_0648_));
 sky130_fd_sc_hd__a22o_1 _3508_ (.A1(\core_1.execute.rf.reg_outputs[3][1] ),
    .A2(_0526_),
    .B1(_0558_),
    .B2(\core_1.execute.rf.reg_outputs[1][1] ),
    .X(_0649_));
 sky130_fd_sc_hd__and4b_1 _3509_ (.A_N(_0538_),
    .B(_0537_),
    .C(_0536_),
    .D(\core_1.execute.rf.reg_outputs[6][1] ),
    .X(_0650_));
 sky130_fd_sc_hd__and4_1 _3510_ (.A(\core_1.execute.rf.reg_outputs[7][1] ),
    .B(_0536_),
    .C(_0537_),
    .D(_0538_),
    .X(_0651_));
 sky130_fd_sc_hd__a2111o_2 _3511_ (.A1(\core_1.execute.rf.reg_outputs[2][1] ),
    .A2(_0522_),
    .B1(_0650_),
    .C1(_0651_),
    .D1(_0569_),
    .X(_0652_));
 sky130_fd_sc_hd__or2_1 _3512_ (.A(net95),
    .B(_0519_),
    .X(_0653_));
 sky130_fd_sc_hd__o31a_1 _3513_ (.A1(_0648_),
    .A2(_0649_),
    .A3(_0652_),
    .B1(_0653_),
    .X(_0654_));
 sky130_fd_sc_hd__buf_6 _3514_ (.A(_0654_),
    .X(net201));
 sky130_fd_sc_hd__a22o_1 _3515_ (.A1(\core_1.execute.rf.reg_outputs[1][0] ),
    .A2(_0558_),
    .B1(_0559_),
    .B2(\core_1.execute.rf.reg_outputs[6][0] ),
    .X(_0655_));
 sky130_fd_sc_hd__a22o_1 _3516_ (.A1(\core_1.execute.rf.reg_outputs[2][0] ),
    .A2(_0521_),
    .B1(_0526_),
    .B2(\core_1.execute.rf.reg_outputs[3][0] ),
    .X(_0656_));
 sky130_fd_sc_hd__and4_1 _3517_ (.A(\core_1.execute.rf.reg_outputs[7][0] ),
    .B(_0523_),
    .C(_0537_),
    .D(_0538_),
    .X(_0657_));
 sky130_fd_sc_hd__and4b_1 _3518_ (.A_N(_0537_),
    .B(_0538_),
    .C(\core_1.execute.rf.reg_outputs[5][0] ),
    .D(_0523_),
    .X(_0658_));
 sky130_fd_sc_hd__a2111o_2 _3519_ (.A1(\core_1.execute.rf.reg_outputs[4][0] ),
    .A2(_0564_),
    .B1(_0657_),
    .C1(_0658_),
    .D1(_0569_),
    .X(_0659_));
 sky130_fd_sc_hd__or2_2 _3520_ (.A(net88),
    .B(_0519_),
    .X(_0660_));
 sky130_fd_sc_hd__o31ai_4 _3521_ (.A1(_0655_),
    .A2(_0656_),
    .A3(_0659_),
    .B1(_0660_),
    .Y(_0661_));
 sky130_fd_sc_hd__inv_4 _3522_ (.A(_0661_),
    .Y(net194));
 sky130_fd_sc_hd__inv_6 _3523_ (.A(net71),
    .Y(_0662_));
 sky130_fd_sc_hd__inv_2 _3524_ (.A(\core_1.fetch.dbg_out ),
    .Y(_0663_));
 sky130_fd_sc_hd__clkbuf_16 _3525_ (.A(\core_1.fetch.out_buffer_valid ),
    .X(_0664_));
 sky130_fd_sc_hd__clkbuf_16 _3526_ (.A(_0664_),
    .X(_0665_));
 sky130_fd_sc_hd__buf_4 _3527_ (.A(_0665_),
    .X(_0666_));
 sky130_fd_sc_hd__o21a_1 _3528_ (.A1(net19),
    .A2(net18),
    .B1(\core_1.execute.irq_en ),
    .X(_0667_));
 sky130_fd_sc_hd__or3_1 _3529_ (.A(net37),
    .B(\core_1.execute.sreg_irq_flags.i_d[2] ),
    .C(_0667_),
    .X(_0668_));
 sky130_fd_sc_hd__or2_1 _3530_ (.A(\core_1.execute.prev_sys ),
    .B(_0668_),
    .X(_0669_));
 sky130_fd_sc_hd__buf_6 _3531_ (.A(_0669_),
    .X(_0670_));
 sky130_fd_sc_hd__buf_4 _3532_ (.A(net105),
    .X(_0671_));
 sky130_fd_sc_hd__nand2_2 _3533_ (.A(\core_1.execute.pc_high_out[2] ),
    .B(_0671_),
    .Y(_0672_));
 sky130_fd_sc_hd__nand2_2 _3534_ (.A(\core_1.execute.pc_high_out[7] ),
    .B(_0671_),
    .Y(_0673_));
 sky130_fd_sc_hd__nand2_2 _3535_ (.A(\core_1.execute.pc_high_out[3] ),
    .B(net105),
    .Y(_0674_));
 sky130_fd_sc_hd__a2bb2o_1 _3536_ (.A1_N(\core_1.execute.prev_pc_high[7] ),
    .A2_N(_0673_),
    .B1(_0674_),
    .B2(\core_1.execute.prev_pc_high[3] ),
    .X(_0675_));
 sky130_fd_sc_hd__a221o_1 _3537_ (.A1(\core_1.execute.prev_pc_high[2] ),
    .A2(_0672_),
    .B1(_0673_),
    .B2(\core_1.execute.prev_pc_high[7] ),
    .C1(_0675_),
    .X(_0676_));
 sky130_fd_sc_hd__nand2_4 _3538_ (.A(\core_1.execute.pc_high_out[6] ),
    .B(_0671_),
    .Y(_0677_));
 sky130_fd_sc_hd__nand2_2 _3539_ (.A(\core_1.execute.pc_high_out[4] ),
    .B(net105),
    .Y(_0678_));
 sky130_fd_sc_hd__o2bb2a_1 _3540_ (.A1_N(\core_1.execute.prev_pc_high[6] ),
    .A2_N(_0677_),
    .B1(_0678_),
    .B2(\core_1.execute.prev_pc_high[4] ),
    .X(_0679_));
 sky130_fd_sc_hd__o221ai_1 _3541_ (.A1(\core_1.execute.prev_pc_high[6] ),
    .A2(_0677_),
    .B1(_0672_),
    .B2(\core_1.execute.prev_pc_high[2] ),
    .C1(_0679_),
    .Y(_0680_));
 sky130_fd_sc_hd__nand2_4 _3542_ (.A(\core_1.execute.pc_high_out[5] ),
    .B(net105),
    .Y(_0681_));
 sky130_fd_sc_hd__xnor2_1 _3543_ (.A(\core_1.execute.prev_pc_high[5] ),
    .B(_0681_),
    .Y(_0682_));
 sky130_fd_sc_hd__nand2_2 _3544_ (.A(\core_1.execute.pc_high_out[1] ),
    .B(net105),
    .Y(_0683_));
 sky130_fd_sc_hd__a2bb2o_1 _3545_ (.A1_N(\core_1.execute.prev_pc_high[1] ),
    .A2_N(_0683_),
    .B1(_0678_),
    .B2(\core_1.execute.prev_pc_high[4] ),
    .X(_0684_));
 sky130_fd_sc_hd__nand2_2 _3546_ (.A(\core_1.execute.pc_high_out[0] ),
    .B(_0671_),
    .Y(_0685_));
 sky130_fd_sc_hd__xnor2_1 _3547_ (.A(\core_1.execute.prev_pc_high[0] ),
    .B(_0685_),
    .Y(_0686_));
 sky130_fd_sc_hd__a2bb2o_1 _3548_ (.A1_N(\core_1.execute.prev_pc_high[3] ),
    .A2_N(_0674_),
    .B1(_0683_),
    .B2(\core_1.execute.prev_pc_high[1] ),
    .X(_0687_));
 sky130_fd_sc_hd__or4_1 _3549_ (.A(_0682_),
    .B(_0684_),
    .C(_0686_),
    .D(_0687_),
    .X(_0688_));
 sky130_fd_sc_hd__or3_4 _3550_ (.A(_0676_),
    .B(_0680_),
    .C(_0688_),
    .X(_0689_));
 sky130_fd_sc_hd__or2_1 _3551_ (.A(_0670_),
    .B(_0689_),
    .X(_0690_));
 sky130_fd_sc_hd__nor2_1 _3552_ (.A(\core_1.execute.hold_valid ),
    .B(\core_1.decode.o_submit ),
    .Y(_0691_));
 sky130_fd_sc_hd__or3_4 _3553_ (.A(\core_1.decode.i_flush ),
    .B(_0690_),
    .C(_0691_),
    .X(_0692_));
 sky130_fd_sc_hd__inv_2 _3554_ (.A(\core_1.execute.next_ready_delayed ),
    .Y(_0693_));
 sky130_fd_sc_hd__mux4_1 _3555_ (.A0(\core_1.ew_reg_ie[0] ),
    .A1(\core_1.ew_reg_ie[1] ),
    .A2(\core_1.ew_reg_ie[2] ),
    .A3(\core_1.ew_reg_ie[3] ),
    .S0(_0533_),
    .S1(_0532_),
    .X(_0694_));
 sky130_fd_sc_hd__clkinv_2 _3556_ (.A(_0546_),
    .Y(_0695_));
 sky130_fd_sc_hd__mux4_1 _3557_ (.A0(\core_1.ew_reg_ie[4] ),
    .A1(\core_1.ew_reg_ie[5] ),
    .A2(\core_1.ew_reg_ie[6] ),
    .A3(\core_1.ew_reg_ie[7] ),
    .S0(_0533_),
    .S1(_0532_),
    .X(_0696_));
 sky130_fd_sc_hd__or2_1 _3558_ (.A(_0695_),
    .B(_0696_),
    .X(_0697_));
 sky130_fd_sc_hd__o211a_1 _3559_ (.A1(_0546_),
    .A2(_0694_),
    .B1(_0697_),
    .C1(\core_1.dec_used_operands[1] ),
    .X(_0698_));
 sky130_fd_sc_hd__buf_4 _3560_ (.A(\core_1.dec_l_reg_sel[2] ),
    .X(_0699_));
 sky130_fd_sc_hd__inv_2 _3561_ (.A(_0699_),
    .Y(_0700_));
 sky130_fd_sc_hd__buf_4 _3562_ (.A(_0700_),
    .X(_0701_));
 sky130_fd_sc_hd__buf_4 _3563_ (.A(\core_1.dec_l_reg_sel[1] ),
    .X(_0702_));
 sky130_fd_sc_hd__buf_4 _3564_ (.A(\core_1.dec_l_reg_sel[0] ),
    .X(_0703_));
 sky130_fd_sc_hd__nand2_4 _3565_ (.A(_0702_),
    .B(_0703_),
    .Y(_0704_));
 sky130_fd_sc_hd__buf_2 _3566_ (.A(\core_1.dec_l_reg_sel[2] ),
    .X(_0705_));
 sky130_fd_sc_hd__buf_4 _3567_ (.A(_0705_),
    .X(_0706_));
 sky130_fd_sc_hd__buf_4 _3568_ (.A(_0703_),
    .X(_0707_));
 sky130_fd_sc_hd__buf_4 _3569_ (.A(_0707_),
    .X(_0708_));
 sky130_fd_sc_hd__buf_4 _3570_ (.A(\core_1.dec_l_reg_sel[1] ),
    .X(_0709_));
 sky130_fd_sc_hd__clkbuf_4 _3571_ (.A(_0709_),
    .X(_0710_));
 sky130_fd_sc_hd__and3b_1 _3572_ (.A_N(_0708_),
    .B(\core_1.ew_reg_ie[3] ),
    .C(_0710_),
    .X(_0711_));
 sky130_fd_sc_hd__nor2_8 _3573_ (.A(_0709_),
    .B(\core_1.dec_l_reg_sel[0] ),
    .Y(_0712_));
 sky130_fd_sc_hd__or2_1 _3574_ (.A(_0710_),
    .B(\core_1.ew_reg_ie[2] ),
    .X(_0713_));
 sky130_fd_sc_hd__a22o_1 _3575_ (.A1(\core_1.ew_reg_ie[1] ),
    .A2(_0712_),
    .B1(_0713_),
    .B2(_0708_),
    .X(_0714_));
 sky130_fd_sc_hd__or3_1 _3576_ (.A(_0706_),
    .B(_0711_),
    .C(_0714_),
    .X(_0715_));
 sky130_fd_sc_hd__and2_1 _3577_ (.A(_0701_),
    .B(_0704_),
    .X(_0716_));
 sky130_fd_sc_hd__mux4_1 _3578_ (.A0(\core_1.ew_reg_ie[5] ),
    .A1(\core_1.ew_reg_ie[6] ),
    .A2(\core_1.ew_reg_ie[7] ),
    .A3(\core_1.ew_reg_ie[4] ),
    .S0(_0708_),
    .S1(_0710_),
    .X(_0717_));
 sky130_fd_sc_hd__o211a_1 _3579_ (.A1(_0716_),
    .A2(_0717_),
    .B1(\core_1.execute.sreg_long_ptr_en ),
    .C1(\core_1.dec_mem_long ),
    .X(_0718_));
 sky130_fd_sc_hd__o211a_1 _3580_ (.A1(_0701_),
    .A2(_0704_),
    .B1(_0715_),
    .C1(_0718_),
    .X(_0719_));
 sky130_fd_sc_hd__or2_1 _3581_ (.A(_0710_),
    .B(_0708_),
    .X(_0720_));
 sky130_fd_sc_hd__or2b_4 _3582_ (.A(_0702_),
    .B_N(_0703_),
    .X(_0721_));
 sky130_fd_sc_hd__or3b_1 _3583_ (.A(_0708_),
    .B(\core_1.ew_reg_ie[2] ),
    .C_N(_0710_),
    .X(_0722_));
 sky130_fd_sc_hd__o221a_1 _3584_ (.A1(\core_1.ew_reg_ie[0] ),
    .A2(_0720_),
    .B1(_0721_),
    .B2(\core_1.ew_reg_ie[1] ),
    .C1(_0722_),
    .X(_0723_));
 sky130_fd_sc_hd__o211a_1 _3585_ (.A1(\core_1.ew_reg_ie[3] ),
    .A2(_0704_),
    .B1(_0723_),
    .C1(_0701_),
    .X(_0724_));
 sky130_fd_sc_hd__or3b_1 _3586_ (.A(_0708_),
    .B(\core_1.ew_reg_ie[6] ),
    .C_N(_0710_),
    .X(_0725_));
 sky130_fd_sc_hd__o221a_1 _3587_ (.A1(\core_1.ew_reg_ie[4] ),
    .A2(_0720_),
    .B1(_0721_),
    .B2(\core_1.ew_reg_ie[5] ),
    .C1(_0725_),
    .X(_0726_));
 sky130_fd_sc_hd__o211a_1 _3588_ (.A1(\core_1.ew_reg_ie[7] ),
    .A2(_0704_),
    .B1(_0726_),
    .C1(_0706_),
    .X(_0727_));
 sky130_fd_sc_hd__o31a_1 _3589_ (.A1(_0719_),
    .A2(_0724_),
    .A3(_0727_),
    .B1(\core_1.dec_used_operands[0] ),
    .X(_0728_));
 sky130_fd_sc_hd__o22a_4 _3590_ (.A1(\core_1.ew_submit ),
    .A2(_0693_),
    .B1(_0698_),
    .B2(_0728_),
    .X(_0729_));
 sky130_fd_sc_hd__inv_2 _3591_ (.A(net20),
    .Y(_0730_));
 sky130_fd_sc_hd__a22o_4 _3592_ (.A1(net156),
    .A2(_0730_),
    .B1(\core_1.ew_mem_access ),
    .B2(\core_1.ew_submit ),
    .X(_0731_));
 sky130_fd_sc_hd__or2_4 _3593_ (.A(\core_1.execute.alu_mul_div.i_div ),
    .B(\core_1.execute.alu_mul_div.i_mod ),
    .X(_0732_));
 sky130_fd_sc_hd__nand2_1 _3594_ (.A(\core_1.decode.o_submit ),
    .B(_0732_),
    .Y(_0733_));
 sky130_fd_sc_hd__nand2_4 _3595_ (.A(\core_1.decode.o_submit ),
    .B(\core_1.execute.alu_mul_div.i_mul ),
    .Y(_0734_));
 sky130_fd_sc_hd__nand2_2 _3596_ (.A(_0733_),
    .B(_0734_),
    .Y(_0735_));
 sky130_fd_sc_hd__or3_4 _3597_ (.A(\core_1.execute.alu_mul_div.comp ),
    .B(_0731_),
    .C(_0735_),
    .X(_0736_));
 sky130_fd_sc_hd__nor3_4 _3598_ (.A(_0729_),
    .B(_0736_),
    .C(_0692_),
    .Y(_0737_));
 sky130_fd_sc_hd__nor2_2 _3599_ (.A(_0692_),
    .B(_0737_),
    .Y(_0738_));
 sky130_fd_sc_hd__nor2_4 _3600_ (.A(\core_1.decode.input_valid ),
    .B(_0738_),
    .Y(_0739_));
 sky130_fd_sc_hd__mux2_8 _3601_ (.A0(net66),
    .A1(\core_1.fetch.out_buffer_data_instr[6] ),
    .S(_0665_),
    .X(_0740_));
 sky130_fd_sc_hd__mux2_8 _3602_ (.A0(net65),
    .A1(\core_1.fetch.out_buffer_data_instr[5] ),
    .S(_0665_),
    .X(_0741_));
 sky130_fd_sc_hd__mux2_8 _3603_ (.A0(net38),
    .A1(\core_1.fetch.out_buffer_data_instr[0] ),
    .S(_0664_),
    .X(_0742_));
 sky130_fd_sc_hd__mux2_8 _3604_ (.A0(net49),
    .A1(\core_1.fetch.out_buffer_data_instr[1] ),
    .S(_0664_),
    .X(_0743_));
 sky130_fd_sc_hd__or2b_1 _3605_ (.A(_0742_),
    .B_N(_0743_),
    .X(_0744_));
 sky130_fd_sc_hd__mux2_8 _3606_ (.A0(net60),
    .A1(\core_1.fetch.out_buffer_data_instr[2] ),
    .S(_0665_),
    .X(_0745_));
 sky130_fd_sc_hd__mux2_8 _3607_ (.A0(net63),
    .A1(\core_1.fetch.out_buffer_data_instr[3] ),
    .S(_0665_),
    .X(_0746_));
 sky130_fd_sc_hd__nand2_1 _3608_ (.A(_0745_),
    .B(_0746_),
    .Y(_0747_));
 sky130_fd_sc_hd__nor2_1 _3609_ (.A(_0744_),
    .B(_0747_),
    .Y(_0748_));
 sky130_fd_sc_hd__mux2_2 _3610_ (.A0(net54),
    .A1(\core_1.fetch.out_buffer_data_instr[24] ),
    .S(\core_1.fetch.out_buffer_valid ),
    .X(_0749_));
 sky130_fd_sc_hd__mux2_4 _3611_ (.A0(net56),
    .A1(\core_1.fetch.out_buffer_data_instr[26] ),
    .S(_0664_),
    .X(_0750_));
 sky130_fd_sc_hd__mux2_2 _3612_ (.A0(net46),
    .A1(\core_1.fetch.out_buffer_data_instr[17] ),
    .S(_0664_),
    .X(_0751_));
 sky130_fd_sc_hd__clkbuf_4 _3613_ (.A(\core_1.fetch.out_buffer_valid ),
    .X(_0752_));
 sky130_fd_sc_hd__or2b_1 _3614_ (.A(\core_1.fetch.out_buffer_data_instr[19] ),
    .B_N(_0752_),
    .X(_0753_));
 sky130_fd_sc_hd__o21a_1 _3615_ (.A1(_0664_),
    .A2(net48),
    .B1(_0753_),
    .X(_0754_));
 sky130_fd_sc_hd__or4b_1 _3616_ (.A(_0743_),
    .B(_0751_),
    .C(_0754_),
    .D_N(_0742_),
    .X(_0755_));
 sky130_fd_sc_hd__mux2_2 _3617_ (.A0(net53),
    .A1(\core_1.fetch.out_buffer_data_instr[23] ),
    .S(_0752_),
    .X(_0756_));
 sky130_fd_sc_hd__or2b_1 _3618_ (.A(\core_1.fetch.out_buffer_data_instr[18] ),
    .B_N(\core_1.fetch.out_buffer_valid ),
    .X(_0757_));
 sky130_fd_sc_hd__o21a_1 _3619_ (.A1(_0752_),
    .A2(net47),
    .B1(_0757_),
    .X(_0758_));
 sky130_fd_sc_hd__mux2_2 _3620_ (.A0(net50),
    .A1(\core_1.fetch.out_buffer_data_instr[20] ),
    .S(_0752_),
    .X(_0759_));
 sky130_fd_sc_hd__mux2_2 _3621_ (.A0(net61),
    .A1(\core_1.fetch.out_buffer_data_instr[30] ),
    .S(\core_1.fetch.out_buffer_valid ),
    .X(_0760_));
 sky130_fd_sc_hd__or4_1 _3622_ (.A(_0756_),
    .B(_0758_),
    .C(_0759_),
    .D(_0760_),
    .X(_0761_));
 sky130_fd_sc_hd__mux2_2 _3623_ (.A0(net51),
    .A1(\core_1.fetch.out_buffer_data_instr[21] ),
    .S(\core_1.fetch.out_buffer_valid ),
    .X(_0762_));
 sky130_fd_sc_hd__mux2_2 _3624_ (.A0(net45),
    .A1(\core_1.fetch.out_buffer_data_instr[16] ),
    .S(\core_1.fetch.out_buffer_valid ),
    .X(_0763_));
 sky130_fd_sc_hd__or2b_1 _3625_ (.A(\core_1.fetch.out_buffer_data_instr[28] ),
    .B_N(\core_1.fetch.out_buffer_valid ),
    .X(_0764_));
 sky130_fd_sc_hd__o21a_2 _3626_ (.A1(_0752_),
    .A2(net58),
    .B1(_0764_),
    .X(_0765_));
 sky130_fd_sc_hd__or2b_1 _3627_ (.A(\core_1.fetch.out_buffer_data_instr[31] ),
    .B_N(\core_1.fetch.out_buffer_valid ),
    .X(_0766_));
 sky130_fd_sc_hd__o21a_1 _3628_ (.A1(_0664_),
    .A2(net62),
    .B1(_0766_),
    .X(_0767_));
 sky130_fd_sc_hd__or4_1 _3629_ (.A(_0762_),
    .B(_0763_),
    .C(_0765_),
    .D(_0767_),
    .X(_0768_));
 sky130_fd_sc_hd__mux2_2 _3630_ (.A0(net52),
    .A1(\core_1.fetch.out_buffer_data_instr[22] ),
    .S(_0752_),
    .X(_0769_));
 sky130_fd_sc_hd__mux2_2 _3631_ (.A0(net57),
    .A1(\core_1.fetch.out_buffer_data_instr[27] ),
    .S(_0752_),
    .X(_0770_));
 sky130_fd_sc_hd__or2b_1 _3632_ (.A(\core_1.fetch.out_buffer_data_instr[25] ),
    .B_N(\core_1.fetch.out_buffer_valid ),
    .X(_0771_));
 sky130_fd_sc_hd__o21a_2 _3633_ (.A1(_0752_),
    .A2(net55),
    .B1(_0771_),
    .X(_0772_));
 sky130_fd_sc_hd__mux2_4 _3634_ (.A0(net59),
    .A1(\core_1.fetch.out_buffer_data_instr[29] ),
    .S(_0752_),
    .X(_0773_));
 sky130_fd_sc_hd__or4_1 _3635_ (.A(_0769_),
    .B(_0770_),
    .C(_0772_),
    .D(_0773_),
    .X(_0774_));
 sky130_fd_sc_hd__or3_1 _3636_ (.A(_0761_),
    .B(_0768_),
    .C(_0774_),
    .X(_0775_));
 sky130_fd_sc_hd__or4_1 _3637_ (.A(_0749_),
    .B(_0750_),
    .C(_0755_),
    .D(_0775_),
    .X(_0776_));
 sky130_fd_sc_hd__a211oi_1 _3638_ (.A1(_0744_),
    .A2(_0776_),
    .B1(_0745_),
    .C1(_0746_),
    .Y(_0777_));
 sky130_fd_sc_hd__nor2_1 _3639_ (.A(_0748_),
    .B(_0777_),
    .Y(_0778_));
 sky130_fd_sc_hd__mux2_8 _3640_ (.A0(net64),
    .A1(\core_1.fetch.out_buffer_data_instr[4] ),
    .S(_0665_),
    .X(_0779_));
 sky130_fd_sc_hd__or4b_1 _3641_ (.A(_0740_),
    .B(_0741_),
    .C(_0778_),
    .D_N(_0779_),
    .X(_0780_));
 sky130_fd_sc_hd__o211a_1 _3642_ (.A1(_0666_),
    .A2(net70),
    .B1(_0739_),
    .C1(_0780_),
    .X(_0781_));
 sky130_fd_sc_hd__a211o_2 _3643_ (.A1(\core_1.fetch.pc_flush_override ),
    .A2(_0663_),
    .B1(_0781_),
    .C1(\core_1.fetch.pc_reset_override ),
    .X(_0782_));
 sky130_fd_sc_hd__and2_1 _3644_ (.A(_0662_),
    .B(_0782_),
    .X(_0783_));
 sky130_fd_sc_hd__clkbuf_4 _3645_ (.A(_0783_),
    .X(_0784_));
 sky130_fd_sc_hd__buf_6 _3646_ (.A(_0784_),
    .X(net177));
 sky130_fd_sc_hd__buf_6 _3647_ (.A(\core_1.decode.i_flush ),
    .X(_0785_));
 sky130_fd_sc_hd__nor2_4 _3648_ (.A(\core_1.fetch.pc_flush_override ),
    .B(_0785_),
    .Y(_0786_));
 sky130_fd_sc_hd__clkbuf_4 _3649_ (.A(_0786_),
    .X(_0787_));
 sky130_fd_sc_hd__o21ai_1 _3650_ (.A1(_0665_),
    .A2(net55),
    .B1(_0771_),
    .Y(_0788_));
 sky130_fd_sc_hd__inv_2 _3651_ (.A(_0749_),
    .Y(_0789_));
 sky130_fd_sc_hd__a22oi_2 _3652_ (.A1(\core_1.fetch.prev_request_pc[9] ),
    .A2(_0788_),
    .B1(_0789_),
    .B2(\core_1.fetch.prev_request_pc[8] ),
    .Y(_0790_));
 sky130_fd_sc_hd__clkinv_2 _3653_ (.A(_0790_),
    .Y(_0791_));
 sky130_fd_sc_hd__inv_2 _3654_ (.A(\core_1.fetch.prev_request_pc[10] ),
    .Y(_0792_));
 sky130_fd_sc_hd__a2bb2o_1 _3655_ (.A1_N(\core_1.fetch.prev_request_pc[9] ),
    .A2_N(_0788_),
    .B1(_0750_),
    .B2(_0792_),
    .X(_0793_));
 sky130_fd_sc_hd__inv_2 _3656_ (.A(\core_1.fetch.prev_request_pc[13] ),
    .Y(_0794_));
 sky130_fd_sc_hd__inv_2 _3657_ (.A(\core_1.fetch.prev_request_pc[14] ),
    .Y(_0795_));
 sky130_fd_sc_hd__a22o_1 _3658_ (.A1(_0794_),
    .A2(_0773_),
    .B1(_0760_),
    .B2(_0795_),
    .X(_0796_));
 sky130_fd_sc_hd__o21ai_1 _3659_ (.A1(_0664_),
    .A2(net58),
    .B1(_0764_),
    .Y(_0797_));
 sky130_fd_sc_hd__nand2_1 _3660_ (.A(\core_1.fetch.prev_request_pc[12] ),
    .B(_0797_),
    .Y(_0798_));
 sky130_fd_sc_hd__o21ai_2 _3661_ (.A1(_0752_),
    .A2(net62),
    .B1(_0766_),
    .Y(_0799_));
 sky130_fd_sc_hd__o2bb2a_1 _3662_ (.A1_N(\core_1.fetch.prev_request_pc[15] ),
    .A2_N(_0799_),
    .B1(_0795_),
    .B2(_0760_),
    .X(_0800_));
 sky130_fd_sc_hd__o221a_1 _3663_ (.A1(\core_1.fetch.prev_request_pc[8] ),
    .A2(_0789_),
    .B1(_0799_),
    .B2(\core_1.fetch.prev_request_pc[15] ),
    .C1(_0800_),
    .X(_0801_));
 sky130_fd_sc_hd__o211a_1 _3664_ (.A1(_0794_),
    .A2(_0773_),
    .B1(_0798_),
    .C1(_0801_),
    .X(_0802_));
 sky130_fd_sc_hd__or2b_1 _3665_ (.A(_0796_),
    .B_N(_0802_),
    .X(_0803_));
 sky130_fd_sc_hd__inv_2 _3666_ (.A(\core_1.fetch.prev_request_pc[11] ),
    .Y(_0804_));
 sky130_fd_sc_hd__a2bb2o_1 _3667_ (.A1_N(\core_1.fetch.prev_request_pc[12] ),
    .A2_N(_0797_),
    .B1(_0804_),
    .B2(_0770_),
    .X(_0805_));
 sky130_fd_sc_hd__o22a_1 _3668_ (.A1(_0804_),
    .A2(_0770_),
    .B1(_0750_),
    .B2(_0792_),
    .X(_0806_));
 sky130_fd_sc_hd__or2b_1 _3669_ (.A(_0805_),
    .B_N(_0806_),
    .X(_0807_));
 sky130_fd_sc_hd__or4_1 _3670_ (.A(_0791_),
    .B(_0793_),
    .C(_0803_),
    .D(_0807_),
    .X(_0808_));
 sky130_fd_sc_hd__inv_2 _3671_ (.A(\core_1.fetch.prev_request_pc[7] ),
    .Y(_0809_));
 sky130_fd_sc_hd__and2_1 _3672_ (.A(_0809_),
    .B(_0756_),
    .X(_0810_));
 sky130_fd_sc_hd__inv_2 _3673_ (.A(\core_1.fetch.prev_request_pc[0] ),
    .Y(_0811_));
 sky130_fd_sc_hd__nor2_1 _3674_ (.A(_0811_),
    .B(_0763_),
    .Y(_0812_));
 sky130_fd_sc_hd__inv_2 _3675_ (.A(\core_1.fetch.prev_request_pc[1] ),
    .Y(_0813_));
 sky130_fd_sc_hd__o21ai_1 _3676_ (.A1(_0664_),
    .A2(net47),
    .B1(_0757_),
    .Y(_0814_));
 sky130_fd_sc_hd__nor2_1 _3677_ (.A(\core_1.fetch.prev_request_pc[2] ),
    .B(_0814_),
    .Y(_0815_));
 sky130_fd_sc_hd__a221o_1 _3678_ (.A1(_0813_),
    .A2(_0751_),
    .B1(_0763_),
    .B2(_0811_),
    .C1(_0815_),
    .X(_0816_));
 sky130_fd_sc_hd__nor2_1 _3679_ (.A(_0813_),
    .B(_0751_),
    .Y(_0817_));
 sky130_fd_sc_hd__inv_2 _3680_ (.A(\core_1.fetch.prev_request_pc[6] ),
    .Y(_0818_));
 sky130_fd_sc_hd__inv_2 _3681_ (.A(\core_1.fetch.prev_request_pc[5] ),
    .Y(_0819_));
 sky130_fd_sc_hd__a22o_1 _3682_ (.A1(_0818_),
    .A2(_0769_),
    .B1(_0762_),
    .B2(_0819_),
    .X(_0820_));
 sky130_fd_sc_hd__o21ai_1 _3683_ (.A1(_0664_),
    .A2(net48),
    .B1(_0753_),
    .Y(_0821_));
 sky130_fd_sc_hd__inv_2 _3684_ (.A(\core_1.fetch.prev_request_pc[4] ),
    .Y(_0822_));
 sky130_fd_sc_hd__a2bb2o_1 _3685_ (.A1_N(\core_1.fetch.prev_request_pc[3] ),
    .A2_N(_0821_),
    .B1(_0759_),
    .B2(_0822_),
    .X(_0823_));
 sky130_fd_sc_hd__o22a_1 _3686_ (.A1(_0818_),
    .A2(_0769_),
    .B1(_0756_),
    .B2(_0809_),
    .X(_0824_));
 sky130_fd_sc_hd__or3b_1 _3687_ (.A(_0820_),
    .B(_0823_),
    .C_N(_0824_),
    .X(_0825_));
 sky130_fd_sc_hd__a22oi_1 _3688_ (.A1(\core_1.fetch.prev_request_pc[3] ),
    .A2(_0821_),
    .B1(_0814_),
    .B2(\core_1.fetch.prev_request_pc[2] ),
    .Y(_0826_));
 sky130_fd_sc_hd__or4b_1 _3689_ (.A(_0816_),
    .B(_0817_),
    .C(_0825_),
    .D_N(_0826_),
    .X(_0827_));
 sky130_fd_sc_hd__o22a_1 _3690_ (.A1(_0819_),
    .A2(_0762_),
    .B1(_0759_),
    .B2(_0822_),
    .X(_0828_));
 sky130_fd_sc_hd__or4b_1 _3691_ (.A(_0810_),
    .B(_0812_),
    .C(_0827_),
    .D_N(_0828_),
    .X(_0829_));
 sky130_fd_sc_hd__or3_1 _3692_ (.A(_0813_),
    .B(_0751_),
    .C(_0815_),
    .X(_0830_));
 sky130_fd_sc_hd__a31o_1 _3693_ (.A1(_0816_),
    .A2(_0826_),
    .A3(_0830_),
    .B1(_0823_),
    .X(_0831_));
 sky130_fd_sc_hd__a21o_1 _3694_ (.A1(_0828_),
    .A2(_0831_),
    .B1(_0820_),
    .X(_0832_));
 sky130_fd_sc_hd__a211o_1 _3695_ (.A1(_0824_),
    .A2(_0832_),
    .B1(_0808_),
    .C1(_0810_),
    .X(_0833_));
 sky130_fd_sc_hd__o21a_1 _3696_ (.A1(_0790_),
    .A2(_0793_),
    .B1(_0806_),
    .X(_0834_));
 sky130_fd_sc_hd__o221a_1 _3697_ (.A1(_0794_),
    .A2(_0773_),
    .B1(_0805_),
    .B2(_0834_),
    .C1(_0798_),
    .X(_0835_));
 sky130_fd_sc_hd__o21ai_1 _3698_ (.A1(_0796_),
    .A2(_0835_),
    .B1(_0800_),
    .Y(_0836_));
 sky130_fd_sc_hd__o21ai_1 _3699_ (.A1(\core_1.fetch.prev_request_pc[15] ),
    .A2(_0799_),
    .B1(_0836_),
    .Y(_0837_));
 sky130_fd_sc_hd__a2bb2o_2 _3700_ (.A1_N(_0808_),
    .A2_N(_0829_),
    .B1(_0833_),
    .B2(_0837_),
    .X(_0838_));
 sky130_fd_sc_hd__mux2_4 _3701_ (.A0(net68),
    .A1(\core_1.fetch.out_buffer_data_instr[8] ),
    .S(_0665_),
    .X(_0839_));
 sky130_fd_sc_hd__mux2_4 _3702_ (.A0(net67),
    .A1(\core_1.fetch.out_buffer_data_instr[7] ),
    .S(_0665_),
    .X(_0840_));
 sky130_fd_sc_hd__mux2_1 _3703_ (.A0(net39),
    .A1(\core_1.fetch.out_buffer_data_instr[10] ),
    .S(_0665_),
    .X(_0841_));
 sky130_fd_sc_hd__mux2_4 _3704_ (.A0(net69),
    .A1(\core_1.fetch.out_buffer_data_instr[9] ),
    .S(_0666_),
    .X(_0842_));
 sky130_fd_sc_hd__o41a_1 _3705_ (.A1(_0839_),
    .A2(_0840_),
    .A3(_0841_),
    .A4(_0842_),
    .B1(_0748_),
    .X(_0843_));
 sky130_fd_sc_hd__or3_1 _3706_ (.A(\core_1.fetch.pc_reset_override ),
    .B(_0740_),
    .C(_0741_),
    .X(_0844_));
 sky130_fd_sc_hd__or4b_2 _3707_ (.A(_0779_),
    .B(_0747_),
    .C(_0844_),
    .D_N(_0743_),
    .X(_0845_));
 sky130_fd_sc_hd__a21oi_4 _3708_ (.A1(_0838_),
    .A2(_0843_),
    .B1(_0845_),
    .Y(_0846_));
 sky130_fd_sc_hd__buf_2 _3709_ (.A(_0846_),
    .X(_0847_));
 sky130_fd_sc_hd__buf_2 _3710_ (.A(_0847_),
    .X(_0848_));
 sky130_fd_sc_hd__or2_2 _3711_ (.A(\core_1.fetch.pc_flush_override ),
    .B(_0785_),
    .X(_0849_));
 sky130_fd_sc_hd__buf_2 _3712_ (.A(_0849_),
    .X(_0850_));
 sky130_fd_sc_hd__a21o_1 _3713_ (.A1(_0767_),
    .A2(_0848_),
    .B1(_0850_),
    .X(_0851_));
 sky130_fd_sc_hd__clkbuf_4 _3714_ (.A(_0847_),
    .X(_0852_));
 sky130_fd_sc_hd__and3_1 _3715_ (.A(\core_1.fetch.prev_request_pc[2] ),
    .B(\core_1.fetch.prev_request_pc[1] ),
    .C(\core_1.fetch.prev_request_pc[0] ),
    .X(_0853_));
 sky130_fd_sc_hd__and2_1 _3716_ (.A(\core_1.fetch.prev_request_pc[3] ),
    .B(_0853_),
    .X(_0854_));
 sky130_fd_sc_hd__and3_1 _3717_ (.A(\core_1.fetch.prev_request_pc[5] ),
    .B(\core_1.fetch.prev_request_pc[4] ),
    .C(_0854_),
    .X(_0855_));
 sky130_fd_sc_hd__and3_1 _3718_ (.A(\core_1.fetch.prev_request_pc[7] ),
    .B(\core_1.fetch.prev_request_pc[6] ),
    .C(_0855_),
    .X(_0856_));
 sky130_fd_sc_hd__and3_1 _3719_ (.A(\core_1.fetch.prev_request_pc[9] ),
    .B(\core_1.fetch.prev_request_pc[8] ),
    .C(_0856_),
    .X(_0857_));
 sky130_fd_sc_hd__nand2_1 _3720_ (.A(\core_1.fetch.prev_request_pc[10] ),
    .B(_0857_),
    .Y(_0858_));
 sky130_fd_sc_hd__nor2_1 _3721_ (.A(_0804_),
    .B(_0858_),
    .Y(_0859_));
 sky130_fd_sc_hd__and2_1 _3722_ (.A(\core_1.fetch.prev_request_pc[12] ),
    .B(_0859_),
    .X(_0860_));
 sky130_fd_sc_hd__nand2_1 _3723_ (.A(\core_1.fetch.prev_request_pc[13] ),
    .B(_0860_),
    .Y(_0861_));
 sky130_fd_sc_hd__nor2_1 _3724_ (.A(_0795_),
    .B(_0861_),
    .Y(_0862_));
 sky130_fd_sc_hd__xnor2_1 _3725_ (.A(\core_1.fetch.prev_request_pc[15] ),
    .B(_0862_),
    .Y(_0863_));
 sky130_fd_sc_hd__nor2_1 _3726_ (.A(_0852_),
    .B(_0863_),
    .Y(_0864_));
 sky130_fd_sc_hd__inv_2 _3727_ (.A(\core_1.fetch.pc_reset_override ),
    .Y(_0865_));
 sky130_fd_sc_hd__clkbuf_4 _3728_ (.A(_0865_),
    .X(_0866_));
 sky130_fd_sc_hd__o221a_1 _3729_ (.A1(net78),
    .A2(_0787_),
    .B1(_0851_),
    .B2(_0864_),
    .C1(_0866_),
    .X(net167));
 sky130_fd_sc_hd__and2_1 _3730_ (.A(_0795_),
    .B(_0861_),
    .X(_0867_));
 sky130_fd_sc_hd__nor3_1 _3731_ (.A(_0852_),
    .B(_0862_),
    .C(_0867_),
    .Y(_0868_));
 sky130_fd_sc_hd__a21o_1 _3732_ (.A1(_0760_),
    .A2(_0848_),
    .B1(_0850_),
    .X(_0869_));
 sky130_fd_sc_hd__o221a_1 _3733_ (.A1(net77),
    .A2(_0787_),
    .B1(_0868_),
    .B2(_0869_),
    .C1(_0866_),
    .X(net166));
 sky130_fd_sc_hd__o21ba_1 _3734_ (.A1(\core_1.fetch.prev_request_pc[13] ),
    .A2(_0860_),
    .B1_N(_0846_),
    .X(_0870_));
 sky130_fd_sc_hd__a221o_1 _3735_ (.A1(_0773_),
    .A2(_0848_),
    .B1(_0861_),
    .B2(_0870_),
    .C1(_0850_),
    .X(_0871_));
 sky130_fd_sc_hd__o211a_1 _3736_ (.A1(net76),
    .A2(_0787_),
    .B1(_0871_),
    .C1(_0866_),
    .X(net165));
 sky130_fd_sc_hd__nor2_1 _3737_ (.A(\core_1.fetch.prev_request_pc[12] ),
    .B(_0859_),
    .Y(_0872_));
 sky130_fd_sc_hd__nor3_1 _3738_ (.A(_0852_),
    .B(_0860_),
    .C(_0872_),
    .Y(_0873_));
 sky130_fd_sc_hd__a21o_1 _3739_ (.A1(_0765_),
    .A2(_0848_),
    .B1(_0850_),
    .X(_0874_));
 sky130_fd_sc_hd__o221a_1 _3740_ (.A1(net75),
    .A2(_0786_),
    .B1(_0873_),
    .B2(_0874_),
    .C1(_0865_),
    .X(net164));
 sky130_fd_sc_hd__and2_1 _3741_ (.A(_0804_),
    .B(_0858_),
    .X(_0875_));
 sky130_fd_sc_hd__nor3_1 _3742_ (.A(_0852_),
    .B(_0859_),
    .C(_0875_),
    .Y(_0876_));
 sky130_fd_sc_hd__a21o_1 _3743_ (.A1(_0770_),
    .A2(_0848_),
    .B1(_0850_),
    .X(_0877_));
 sky130_fd_sc_hd__o221a_1 _3744_ (.A1(net74),
    .A2(_0786_),
    .B1(_0876_),
    .B2(_0877_),
    .C1(_0865_),
    .X(net163));
 sky130_fd_sc_hd__o21ba_1 _3745_ (.A1(\core_1.fetch.prev_request_pc[10] ),
    .A2(_0857_),
    .B1_N(_0846_),
    .X(_0878_));
 sky130_fd_sc_hd__a221o_1 _3746_ (.A1(_0750_),
    .A2(_0848_),
    .B1(_0858_),
    .B2(_0878_),
    .C1(_0849_),
    .X(_0879_));
 sky130_fd_sc_hd__o211a_1 _3747_ (.A1(net73),
    .A2(_0787_),
    .B1(_0879_),
    .C1(_0866_),
    .X(net162));
 sky130_fd_sc_hd__and2_1 _3748_ (.A(\core_1.fetch.prev_request_pc[8] ),
    .B(_0856_),
    .X(_0880_));
 sky130_fd_sc_hd__nor2_1 _3749_ (.A(\core_1.fetch.prev_request_pc[9] ),
    .B(_0880_),
    .Y(_0881_));
 sky130_fd_sc_hd__o31a_1 _3750_ (.A1(_0846_),
    .A2(_0857_),
    .A3(_0881_),
    .B1(_0786_),
    .X(_0882_));
 sky130_fd_sc_hd__a21bo_1 _3751_ (.A1(_0772_),
    .A2(_0852_),
    .B1_N(_0882_),
    .X(_0883_));
 sky130_fd_sc_hd__o211a_1 _3752_ (.A1(net87),
    .A2(_0787_),
    .B1(_0883_),
    .C1(_0866_),
    .X(net176));
 sky130_fd_sc_hd__nor2_1 _3753_ (.A(\core_1.fetch.prev_request_pc[8] ),
    .B(_0856_),
    .Y(_0884_));
 sky130_fd_sc_hd__o31a_1 _3754_ (.A1(_0846_),
    .A2(_0880_),
    .A3(_0884_),
    .B1(_0786_),
    .X(_0885_));
 sky130_fd_sc_hd__a21bo_1 _3755_ (.A1(_0749_),
    .A2(_0852_),
    .B1_N(_0885_),
    .X(_0886_));
 sky130_fd_sc_hd__o211a_2 _3756_ (.A1(net86),
    .A2(_0787_),
    .B1(_0886_),
    .C1(_0866_),
    .X(net175));
 sky130_fd_sc_hd__and2_1 _3757_ (.A(\core_1.fetch.prev_request_pc[6] ),
    .B(_0855_),
    .X(_0887_));
 sky130_fd_sc_hd__nor2_1 _3758_ (.A(\core_1.fetch.prev_request_pc[7] ),
    .B(_0887_),
    .Y(_0888_));
 sky130_fd_sc_hd__nor3_1 _3759_ (.A(_0847_),
    .B(_0856_),
    .C(_0888_),
    .Y(_0889_));
 sky130_fd_sc_hd__a21o_1 _3760_ (.A1(_0756_),
    .A2(_0847_),
    .B1(_0849_),
    .X(_0890_));
 sky130_fd_sc_hd__o221a_2 _3761_ (.A1(net85),
    .A2(_0786_),
    .B1(_0889_),
    .B2(_0890_),
    .C1(_0865_),
    .X(net174));
 sky130_fd_sc_hd__nor2_1 _3762_ (.A(\core_1.fetch.prev_request_pc[6] ),
    .B(_0855_),
    .Y(_0891_));
 sky130_fd_sc_hd__nor3_1 _3763_ (.A(_0847_),
    .B(_0887_),
    .C(_0891_),
    .Y(_0892_));
 sky130_fd_sc_hd__a21o_1 _3764_ (.A1(_0769_),
    .A2(_0847_),
    .B1(_0849_),
    .X(_0893_));
 sky130_fd_sc_hd__o221a_4 _3765_ (.A1(net84),
    .A2(_0786_),
    .B1(_0892_),
    .B2(_0893_),
    .C1(_0865_),
    .X(net173));
 sky130_fd_sc_hd__a21oi_1 _3766_ (.A1(\core_1.fetch.prev_request_pc[4] ),
    .A2(_0854_),
    .B1(\core_1.fetch.prev_request_pc[5] ),
    .Y(_0894_));
 sky130_fd_sc_hd__nor3_1 _3767_ (.A(_0852_),
    .B(_0855_),
    .C(_0894_),
    .Y(_0895_));
 sky130_fd_sc_hd__a21o_1 _3768_ (.A1(_0762_),
    .A2(_0848_),
    .B1(_0850_),
    .X(_0896_));
 sky130_fd_sc_hd__o221a_4 _3769_ (.A1(net83),
    .A2(_0787_),
    .B1(_0895_),
    .B2(_0896_),
    .C1(_0866_),
    .X(net172));
 sky130_fd_sc_hd__xnor2_1 _3770_ (.A(\core_1.fetch.prev_request_pc[4] ),
    .B(_0854_),
    .Y(_0897_));
 sky130_fd_sc_hd__nor2_1 _3771_ (.A(_0852_),
    .B(_0897_),
    .Y(_0898_));
 sky130_fd_sc_hd__a21o_1 _3772_ (.A1(_0759_),
    .A2(_0848_),
    .B1(_0850_),
    .X(_0899_));
 sky130_fd_sc_hd__o221a_4 _3773_ (.A1(net82),
    .A2(_0787_),
    .B1(_0898_),
    .B2(_0899_),
    .C1(_0866_),
    .X(net171));
 sky130_fd_sc_hd__nor2_1 _3774_ (.A(\core_1.fetch.prev_request_pc[3] ),
    .B(_0853_),
    .Y(_0900_));
 sky130_fd_sc_hd__nor3_1 _3775_ (.A(_0847_),
    .B(_0854_),
    .C(_0900_),
    .Y(_0901_));
 sky130_fd_sc_hd__a21o_1 _3776_ (.A1(_0754_),
    .A2(_0847_),
    .B1(_0849_),
    .X(_0902_));
 sky130_fd_sc_hd__o221a_4 _3777_ (.A1(net81),
    .A2(_0786_),
    .B1(_0901_),
    .B2(_0902_),
    .C1(_0865_),
    .X(net170));
 sky130_fd_sc_hd__a21oi_1 _3778_ (.A1(\core_1.fetch.prev_request_pc[1] ),
    .A2(\core_1.fetch.prev_request_pc[0] ),
    .B1(\core_1.fetch.prev_request_pc[2] ),
    .Y(_0903_));
 sky130_fd_sc_hd__nor3_1 _3779_ (.A(_0852_),
    .B(_0853_),
    .C(_0903_),
    .Y(_0904_));
 sky130_fd_sc_hd__a21o_1 _3780_ (.A1(_0758_),
    .A2(_0848_),
    .B1(_0850_),
    .X(_0905_));
 sky130_fd_sc_hd__o221a_4 _3781_ (.A1(net80),
    .A2(_0787_),
    .B1(_0904_),
    .B2(_0905_),
    .C1(_0866_),
    .X(net169));
 sky130_fd_sc_hd__xnor2_1 _3782_ (.A(\core_1.fetch.prev_request_pc[1] ),
    .B(\core_1.fetch.prev_request_pc[0] ),
    .Y(_0906_));
 sky130_fd_sc_hd__nor2_1 _3783_ (.A(_0852_),
    .B(_0906_),
    .Y(_0907_));
 sky130_fd_sc_hd__a21o_1 _3784_ (.A1(_0751_),
    .A2(_0848_),
    .B1(_0850_),
    .X(_0908_));
 sky130_fd_sc_hd__o221a_4 _3785_ (.A1(net79),
    .A2(_0787_),
    .B1(_0907_),
    .B2(_0908_),
    .C1(_0866_),
    .X(net168));
 sky130_fd_sc_hd__nor2_1 _3786_ (.A(\core_1.fetch.prev_request_pc[0] ),
    .B(_0847_),
    .Y(_0909_));
 sky130_fd_sc_hd__a21o_1 _3787_ (.A1(_0763_),
    .A2(_0847_),
    .B1(_0849_),
    .X(_0910_));
 sky130_fd_sc_hd__o221a_4 _3788_ (.A1(net211),
    .A2(_0786_),
    .B1(_0909_),
    .B2(_0910_),
    .C1(_0865_),
    .X(net161));
 sky130_fd_sc_hd__inv_2 _3789_ (.A(_0685_),
    .Y(net108));
 sky130_fd_sc_hd__inv_2 _3790_ (.A(_0683_),
    .Y(net109));
 sky130_fd_sc_hd__inv_2 _3791_ (.A(_0672_),
    .Y(net110));
 sky130_fd_sc_hd__inv_2 _3792_ (.A(_0674_),
    .Y(net111));
 sky130_fd_sc_hd__inv_2 _3793_ (.A(_0678_),
    .Y(net112));
 sky130_fd_sc_hd__inv_2 _3794_ (.A(_0681_),
    .Y(net113));
 sky130_fd_sc_hd__inv_2 _3795_ (.A(_0677_),
    .Y(net114));
 sky130_fd_sc_hd__clkinv_2 _3796_ (.A(_0673_),
    .Y(net115));
 sky130_fd_sc_hd__nor2_2 _3797_ (.A(\core_1.decode.input_valid ),
    .B(\core_1.decode.i_submit ),
    .Y(_0911_));
 sky130_fd_sc_hd__nor3_4 _3798_ (.A(_0785_),
    .B(_0738_),
    .C(_0911_),
    .Y(_0912_));
 sky130_fd_sc_hd__nor2_4 _3799_ (.A(net71),
    .B(_0912_),
    .Y(_0913_));
 sky130_fd_sc_hd__clkbuf_4 _3800_ (.A(_0913_),
    .X(_0914_));
 sky130_fd_sc_hd__or3_4 _3801_ (.A(_0785_),
    .B(_0738_),
    .C(_0911_),
    .X(_0915_));
 sky130_fd_sc_hd__nor2_8 _3802_ (.A(net71),
    .B(_0915_),
    .Y(_0916_));
 sky130_fd_sc_hd__clkbuf_4 _3803_ (.A(_0916_),
    .X(_0917_));
 sky130_fd_sc_hd__clkbuf_4 _3804_ (.A(_0917_),
    .X(_0015_));
 sky130_fd_sc_hd__inv_2 _3805_ (.A(\core_1.decode.i_instr_l[1] ),
    .Y(_0918_));
 sky130_fd_sc_hd__nor2_2 _3806_ (.A(_0918_),
    .B(\core_1.decode.i_instr_l[0] ),
    .Y(_0919_));
 sky130_fd_sc_hd__or3b_2 _3807_ (.A(\core_1.decode.i_instr_l[6] ),
    .B(\core_1.decode.i_instr_l[5] ),
    .C_N(\core_1.decode.i_instr_l[4] ),
    .X(_0920_));
 sky130_fd_sc_hd__clkbuf_4 _3808_ (.A(_0920_),
    .X(_0921_));
 sky130_fd_sc_hd__nand2b_2 _3809_ (.A_N(\core_1.decode.i_instr_l[2] ),
    .B(\core_1.decode.i_instr_l[3] ),
    .Y(_0922_));
 sky130_fd_sc_hd__nor2_1 _3810_ (.A(_0921_),
    .B(_0922_),
    .Y(_0923_));
 sky130_fd_sc_hd__or3b_1 _3811_ (.A(\core_1.decode.i_instr_l[6] ),
    .B(\core_1.decode.i_instr_l[4] ),
    .C_N(\core_1.decode.i_instr_l[5] ),
    .X(_0924_));
 sky130_fd_sc_hd__buf_2 _3812_ (.A(_0924_),
    .X(_0925_));
 sky130_fd_sc_hd__nor2_1 _3813_ (.A(\core_1.decode.i_instr_l[1] ),
    .B(\core_1.decode.i_instr_l[0] ),
    .Y(_0926_));
 sky130_fd_sc_hd__nor2b_2 _3814_ (.A(\core_1.decode.i_instr_l[3] ),
    .B_N(\core_1.decode.i_instr_l[2] ),
    .Y(_0927_));
 sky130_fd_sc_hd__nand2_1 _3815_ (.A(_0926_),
    .B(_0927_),
    .Y(_0928_));
 sky130_fd_sc_hd__nor2_1 _3816_ (.A(_0925_),
    .B(_0928_),
    .Y(_0929_));
 sky130_fd_sc_hd__a21o_1 _3817_ (.A1(_0919_),
    .A2(_0923_),
    .B1(_0929_),
    .X(_0930_));
 sky130_fd_sc_hd__a22o_1 _3818_ (.A1(\core_1.decode.oc_alu_mode[1] ),
    .A2(_0914_),
    .B1(_0015_),
    .B2(_0930_),
    .X(_0004_));
 sky130_fd_sc_hd__clkbuf_4 _3819_ (.A(\core_1.decode.oc_alu_mode[6] ),
    .X(_0931_));
 sky130_fd_sc_hd__inv_2 _3820_ (.A(\core_1.decode.i_instr_l[0] ),
    .Y(_0932_));
 sky130_fd_sc_hd__nor2_2 _3821_ (.A(\core_1.decode.i_instr_l[1] ),
    .B(_0932_),
    .Y(_0933_));
 sky130_fd_sc_hd__nand2_1 _3822_ (.A(_0927_),
    .B(_0933_),
    .Y(_0934_));
 sky130_fd_sc_hd__or3_2 _3823_ (.A(\core_1.decode.i_instr_l[1] ),
    .B(\core_1.decode.i_instr_l[0] ),
    .C(_0922_),
    .X(_0935_));
 sky130_fd_sc_hd__a21oi_1 _3824_ (.A1(_0934_),
    .A2(_0935_),
    .B1(_0921_),
    .Y(_0936_));
 sky130_fd_sc_hd__a22o_1 _3825_ (.A1(_0931_),
    .A2(_0914_),
    .B1(_0015_),
    .B2(_0936_),
    .X(_0009_));
 sky130_fd_sc_hd__clkbuf_4 _3826_ (.A(\core_1.decode.oc_alu_mode[7] ),
    .X(_0937_));
 sky130_fd_sc_hd__nor3_4 _3827_ (.A(\core_1.decode.i_instr_l[6] ),
    .B(\core_1.decode.i_instr_l[4] ),
    .C(\core_1.decode.i_instr_l[5] ),
    .Y(_0938_));
 sky130_fd_sc_hd__and2_1 _3828_ (.A(\core_1.decode.i_instr_l[3] ),
    .B(\core_1.decode.i_instr_l[2] ),
    .X(_0939_));
 sky130_fd_sc_hd__and3_2 _3829_ (.A(_0919_),
    .B(_0938_),
    .C(_0939_),
    .X(_0940_));
 sky130_fd_sc_hd__nor2_1 _3830_ (.A(\core_1.decode.i_instr_l[3] ),
    .B(\core_1.decode.i_instr_l[2] ),
    .Y(_0941_));
 sky130_fd_sc_hd__nand2_1 _3831_ (.A(\core_1.decode.i_instr_l[1] ),
    .B(_0941_),
    .Y(_0942_));
 sky130_fd_sc_hd__or2_1 _3832_ (.A(\core_1.decode.i_instr_l[0] ),
    .B(_0942_),
    .X(_0943_));
 sky130_fd_sc_hd__nand2_1 _3833_ (.A(\core_1.decode.i_instr_l[3] ),
    .B(\core_1.decode.i_instr_l[2] ),
    .Y(_0944_));
 sky130_fd_sc_hd__or3_2 _3834_ (.A(_0918_),
    .B(_0932_),
    .C(_0944_),
    .X(_0945_));
 sky130_fd_sc_hd__or3_1 _3835_ (.A(\core_1.decode.i_instr_l[6] ),
    .B(\core_1.decode.i_instr_l[4] ),
    .C(\core_1.decode.i_instr_l[5] ),
    .X(_0946_));
 sky130_fd_sc_hd__buf_2 _3836_ (.A(_0946_),
    .X(_0947_));
 sky130_fd_sc_hd__a31o_1 _3837_ (.A1(_0928_),
    .A2(_0943_),
    .A3(_0945_),
    .B1(_0947_),
    .X(_0948_));
 sky130_fd_sc_hd__or2b_1 _3838_ (.A(_0940_),
    .B_N(_0948_),
    .X(_0949_));
 sky130_fd_sc_hd__nand2_1 _3839_ (.A(_0933_),
    .B(_0941_),
    .Y(_0950_));
 sky130_fd_sc_hd__nor2_1 _3840_ (.A(_0925_),
    .B(_0950_),
    .Y(_0951_));
 sky130_fd_sc_hd__a31o_1 _3841_ (.A1(_0927_),
    .A2(_0933_),
    .A3(_0938_),
    .B1(_0951_),
    .X(_0952_));
 sky130_fd_sc_hd__nor2_1 _3842_ (.A(_0920_),
    .B(_0945_),
    .Y(_0953_));
 sky130_fd_sc_hd__or3_1 _3843_ (.A(_0949_),
    .B(_0952_),
    .C(_0953_),
    .X(_0954_));
 sky130_fd_sc_hd__a22o_1 _3844_ (.A1(_0937_),
    .A2(_0914_),
    .B1(_0015_),
    .B2(_0954_),
    .X(_0010_));
 sky130_fd_sc_hd__buf_4 _3845_ (.A(_0916_),
    .X(_0955_));
 sky130_fd_sc_hd__and3b_1 _3846_ (.A_N(_0920_),
    .B(_0939_),
    .C(_0918_),
    .X(_0956_));
 sky130_fd_sc_hd__clkbuf_4 _3847_ (.A(_0913_),
    .X(_0957_));
 sky130_fd_sc_hd__clkbuf_4 _3848_ (.A(\core_1.execute.alu_mul_div.i_mul ),
    .X(_0958_));
 sky130_fd_sc_hd__clkbuf_4 _3849_ (.A(_0958_),
    .X(_0959_));
 sky130_fd_sc_hd__a32o_1 _3850_ (.A1(_0932_),
    .A2(_0955_),
    .A3(_0956_),
    .B1(_0957_),
    .B2(_0959_),
    .X(_0011_));
 sky130_fd_sc_hd__clkbuf_4 _3851_ (.A(\core_1.decode.oc_alu_mode[9] ),
    .X(_0960_));
 sky130_fd_sc_hd__and3_1 _3852_ (.A(\core_1.decode.i_instr_l[1] ),
    .B(\core_1.decode.i_instr_l[0] ),
    .C(_0927_),
    .X(_0961_));
 sky130_fd_sc_hd__or2b_1 _3853_ (.A(_0920_),
    .B_N(_0961_),
    .X(_0962_));
 sky130_fd_sc_hd__o21ai_1 _3854_ (.A1(_0928_),
    .A2(_0921_),
    .B1(_0962_),
    .Y(_0963_));
 sky130_fd_sc_hd__a22o_1 _3855_ (.A1(_0960_),
    .A2(_0914_),
    .B1(_0015_),
    .B2(_0963_),
    .X(_0012_));
 sky130_fd_sc_hd__buf_4 _3856_ (.A(\core_1.execute.alu_mul_div.i_mod ),
    .X(_0964_));
 sky130_fd_sc_hd__and3b_1 _3857_ (.A_N(_0925_),
    .B(_0926_),
    .C(_0939_),
    .X(_0965_));
 sky130_fd_sc_hd__a22o_1 _3858_ (.A1(_0964_),
    .A2(_0914_),
    .B1(_0015_),
    .B2(_0965_),
    .X(_0000_));
 sky130_fd_sc_hd__buf_4 _3859_ (.A(\core_1.decode.oc_alu_mode[4] ),
    .X(_0966_));
 sky130_fd_sc_hd__or2_1 _3860_ (.A(_0932_),
    .B(_0942_),
    .X(_0967_));
 sky130_fd_sc_hd__a21oi_1 _3861_ (.A1(_0935_),
    .A2(_0967_),
    .B1(_0947_),
    .Y(_0968_));
 sky130_fd_sc_hd__nor3_2 _3862_ (.A(_0932_),
    .B(_0922_),
    .C(_0947_),
    .Y(_0969_));
 sky130_fd_sc_hd__and2_1 _3863_ (.A(_0918_),
    .B(_0969_),
    .X(_0970_));
 sky130_fd_sc_hd__and2_1 _3864_ (.A(_0938_),
    .B(_0961_),
    .X(_0971_));
 sky130_fd_sc_hd__or2_1 _3865_ (.A(_0970_),
    .B(_0971_),
    .X(_0972_));
 sky130_fd_sc_hd__or2_1 _3866_ (.A(_0968_),
    .B(_0972_),
    .X(_0973_));
 sky130_fd_sc_hd__nor2_1 _3867_ (.A(_0925_),
    .B(_0943_),
    .Y(_0974_));
 sky130_fd_sc_hd__nand2_2 _3868_ (.A(_0927_),
    .B(_0919_),
    .Y(_0975_));
 sky130_fd_sc_hd__nor2_1 _3869_ (.A(_0947_),
    .B(_0975_),
    .Y(_0976_));
 sky130_fd_sc_hd__or2_1 _3870_ (.A(_0974_),
    .B(_0976_),
    .X(_0977_));
 sky130_fd_sc_hd__and3b_1 _3871_ (.A_N(_0925_),
    .B(_0926_),
    .C(_0941_),
    .X(_0978_));
 sky130_fd_sc_hd__nor2_2 _3872_ (.A(_0925_),
    .B(_0922_),
    .Y(_0979_));
 sky130_fd_sc_hd__or4_1 _3873_ (.A(_0973_),
    .B(_0977_),
    .C(_0978_),
    .D(_0979_),
    .X(_0980_));
 sky130_fd_sc_hd__a22o_1 _3874_ (.A1(_0966_),
    .A2(_0914_),
    .B1(_0015_),
    .B2(_0980_),
    .X(_0007_));
 sky130_fd_sc_hd__buf_4 _3875_ (.A(\core_1.decode.oc_alu_mode[11] ),
    .X(_0981_));
 sky130_fd_sc_hd__and3_1 _3876_ (.A(_0933_),
    .B(_0938_),
    .C(_0939_),
    .X(_0982_));
 sky130_fd_sc_hd__a21o_1 _3877_ (.A1(\core_1.decode.i_instr_l[1] ),
    .A2(_0969_),
    .B1(_0982_),
    .X(_0983_));
 sky130_fd_sc_hd__inv_2 _3878_ (.A(_0919_),
    .Y(_0984_));
 sky130_fd_sc_hd__nor3_1 _3879_ (.A(_0984_),
    .B(_0922_),
    .C(_0947_),
    .Y(_0985_));
 sky130_fd_sc_hd__a31o_1 _3880_ (.A1(_0926_),
    .A2(_0938_),
    .A3(_0939_),
    .B1(_0985_),
    .X(_0986_));
 sky130_fd_sc_hd__or2_1 _3881_ (.A(_0983_),
    .B(_0986_),
    .X(_0987_));
 sky130_fd_sc_hd__a22o_1 _3882_ (.A1(_0981_),
    .A2(_0914_),
    .B1(_0015_),
    .B2(_0987_),
    .X(_0001_));
 sky130_fd_sc_hd__buf_4 _3883_ (.A(\core_1.decode.oc_alu_mode[12] ),
    .X(_0988_));
 sky130_fd_sc_hd__nor2_1 _3884_ (.A(_0925_),
    .B(_0934_),
    .Y(_0989_));
 sky130_fd_sc_hd__nor2_1 _3885_ (.A(_0925_),
    .B(_0975_),
    .Y(_0990_));
 sky130_fd_sc_hd__or2_1 _3886_ (.A(_0989_),
    .B(_0990_),
    .X(_0991_));
 sky130_fd_sc_hd__a22o_1 _3887_ (.A1(_0988_),
    .A2(_0914_),
    .B1(_0015_),
    .B2(_0991_),
    .X(_0002_));
 sky130_fd_sc_hd__clkbuf_4 _3888_ (.A(\core_1.execute.alu_mul_div.i_div ),
    .X(_0992_));
 sky130_fd_sc_hd__a32o_1 _3889_ (.A1(\core_1.decode.i_instr_l[0] ),
    .A2(_0955_),
    .A3(_0956_),
    .B1(_0957_),
    .B2(_0992_),
    .X(_0008_));
 sky130_fd_sc_hd__buf_4 _3890_ (.A(_0913_),
    .X(_0993_));
 sky130_fd_sc_hd__nor2_1 _3891_ (.A(_0925_),
    .B(_0967_),
    .Y(_0994_));
 sky130_fd_sc_hd__a21o_1 _3892_ (.A1(_0923_),
    .A2(_0933_),
    .B1(_0994_),
    .X(_0995_));
 sky130_fd_sc_hd__a22o_1 _3893_ (.A1(\core_1.decode.oc_alu_mode[13] ),
    .A2(_0993_),
    .B1(_0015_),
    .B2(_0995_),
    .X(_0003_));
 sky130_fd_sc_hd__or2b_1 _3894_ (.A(_0925_),
    .B_N(_0961_),
    .X(_0996_));
 sky130_fd_sc_hd__nand2_1 _3895_ (.A(_0912_),
    .B(_0996_),
    .Y(_0997_));
 sky130_fd_sc_hd__clkbuf_8 _3896_ (.A(_0662_),
    .X(_0998_));
 sky130_fd_sc_hd__buf_4 _3897_ (.A(_0998_),
    .X(_0999_));
 sky130_fd_sc_hd__o211a_1 _3898_ (.A1(\core_1.decode.oc_alu_mode[3] ),
    .A2(_0912_),
    .B1(_0997_),
    .C1(_0999_),
    .X(_0006_));
 sky130_fd_sc_hd__buf_4 _3899_ (.A(\core_1.decode.oc_alu_mode[2] ),
    .X(_1000_));
 sky130_fd_sc_hd__buf_4 _3900_ (.A(_0917_),
    .X(_1001_));
 sky130_fd_sc_hd__nor2_1 _3901_ (.A(_0921_),
    .B(_0975_),
    .Y(_1002_));
 sky130_fd_sc_hd__and3_1 _3902_ (.A(\core_1.decode.i_instr_l[1] ),
    .B(\core_1.decode.i_instr_l[0] ),
    .C(_0923_),
    .X(_1003_));
 sky130_fd_sc_hd__nor2_1 _3903_ (.A(_0921_),
    .B(_0967_),
    .Y(_1004_));
 sky130_fd_sc_hd__or3_1 _3904_ (.A(_1002_),
    .B(_1003_),
    .C(_1004_),
    .X(_1005_));
 sky130_fd_sc_hd__a22o_1 _3905_ (.A1(_1000_),
    .A2(_0993_),
    .B1(_1001_),
    .B2(_1005_),
    .X(_0005_));
 sky130_fd_sc_hd__mux2_1 _3906_ (.A0(\core_1.fetch.prev_req_branch_pred ),
    .A1(_0846_),
    .S(net70),
    .X(_1006_));
 sky130_fd_sc_hd__clkbuf_1 _3907_ (.A(_1006_),
    .X(\core_1.fetch.current_req_branch_pred ));
 sky130_fd_sc_hd__nand2_4 _3908_ (.A(\core_1.ew_addr[0] ),
    .B(\core_1.ew_mem_width ),
    .Y(_1007_));
 sky130_fd_sc_hd__clkbuf_4 _3909_ (.A(_1007_),
    .X(_1008_));
 sky130_fd_sc_hd__clkbuf_4 _3910_ (.A(_1008_),
    .X(net157));
 sky130_fd_sc_hd__and2_1 _3911_ (.A(\core_1.ew_data[0] ),
    .B(net157),
    .X(_1009_));
 sky130_fd_sc_hd__clkbuf_1 _3912_ (.A(_1009_),
    .X(net139));
 sky130_fd_sc_hd__and2_1 _3913_ (.A(\core_1.ew_data[1] ),
    .B(net157),
    .X(_1010_));
 sky130_fd_sc_hd__clkbuf_1 _3914_ (.A(_1010_),
    .X(net146));
 sky130_fd_sc_hd__and2_1 _3915_ (.A(\core_1.ew_data[2] ),
    .B(net157),
    .X(_1011_));
 sky130_fd_sc_hd__clkbuf_1 _3916_ (.A(_1011_),
    .X(net147));
 sky130_fd_sc_hd__and2_1 _3917_ (.A(\core_1.ew_data[3] ),
    .B(net157),
    .X(_1012_));
 sky130_fd_sc_hd__clkbuf_1 _3918_ (.A(_1012_),
    .X(net148));
 sky130_fd_sc_hd__and2_1 _3919_ (.A(\core_1.ew_data[4] ),
    .B(net157),
    .X(_1013_));
 sky130_fd_sc_hd__clkbuf_1 _3920_ (.A(_1013_),
    .X(net149));
 sky130_fd_sc_hd__and2_1 _3921_ (.A(\core_1.ew_data[5] ),
    .B(net157),
    .X(_1014_));
 sky130_fd_sc_hd__clkbuf_1 _3922_ (.A(_1014_),
    .X(net150));
 sky130_fd_sc_hd__and2_1 _3923_ (.A(\core_1.ew_data[6] ),
    .B(net157),
    .X(_1015_));
 sky130_fd_sc_hd__clkbuf_1 _3924_ (.A(_1015_),
    .X(net151));
 sky130_fd_sc_hd__and2_1 _3925_ (.A(\core_1.ew_data[7] ),
    .B(net157),
    .X(_1016_));
 sky130_fd_sc_hd__clkbuf_1 _3926_ (.A(_1016_),
    .X(net152));
 sky130_fd_sc_hd__mux2_1 _3927_ (.A0(\core_1.ew_data[0] ),
    .A1(\core_1.ew_data[8] ),
    .S(net157),
    .X(_1017_));
 sky130_fd_sc_hd__clkbuf_1 _3928_ (.A(_1017_),
    .X(net153));
 sky130_fd_sc_hd__mux2_1 _3929_ (.A0(\core_1.ew_data[1] ),
    .A1(\core_1.ew_data[9] ),
    .S(_1008_),
    .X(_1018_));
 sky130_fd_sc_hd__clkbuf_1 _3930_ (.A(_1018_),
    .X(net154));
 sky130_fd_sc_hd__mux2_1 _3931_ (.A0(\core_1.ew_data[2] ),
    .A1(\core_1.ew_data[10] ),
    .S(_1008_),
    .X(_1019_));
 sky130_fd_sc_hd__clkbuf_1 _3932_ (.A(_1019_),
    .X(net140));
 sky130_fd_sc_hd__mux2_1 _3933_ (.A0(\core_1.ew_data[3] ),
    .A1(\core_1.ew_data[11] ),
    .S(_1008_),
    .X(_1020_));
 sky130_fd_sc_hd__clkbuf_1 _3934_ (.A(_1020_),
    .X(net141));
 sky130_fd_sc_hd__mux2_1 _3935_ (.A0(\core_1.ew_data[4] ),
    .A1(\core_1.ew_data[12] ),
    .S(_1008_),
    .X(_1021_));
 sky130_fd_sc_hd__clkbuf_1 _3936_ (.A(_1021_),
    .X(net142));
 sky130_fd_sc_hd__mux2_1 _3937_ (.A0(\core_1.ew_data[5] ),
    .A1(\core_1.ew_data[13] ),
    .S(_1008_),
    .X(_1022_));
 sky130_fd_sc_hd__clkbuf_1 _3938_ (.A(_1022_),
    .X(net143));
 sky130_fd_sc_hd__mux2_1 _3939_ (.A0(\core_1.ew_data[6] ),
    .A1(\core_1.ew_data[14] ),
    .S(_1008_),
    .X(_1023_));
 sky130_fd_sc_hd__clkbuf_1 _3940_ (.A(_1023_),
    .X(net144));
 sky130_fd_sc_hd__mux2_1 _3941_ (.A0(\core_1.ew_data[7] ),
    .A1(\core_1.ew_data[15] ),
    .S(_1008_),
    .X(_1024_));
 sky130_fd_sc_hd__clkbuf_1 _3942_ (.A(_1024_),
    .X(net145));
 sky130_fd_sc_hd__or2b_1 _3943_ (.A(\core_1.ew_addr[0] ),
    .B_N(\core_1.ew_mem_width ),
    .X(_1025_));
 sky130_fd_sc_hd__clkbuf_1 _3944_ (.A(_1025_),
    .X(net158));
 sky130_fd_sc_hd__inv_2 _3945_ (.A(net17),
    .Y(net160));
 sky130_fd_sc_hd__nor2_2 _3946_ (.A(_0785_),
    .B(\core_1.fetch.flush_event_invalidate ),
    .Y(_1026_));
 sky130_fd_sc_hd__o211ai_4 _3947_ (.A1(_0666_),
    .A2(net70),
    .B1(_0739_),
    .C1(_1026_),
    .Y(_1027_));
 sky130_fd_sc_hd__inv_2 _3948_ (.A(_1027_),
    .Y(\core_1.fetch.submitable ));
 sky130_fd_sc_hd__and2_2 _3949_ (.A(net155),
    .B(\core_1.ew_addr_high[0] ),
    .X(_1028_));
 sky130_fd_sc_hd__clkbuf_1 _3950_ (.A(_1028_),
    .X(net122));
 sky130_fd_sc_hd__clkbuf_8 _3951_ (.A(_0737_),
    .X(_1029_));
 sky130_fd_sc_hd__clkbuf_4 _3952_ (.A(_1029_),
    .X(_1030_));
 sky130_fd_sc_hd__inv_2 _3953_ (.A(\core_1.execute.alu_flag_reg.o_d[2] ),
    .Y(_1031_));
 sky130_fd_sc_hd__xor2_1 _3954_ (.A(\core_1.dec_jump_cond_code[1] ),
    .B(\core_1.dec_jump_cond_code[0] ),
    .X(_1032_));
 sky130_fd_sc_hd__inv_2 _3955_ (.A(\core_1.execute.alu_flag_reg.o_d[0] ),
    .Y(_1033_));
 sky130_fd_sc_hd__o221a_1 _3956_ (.A1(_1031_),
    .A2(\core_1.dec_jump_cond_code[0] ),
    .B1(_1032_),
    .B2(_1033_),
    .C1(\core_1.dec_jump_cond_code[2] ),
    .X(_1034_));
 sky130_fd_sc_hd__inv_2 _3957_ (.A(\core_1.dec_jump_cond_code[0] ),
    .Y(_1035_));
 sky130_fd_sc_hd__or4_1 _3958_ (.A(\core_1.execute.alu_flag_reg.o_d[2] ),
    .B(\core_1.execute.alu_flag_reg.o_d[0] ),
    .C(\core_1.dec_jump_cond_code[1] ),
    .D(_1035_),
    .X(_1036_));
 sky130_fd_sc_hd__a31o_1 _3959_ (.A1(_1033_),
    .A2(\core_1.dec_jump_cond_code[1] ),
    .A3(_1035_),
    .B1(\core_1.dec_jump_cond_code[2] ),
    .X(_1037_));
 sky130_fd_sc_hd__mux2_1 _3960_ (.A0(\core_1.execute.alu_flag_reg.o_d[1] ),
    .A1(\core_1.execute.alu_flag_reg.o_d[2] ),
    .S(\core_1.dec_jump_cond_code[1] ),
    .X(_1038_));
 sky130_fd_sc_hd__nor2_1 _3961_ (.A(_1035_),
    .B(_1038_),
    .Y(_1039_));
 sky130_fd_sc_hd__o2bb2a_1 _3962_ (.A1_N(_1034_),
    .A2_N(_1036_),
    .B1(_1037_),
    .B2(_1039_),
    .X(_1040_));
 sky130_fd_sc_hd__a21o_1 _3963_ (.A1(\core_1.execute.alu_flag_reg.o_d[0] ),
    .A2(_1035_),
    .B1(\core_1.execute.alu_flag_reg.o_d[1] ),
    .X(_1041_));
 sky130_fd_sc_hd__or4_1 _3964_ (.A(\core_1.execute.alu_flag_reg.o_d[3] ),
    .B(\core_1.dec_jump_cond_code[2] ),
    .C(\core_1.dec_jump_cond_code[1] ),
    .D(\core_1.dec_jump_cond_code[0] ),
    .X(_1042_));
 sky130_fd_sc_hd__o31ai_1 _3965_ (.A1(\core_1.execute.alu_flag_reg.o_d[4] ),
    .A2(\core_1.dec_jump_cond_code[1] ),
    .A3(_1035_),
    .B1(_1042_),
    .Y(_1043_));
 sky130_fd_sc_hd__nor2_1 _3966_ (.A(\core_1.execute.alu_flag_reg.o_d[1] ),
    .B(\core_1.execute.alu_flag_reg.o_d[0] ),
    .Y(_1044_));
 sky130_fd_sc_hd__o21a_1 _3967_ (.A1(\core_1.dec_jump_cond_code[0] ),
    .A2(_1044_),
    .B1(\core_1.dec_jump_cond_code[2] ),
    .X(_1045_));
 sky130_fd_sc_hd__a211o_1 _3968_ (.A1(\core_1.dec_jump_cond_code[1] ),
    .A2(_1041_),
    .B1(_1043_),
    .C1(_1045_),
    .X(_1046_));
 sky130_fd_sc_hd__mux2_1 _3969_ (.A0(_1040_),
    .A1(_1046_),
    .S(\core_1.dec_jump_cond_code[3] ),
    .X(_1047_));
 sky130_fd_sc_hd__xnor2_1 _3970_ (.A(\core_1.de_jmp_pred ),
    .B(_1047_),
    .Y(_1048_));
 sky130_fd_sc_hd__inv_2 _3971_ (.A(\core_1.execute.sreg_jtr_buff.o_d[0] ),
    .Y(_1049_));
 sky130_fd_sc_hd__inv_2 _3972_ (.A(net186),
    .Y(_1050_));
 sky130_fd_sc_hd__nor4_4 _3973_ (.A(net189),
    .B(net188),
    .C(net191),
    .D(net190),
    .Y(_1051_));
 sky130_fd_sc_hd__and3b_2 _3974_ (.A_N(net187),
    .B(_1050_),
    .C(_1051_),
    .X(_1052_));
 sky130_fd_sc_hd__nor4_4 _3975_ (.A(net182),
    .B(net181),
    .C(net184),
    .D(net183),
    .Y(_1053_));
 sky130_fd_sc_hd__nor4_4 _3976_ (.A(net193),
    .B(net192),
    .C(net180),
    .D(net179),
    .Y(_1054_));
 sky130_fd_sc_hd__and4bb_1 _3977_ (.A_N(net185),
    .B_N(net178),
    .C(_1053_),
    .D(_1054_),
    .X(_1055_));
 sky130_fd_sc_hd__buf_2 _3978_ (.A(_1055_),
    .X(_1056_));
 sky130_fd_sc_hd__buf_6 _3979_ (.A(\core_1.dec_sreg_irt ),
    .X(_1057_));
 sky130_fd_sc_hd__a31o_1 _3980_ (.A1(\core_1.dec_sreg_store ),
    .A2(_1052_),
    .A3(_1056_),
    .B1(_1057_),
    .X(_1058_));
 sky130_fd_sc_hd__o21a_2 _3981_ (.A1(\core_1.dec_jump_cond_code[4] ),
    .A2(_1058_),
    .B1(_0737_),
    .X(_1059_));
 sky130_fd_sc_hd__nor2_1 _3982_ (.A(net180),
    .B(net179),
    .Y(_1060_));
 sky130_fd_sc_hd__and4b_1 _3983_ (.A_N(net193),
    .B(net192),
    .C(_1060_),
    .D(\core_1.dec_sreg_store ),
    .X(_1061_));
 sky130_fd_sc_hd__and4_1 _3984_ (.A(_0737_),
    .B(_1051_),
    .C(_1053_),
    .D(_1061_),
    .X(_1062_));
 sky130_fd_sc_hd__a211o_1 _3985_ (.A1(_1049_),
    .A2(_1059_),
    .B1(_1062_),
    .C1(_0670_),
    .X(_1063_));
 sky130_fd_sc_hd__nand2_1 _3986_ (.A(\core_1.execute.sreg_jtr_buff.o_d[0] ),
    .B(_1059_),
    .Y(_1064_));
 sky130_fd_sc_hd__nor2_1 _3987_ (.A(net106),
    .B(_1064_),
    .Y(_1065_));
 sky130_fd_sc_hd__a211o_1 _3988_ (.A1(net106),
    .A2(_1063_),
    .B1(_1065_),
    .C1(_0689_),
    .X(_1066_));
 sky130_fd_sc_hd__a211o_1 _3989_ (.A1(\core_1.dec_jump_cond_code[4] ),
    .A2(_1048_),
    .B1(_1066_),
    .C1(_1058_),
    .X(_1067_));
 sky130_fd_sc_hd__a21o_1 _3990_ (.A1(_1030_),
    .A2(_1067_),
    .B1(_0690_),
    .X(_0013_));
 sky130_fd_sc_hd__buf_4 _3991_ (.A(_0662_),
    .X(_1068_));
 sky130_fd_sc_hd__and2_1 _3992_ (.A(_1068_),
    .B(_1066_),
    .X(_1069_));
 sky130_fd_sc_hd__clkbuf_1 _3993_ (.A(_1069_),
    .X(_0014_));
 sky130_fd_sc_hd__or3_1 _3994_ (.A(_0785_),
    .B(_0690_),
    .C(_0691_),
    .X(_1070_));
 sky130_fd_sc_hd__nor3_4 _3995_ (.A(_1070_),
    .B(_0729_),
    .C(_0736_),
    .Y(_1071_));
 sky130_fd_sc_hd__and3_1 _3996_ (.A(\core_1.execute.sreg_priv_control.o_d[0] ),
    .B(\core_1.dec_sreg_store ),
    .C(_1071_),
    .X(_1072_));
 sky130_fd_sc_hd__clkbuf_2 _3997_ (.A(_1072_),
    .X(net210));
 sky130_fd_sc_hd__or4_2 _3998_ (.A(_0915_),
    .B(_0984_),
    .C(_0921_),
    .D(_0944_),
    .X(_1073_));
 sky130_fd_sc_hd__or4_1 _3999_ (.A(_0918_),
    .B(_0915_),
    .C(_0947_),
    .D(_0944_),
    .X(_1074_));
 sky130_fd_sc_hd__buf_4 _4000_ (.A(_0998_),
    .X(_1075_));
 sky130_fd_sc_hd__o2111a_1 _4001_ (.A1(\core_1.dec_pc_inc ),
    .A2(_0912_),
    .B1(_1073_),
    .C1(_1074_),
    .D1(_1075_),
    .X(_0016_));
 sky130_fd_sc_hd__buf_4 _4002_ (.A(\core_1.dec_r_bus_imm ),
    .X(_1076_));
 sky130_fd_sc_hd__buf_6 _4003_ (.A(_1076_),
    .X(_1077_));
 sky130_fd_sc_hd__or2_1 _4004_ (.A(_0953_),
    .B(_0978_),
    .X(_1078_));
 sky130_fd_sc_hd__a31o_1 _4005_ (.A1(_0934_),
    .A2(_0942_),
    .A3(_0975_),
    .B1(_0947_),
    .X(_1079_));
 sky130_fd_sc_hd__or4b_1 _4006_ (.A(_0951_),
    .B(_0974_),
    .C(_1078_),
    .D_N(_1079_),
    .X(_1080_));
 sky130_fd_sc_hd__nor2_1 _4007_ (.A(_0935_),
    .B(_0947_),
    .Y(_1081_));
 sky130_fd_sc_hd__or4_1 _4008_ (.A(_1081_),
    .B(_0976_),
    .C(_0979_),
    .D(_0983_),
    .X(_1082_));
 sky130_fd_sc_hd__o21ai_1 _4009_ (.A1(_0920_),
    .A2(_0935_),
    .B1(_0962_),
    .Y(_1083_));
 sky130_fd_sc_hd__or4_1 _4010_ (.A(_1002_),
    .B(_1003_),
    .C(_1082_),
    .D(_1083_),
    .X(_1084_));
 sky130_fd_sc_hd__or2_1 _4011_ (.A(_0929_),
    .B(_0994_),
    .X(_1085_));
 sky130_fd_sc_hd__or3_1 _4012_ (.A(_0990_),
    .B(_1003_),
    .C(_1085_),
    .X(_1086_));
 sky130_fd_sc_hd__or4_1 _4013_ (.A(_0949_),
    .B(_1080_),
    .C(_1084_),
    .D(_1086_),
    .X(_1087_));
 sky130_fd_sc_hd__a22o_1 _4014_ (.A1(_1077_),
    .A2(_0993_),
    .B1(_1001_),
    .B2(_1087_),
    .X(_0017_));
 sky130_fd_sc_hd__o21a_1 _4015_ (.A1(_0919_),
    .A2(_0933_),
    .B1(_0923_),
    .X(_1088_));
 sky130_fd_sc_hd__or3_1 _4016_ (.A(_0994_),
    .B(_1003_),
    .C(_1088_),
    .X(_1089_));
 sky130_fd_sc_hd__or3b_1 _4017_ (.A(_0991_),
    .B(_1085_),
    .C_N(_0996_),
    .X(_1090_));
 sky130_fd_sc_hd__nor2_1 _4018_ (.A(_0921_),
    .B(_0934_),
    .Y(_1091_));
 sky130_fd_sc_hd__or3_1 _4019_ (.A(_1091_),
    .B(_1002_),
    .C(_1083_),
    .X(_1092_));
 sky130_fd_sc_hd__a21oi_1 _4020_ (.A1(_0928_),
    .A2(_0967_),
    .B1(_0921_),
    .Y(_1093_));
 sky130_fd_sc_hd__or4_1 _4021_ (.A(_1081_),
    .B(_0972_),
    .C(_1092_),
    .D(_1093_),
    .X(_1094_));
 sky130_fd_sc_hd__or4_2 _4022_ (.A(_0987_),
    .B(_1089_),
    .C(_1090_),
    .D(_1094_),
    .X(_1095_));
 sky130_fd_sc_hd__a22o_1 _4023_ (.A1(\core_1.dec_alu_flags_ie ),
    .A2(_0993_),
    .B1(_1001_),
    .B2(_1095_),
    .X(_0018_));
 sky130_fd_sc_hd__a22o_1 _4024_ (.A1(\core_1.dec_alu_carry_en ),
    .A2(_0993_),
    .B1(_1001_),
    .B2(_0969_),
    .X(_0019_));
 sky130_fd_sc_hd__a21o_2 _4025_ (.A1(\core_1.decode.i_instr_l[0] ),
    .A2(_0979_),
    .B1(_0977_),
    .X(_1096_));
 sky130_fd_sc_hd__or3_1 _4026_ (.A(_0956_),
    .B(_1083_),
    .C(_1089_),
    .X(_1097_));
 sky130_fd_sc_hd__inv_2 _4027_ (.A(_0950_),
    .Y(_1098_));
 sky130_fd_sc_hd__a221o_1 _4028_ (.A1(_0938_),
    .A2(_1098_),
    .B1(_0979_),
    .B2(_0932_),
    .C1(_0978_),
    .X(_1099_));
 sky130_fd_sc_hd__or4_1 _4029_ (.A(_0965_),
    .B(_0973_),
    .C(_1090_),
    .D(_1099_),
    .X(_1100_));
 sky130_fd_sc_hd__or3_4 _4030_ (.A(_1095_),
    .B(_1097_),
    .C(_1100_),
    .X(_1101_));
 sky130_fd_sc_hd__a22o_1 _4031_ (.A1(\core_1.decode.i_instr_l[13] ),
    .A2(_1096_),
    .B1(_1101_),
    .B2(\core_1.decode.i_instr_l[10] ),
    .X(_1102_));
 sky130_fd_sc_hd__a22o_1 _4032_ (.A1(_0708_),
    .A2(_0993_),
    .B1(_1001_),
    .B2(_1102_),
    .X(_0020_));
 sky130_fd_sc_hd__a22o_1 _4033_ (.A1(\core_1.decode.i_instr_l[14] ),
    .A2(_1096_),
    .B1(_1101_),
    .B2(\core_1.decode.i_instr_l[11] ),
    .X(_1103_));
 sky130_fd_sc_hd__a22o_1 _4034_ (.A1(_0710_),
    .A2(_0993_),
    .B1(_1001_),
    .B2(_1103_),
    .X(_0021_));
 sky130_fd_sc_hd__a22o_1 _4035_ (.A1(\core_1.decode.i_instr_l[15] ),
    .A2(_1096_),
    .B1(_1101_),
    .B2(\core_1.decode.i_instr_l[12] ),
    .X(_1104_));
 sky130_fd_sc_hd__a22o_1 _4036_ (.A1(_0706_),
    .A2(_0993_),
    .B1(_1001_),
    .B2(_1104_),
    .X(_0022_));
 sky130_fd_sc_hd__nor2_1 _4037_ (.A(_0921_),
    .B(_0950_),
    .Y(_1105_));
 sky130_fd_sc_hd__or2_1 _4038_ (.A(_0952_),
    .B(_1096_),
    .X(_1106_));
 sky130_fd_sc_hd__or2_4 _4039_ (.A(_1105_),
    .B(_1106_),
    .X(_1107_));
 sky130_fd_sc_hd__or4_1 _4040_ (.A(_1091_),
    .B(_0956_),
    .C(_0965_),
    .D(_0989_),
    .X(_1108_));
 sky130_fd_sc_hd__or3_1 _4041_ (.A(_1093_),
    .B(_1088_),
    .C(_1108_),
    .X(_1109_));
 sky130_fd_sc_hd__or4_4 _4042_ (.A(_0969_),
    .B(_0971_),
    .C(_0986_),
    .D(_1109_),
    .X(_1110_));
 sky130_fd_sc_hd__a22o_1 _4043_ (.A1(\core_1.decode.i_instr_l[10] ),
    .A2(_1107_),
    .B1(_1110_),
    .B2(\core_1.decode.i_instr_l[13] ),
    .X(_1111_));
 sky130_fd_sc_hd__a22o_1 _4044_ (.A1(_0533_),
    .A2(_0993_),
    .B1(_1001_),
    .B2(_1111_),
    .X(_0023_));
 sky130_fd_sc_hd__a22o_1 _4045_ (.A1(\core_1.decode.i_instr_l[11] ),
    .A2(_1107_),
    .B1(_1110_),
    .B2(\core_1.decode.i_instr_l[14] ),
    .X(_1112_));
 sky130_fd_sc_hd__a22o_1 _4046_ (.A1(_0532_),
    .A2(_0993_),
    .B1(_1001_),
    .B2(_1112_),
    .X(_0024_));
 sky130_fd_sc_hd__clkbuf_4 _4047_ (.A(_0913_),
    .X(_1113_));
 sky130_fd_sc_hd__a22o_1 _4048_ (.A1(\core_1.decode.i_instr_l[12] ),
    .A2(_1107_),
    .B1(_1110_),
    .B2(\core_1.decode.i_instr_l[15] ),
    .X(_1114_));
 sky130_fd_sc_hd__a22o_1 _4049_ (.A1(_0546_),
    .A2(_1113_),
    .B1(_1001_),
    .B2(_1114_),
    .X(_0025_));
 sky130_fd_sc_hd__and4b_1 _4050_ (.A_N(_0920_),
    .B(_0941_),
    .C(_0918_),
    .D(_0932_),
    .X(_1115_));
 sky130_fd_sc_hd__or4_1 _4051_ (.A(_0970_),
    .B(_0985_),
    .C(_1078_),
    .D(_1115_),
    .X(_1116_));
 sky130_fd_sc_hd__or4b_1 _4052_ (.A(_1092_),
    .B(_1093_),
    .C(_1116_),
    .D_N(_0948_),
    .X(_1117_));
 sky130_fd_sc_hd__or3_2 _4053_ (.A(_1100_),
    .B(_1109_),
    .C(_1117_),
    .X(_1118_));
 sky130_fd_sc_hd__and2b_1 _4054_ (.A_N(\core_1.decode.i_instr_l[8] ),
    .B(_1118_),
    .X(_1119_));
 sky130_fd_sc_hd__and3b_1 _4055_ (.A_N(\core_1.decode.i_instr_l[7] ),
    .B(_0912_),
    .C(_1119_),
    .X(_1120_));
 sky130_fd_sc_hd__buf_6 _4056_ (.A(net71),
    .X(_1121_));
 sky130_fd_sc_hd__buf_8 _4057_ (.A(_1121_),
    .X(_1122_));
 sky130_fd_sc_hd__nor2_2 _4058_ (.A(_1122_),
    .B(\core_1.decode.i_instr_l[9] ),
    .Y(_1123_));
 sky130_fd_sc_hd__a22o_1 _4059_ (.A1(\core_1.dec_rf_ie[0] ),
    .A2(_1113_),
    .B1(_1120_),
    .B2(_1123_),
    .X(_0026_));
 sky130_fd_sc_hd__and3_1 _4060_ (.A(\core_1.decode.i_instr_l[7] ),
    .B(_0912_),
    .C(_1119_),
    .X(_1124_));
 sky130_fd_sc_hd__a22o_1 _4061_ (.A1(\core_1.dec_rf_ie[1] ),
    .A2(_1113_),
    .B1(_1123_),
    .B2(_1124_),
    .X(_0027_));
 sky130_fd_sc_hd__and4b_1 _4062_ (.A_N(\core_1.decode.i_instr_l[7] ),
    .B(_0912_),
    .C(_1118_),
    .D(\core_1.decode.i_instr_l[8] ),
    .X(_1125_));
 sky130_fd_sc_hd__a22o_1 _4063_ (.A1(\core_1.dec_rf_ie[2] ),
    .A2(_1113_),
    .B1(_1123_),
    .B2(_1125_),
    .X(_0028_));
 sky130_fd_sc_hd__and4_1 _4064_ (.A(\core_1.decode.i_instr_l[8] ),
    .B(\core_1.decode.i_instr_l[7] ),
    .C(_0912_),
    .D(_1118_),
    .X(_1126_));
 sky130_fd_sc_hd__a22o_1 _4065_ (.A1(\core_1.dec_rf_ie[3] ),
    .A2(_1113_),
    .B1(_1123_),
    .B2(_1126_),
    .X(_0029_));
 sky130_fd_sc_hd__and2_1 _4066_ (.A(_0998_),
    .B(\core_1.decode.i_instr_l[9] ),
    .X(_1127_));
 sky130_fd_sc_hd__a22o_1 _4067_ (.A1(\core_1.dec_rf_ie[4] ),
    .A2(_1113_),
    .B1(_1120_),
    .B2(_1127_),
    .X(_0030_));
 sky130_fd_sc_hd__a22o_1 _4068_ (.A1(\core_1.dec_rf_ie[5] ),
    .A2(_1113_),
    .B1(_1124_),
    .B2(_1127_),
    .X(_0031_));
 sky130_fd_sc_hd__a22o_1 _4069_ (.A1(\core_1.dec_rf_ie[6] ),
    .A2(_1113_),
    .B1(_1125_),
    .B2(_1127_),
    .X(_0032_));
 sky130_fd_sc_hd__a22o_1 _4070_ (.A1(\core_1.dec_rf_ie[7] ),
    .A2(_1113_),
    .B1(_1126_),
    .B2(_1127_),
    .X(_0033_));
 sky130_fd_sc_hd__a32o_1 _4071_ (.A1(\core_1.decode.i_instr_l[7] ),
    .A2(_0917_),
    .A3(_0940_),
    .B1(_0957_),
    .B2(\core_1.dec_jump_cond_code[0] ),
    .X(_0034_));
 sky130_fd_sc_hd__a32o_1 _4072_ (.A1(\core_1.decode.i_instr_l[8] ),
    .A2(_0917_),
    .A3(_0940_),
    .B1(_0913_),
    .B2(\core_1.dec_jump_cond_code[1] ),
    .X(_0035_));
 sky130_fd_sc_hd__a32o_1 _4073_ (.A1(\core_1.decode.i_instr_l[9] ),
    .A2(_0917_),
    .A3(_0940_),
    .B1(_0913_),
    .B2(\core_1.dec_jump_cond_code[2] ),
    .X(_0036_));
 sky130_fd_sc_hd__a32o_1 _4074_ (.A1(\core_1.decode.i_instr_l[10] ),
    .A2(_0917_),
    .A3(_0940_),
    .B1(_0913_),
    .B2(\core_1.dec_jump_cond_code[3] ),
    .X(_0037_));
 sky130_fd_sc_hd__buf_4 _4075_ (.A(_1121_),
    .X(_1128_));
 sky130_fd_sc_hd__a2bb2o_1 _4076_ (.A1_N(_1128_),
    .A2_N(_1074_),
    .B1(_0914_),
    .B2(\core_1.dec_jump_cond_code[4] ),
    .X(_0038_));
 sky130_fd_sc_hd__mux2_1 _4077_ (.A0(net178),
    .A1(\core_1.decode.i_imm_pass[0] ),
    .S(_0917_),
    .X(_1129_));
 sky130_fd_sc_hd__clkbuf_1 _4078_ (.A(_1129_),
    .X(_0039_));
 sky130_fd_sc_hd__mux2_1 _4079_ (.A0(net185),
    .A1(\core_1.decode.i_imm_pass[1] ),
    .S(_0917_),
    .X(_1130_));
 sky130_fd_sc_hd__clkbuf_1 _4080_ (.A(_1130_),
    .X(_0040_));
 sky130_fd_sc_hd__mux2_1 _4081_ (.A0(net186),
    .A1(\core_1.decode.i_imm_pass[2] ),
    .S(_0917_),
    .X(_1131_));
 sky130_fd_sc_hd__clkbuf_1 _4082_ (.A(_1131_),
    .X(_0041_));
 sky130_fd_sc_hd__mux2_1 _4083_ (.A0(net187),
    .A1(\core_1.decode.i_imm_pass[3] ),
    .S(_0917_),
    .X(_1132_));
 sky130_fd_sc_hd__clkbuf_1 _4084_ (.A(_1132_),
    .X(_0042_));
 sky130_fd_sc_hd__buf_4 _4085_ (.A(_0916_),
    .X(_1133_));
 sky130_fd_sc_hd__mux2_1 _4086_ (.A0(net188),
    .A1(\core_1.decode.i_imm_pass[4] ),
    .S(_1133_),
    .X(_1134_));
 sky130_fd_sc_hd__clkbuf_1 _4087_ (.A(_1134_),
    .X(_0043_));
 sky130_fd_sc_hd__mux2_1 _4088_ (.A0(net189),
    .A1(\core_1.decode.i_imm_pass[5] ),
    .S(_1133_),
    .X(_1135_));
 sky130_fd_sc_hd__clkbuf_1 _4089_ (.A(_1135_),
    .X(_0044_));
 sky130_fd_sc_hd__mux2_1 _4090_ (.A0(net190),
    .A1(\core_1.decode.i_imm_pass[6] ),
    .S(_1133_),
    .X(_1136_));
 sky130_fd_sc_hd__clkbuf_1 _4091_ (.A(_1136_),
    .X(_0045_));
 sky130_fd_sc_hd__mux2_1 _4092_ (.A0(net191),
    .A1(\core_1.decode.i_imm_pass[7] ),
    .S(_1133_),
    .X(_1137_));
 sky130_fd_sc_hd__clkbuf_1 _4093_ (.A(_1137_),
    .X(_0046_));
 sky130_fd_sc_hd__mux2_1 _4094_ (.A0(net192),
    .A1(\core_1.decode.i_imm_pass[8] ),
    .S(_1133_),
    .X(_1138_));
 sky130_fd_sc_hd__clkbuf_1 _4095_ (.A(_1138_),
    .X(_0047_));
 sky130_fd_sc_hd__mux2_1 _4096_ (.A0(net193),
    .A1(\core_1.decode.i_imm_pass[9] ),
    .S(_1133_),
    .X(_1139_));
 sky130_fd_sc_hd__clkbuf_1 _4097_ (.A(_1139_),
    .X(_0048_));
 sky130_fd_sc_hd__mux2_1 _4098_ (.A0(net179),
    .A1(\core_1.decode.i_imm_pass[10] ),
    .S(_1133_),
    .X(_1140_));
 sky130_fd_sc_hd__clkbuf_1 _4099_ (.A(_1140_),
    .X(_0049_));
 sky130_fd_sc_hd__mux2_1 _4100_ (.A0(net180),
    .A1(\core_1.decode.i_imm_pass[11] ),
    .S(_1133_),
    .X(_1141_));
 sky130_fd_sc_hd__clkbuf_1 _4101_ (.A(_1141_),
    .X(_0050_));
 sky130_fd_sc_hd__mux2_1 _4102_ (.A0(net181),
    .A1(\core_1.decode.i_imm_pass[12] ),
    .S(_1133_),
    .X(_1142_));
 sky130_fd_sc_hd__clkbuf_1 _4103_ (.A(_1142_),
    .X(_0051_));
 sky130_fd_sc_hd__mux2_1 _4104_ (.A0(net182),
    .A1(\core_1.decode.i_imm_pass[13] ),
    .S(_1133_),
    .X(_1143_));
 sky130_fd_sc_hd__clkbuf_1 _4105_ (.A(_1143_),
    .X(_0052_));
 sky130_fd_sc_hd__mux2_1 _4106_ (.A0(net183),
    .A1(\core_1.decode.i_imm_pass[14] ),
    .S(_0916_),
    .X(_1144_));
 sky130_fd_sc_hd__clkbuf_1 _4107_ (.A(_1144_),
    .X(_0053_));
 sky130_fd_sc_hd__mux2_1 _4108_ (.A0(net184),
    .A1(\core_1.decode.i_imm_pass[15] ),
    .S(_0916_),
    .X(_1145_));
 sky130_fd_sc_hd__clkbuf_1 _4109_ (.A(_1145_),
    .X(_0054_));
 sky130_fd_sc_hd__buf_4 _4110_ (.A(\core_1.dec_mem_access ),
    .X(_1146_));
 sky130_fd_sc_hd__buf_6 _4111_ (.A(_1146_),
    .X(_1147_));
 sky130_fd_sc_hd__or2_1 _4112_ (.A(_0979_),
    .B(_1080_),
    .X(_1148_));
 sky130_fd_sc_hd__a22o_1 _4113_ (.A1(_1147_),
    .A2(_1113_),
    .B1(_0955_),
    .B2(_1148_),
    .X(_0055_));
 sky130_fd_sc_hd__a22o_1 _4114_ (.A1(\core_1.dec_mem_we ),
    .A2(_0957_),
    .B1(_0955_),
    .B2(_1106_),
    .X(_0056_));
 sky130_fd_sc_hd__or4_1 _4115_ (.A(_0968_),
    .B(_0982_),
    .C(_1002_),
    .D(_1083_),
    .X(_1149_));
 sky130_fd_sc_hd__or4_1 _4116_ (.A(_0997_),
    .B(_1086_),
    .C(_1099_),
    .D(_1149_),
    .X(_1150_));
 sky130_fd_sc_hd__or2_1 _4117_ (.A(\core_1.dec_used_operands[0] ),
    .B(_0912_),
    .X(_1151_));
 sky130_fd_sc_hd__o311a_1 _4118_ (.A1(_1096_),
    .A2(_1110_),
    .A3(_1150_),
    .B1(_1151_),
    .C1(_1075_),
    .X(_0057_));
 sky130_fd_sc_hd__o21ba_1 _4119_ (.A1(_1107_),
    .A2(_1110_),
    .B1_N(_1150_),
    .X(_1152_));
 sky130_fd_sc_hd__a22o_1 _4120_ (.A1(\core_1.dec_used_operands[1] ),
    .A2(_0957_),
    .B1(_1152_),
    .B2(_1075_),
    .X(_0058_));
 sky130_fd_sc_hd__a22o_1 _4121_ (.A1(\core_1.dec_sreg_load ),
    .A2(_0957_),
    .B1(_0955_),
    .B2(_1115_),
    .X(_0059_));
 sky130_fd_sc_hd__buf_4 _4122_ (.A(\core_1.dec_sreg_store ),
    .X(_1153_));
 sky130_fd_sc_hd__a22o_1 _4123_ (.A1(_1153_),
    .A2(_0957_),
    .B1(_0955_),
    .B2(_1105_),
    .X(_0060_));
 sky130_fd_sc_hd__inv_2 _4124_ (.A(_0945_),
    .Y(_1154_));
 sky130_fd_sc_hd__a32o_1 _4125_ (.A1(_0955_),
    .A2(_0938_),
    .A3(_1154_),
    .B1(_0913_),
    .B2(\core_1.dec_sreg_jal_over ),
    .X(_0061_));
 sky130_fd_sc_hd__buf_4 _4126_ (.A(_1057_),
    .X(_1155_));
 sky130_fd_sc_hd__a2bb2o_1 _4127_ (.A1_N(_1128_),
    .A2_N(_1073_),
    .B1(_0914_),
    .B2(_1155_),
    .X(_0062_));
 sky130_fd_sc_hd__nor2_1 _4128_ (.A(_0921_),
    .B(_0943_),
    .Y(_1156_));
 sky130_fd_sc_hd__a22o_1 _4129_ (.A1(\core_1.dec_sys ),
    .A2(_0957_),
    .B1(_0955_),
    .B2(_1156_),
    .X(_0063_));
 sky130_fd_sc_hd__a2111o_1 _4130_ (.A1(\core_1.decode.i_instr_l[1] ),
    .A2(_0979_),
    .B1(_1078_),
    .C1(_0951_),
    .D1(_0974_),
    .X(_1157_));
 sky130_fd_sc_hd__a22o_1 _4131_ (.A1(\core_1.dec_mem_width ),
    .A2(_0957_),
    .B1(_0955_),
    .B2(_1157_),
    .X(_0064_));
 sky130_fd_sc_hd__a22o_1 _4132_ (.A1(\core_1.dec_mem_long ),
    .A2(_0957_),
    .B1(_0955_),
    .B2(_0979_),
    .X(_0065_));
 sky130_fd_sc_hd__or2_1 _4133_ (.A(_1070_),
    .B(_1071_),
    .X(_1158_));
 sky130_fd_sc_hd__nor4_1 _4134_ (.A(_0785_),
    .B(_1122_),
    .C(_1158_),
    .D(_0911_),
    .Y(_0066_));
 sky130_fd_sc_hd__and4b_1 _4135_ (.A_N(net185),
    .B(net178),
    .C(_1053_),
    .D(_1054_),
    .X(_1159_));
 sky130_fd_sc_hd__buf_2 _4136_ (.A(_1159_),
    .X(_1160_));
 sky130_fd_sc_hd__and2_2 _4137_ (.A(_1052_),
    .B(_1160_),
    .X(_1161_));
 sky130_fd_sc_hd__buf_4 _4138_ (.A(_1161_),
    .X(_1162_));
 sky130_fd_sc_hd__nand2_2 _4139_ (.A(net210),
    .B(_1162_),
    .Y(_1163_));
 sky130_fd_sc_hd__nor2_8 _4140_ (.A(_1057_),
    .B(_1163_),
    .Y(_1164_));
 sky130_fd_sc_hd__nor2_4 _4141_ (.A(_0670_),
    .B(_1164_),
    .Y(_1165_));
 sky130_fd_sc_hd__buf_4 _4142_ (.A(_1165_),
    .X(_1166_));
 sky130_fd_sc_hd__buf_4 _4143_ (.A(_1164_),
    .X(_1167_));
 sky130_fd_sc_hd__or2_1 _4144_ (.A(net71),
    .B(_0670_),
    .X(_1168_));
 sky130_fd_sc_hd__a21o_1 _4145_ (.A1(net194),
    .A2(_1167_),
    .B1(_1168_),
    .X(_1169_));
 sky130_fd_sc_hd__a21o_1 _4146_ (.A1(\core_1.execute.sreg_priv_control.o_d[0] ),
    .A2(_1166_),
    .B1(_1169_),
    .X(_0067_));
 sky130_fd_sc_hd__a22o_1 _4147_ (.A1(net201),
    .A2(_1167_),
    .B1(_1166_),
    .B2(\core_1.execute.sreg_data_page ),
    .X(_1170_));
 sky130_fd_sc_hd__and2_1 _4148_ (.A(_1068_),
    .B(_1170_),
    .X(_1171_));
 sky130_fd_sc_hd__clkbuf_1 _4149_ (.A(_1171_),
    .X(_0068_));
 sky130_fd_sc_hd__a22o_1 _4150_ (.A1(net203),
    .A2(_1167_),
    .B1(_1166_),
    .B2(\core_1.execute.sreg_long_ptr_en ),
    .X(_1172_));
 sky130_fd_sc_hd__and2_1 _4151_ (.A(_1068_),
    .B(_1172_),
    .X(_1173_));
 sky130_fd_sc_hd__clkbuf_1 _4152_ (.A(_1173_),
    .X(_0069_));
 sky130_fd_sc_hd__a22o_1 _4153_ (.A1(net204),
    .A2(_1167_),
    .B1(_1166_),
    .B2(\core_1.execute.sreg_priv_control.o_d[4] ),
    .X(_1174_));
 sky130_fd_sc_hd__and2_1 _4154_ (.A(_1068_),
    .B(_1174_),
    .X(_1175_));
 sky130_fd_sc_hd__clkbuf_1 _4155_ (.A(_1175_),
    .X(_0070_));
 sky130_fd_sc_hd__a22o_1 _4156_ (.A1(net205),
    .A2(_1167_),
    .B1(_1166_),
    .B2(\core_1.execute.sreg_priv_control.o_d[5] ),
    .X(_1176_));
 sky130_fd_sc_hd__and2_1 _4157_ (.A(_1068_),
    .B(_1176_),
    .X(_1177_));
 sky130_fd_sc_hd__clkbuf_1 _4158_ (.A(_1177_),
    .X(_0071_));
 sky130_fd_sc_hd__a22o_1 _4159_ (.A1(net206),
    .A2(_1167_),
    .B1(_1166_),
    .B2(\core_1.execute.sreg_priv_control.o_d[6] ),
    .X(_1178_));
 sky130_fd_sc_hd__and2_1 _4160_ (.A(_1068_),
    .B(_1178_),
    .X(_1179_));
 sky130_fd_sc_hd__clkbuf_1 _4161_ (.A(_1179_),
    .X(_0072_));
 sky130_fd_sc_hd__a22o_1 _4162_ (.A1(net207),
    .A2(_1167_),
    .B1(_1166_),
    .B2(\core_1.execute.sreg_priv_control.o_d[7] ),
    .X(_1180_));
 sky130_fd_sc_hd__and2_1 _4163_ (.A(_1068_),
    .B(_1180_),
    .X(_1181_));
 sky130_fd_sc_hd__clkbuf_1 _4164_ (.A(_1181_),
    .X(_0073_));
 sky130_fd_sc_hd__a22o_1 _4165_ (.A1(net208),
    .A2(_1167_),
    .B1(_1166_),
    .B2(\core_1.execute.sreg_priv_control.o_d[8] ),
    .X(_1182_));
 sky130_fd_sc_hd__and2_1 _4166_ (.A(_1068_),
    .B(_1182_),
    .X(_1183_));
 sky130_fd_sc_hd__clkbuf_1 _4167_ (.A(_1183_),
    .X(_0074_));
 sky130_fd_sc_hd__buf_6 _4168_ (.A(_0998_),
    .X(_1184_));
 sky130_fd_sc_hd__a22o_1 _4169_ (.A1(net209),
    .A2(_1167_),
    .B1(_1166_),
    .B2(\core_1.execute.sreg_priv_control.o_d[9] ),
    .X(_1185_));
 sky130_fd_sc_hd__and2_1 _4170_ (.A(_1184_),
    .B(_1185_),
    .X(_1186_));
 sky130_fd_sc_hd__clkbuf_1 _4171_ (.A(_1186_),
    .X(_0075_));
 sky130_fd_sc_hd__a22o_1 _4172_ (.A1(net195),
    .A2(_1167_),
    .B1(_1166_),
    .B2(\core_1.execute.sreg_priv_control.o_d[10] ),
    .X(_1187_));
 sky130_fd_sc_hd__and2_1 _4173_ (.A(_1184_),
    .B(_1187_),
    .X(_1188_));
 sky130_fd_sc_hd__clkbuf_1 _4174_ (.A(_1188_),
    .X(_0076_));
 sky130_fd_sc_hd__a22o_1 _4175_ (.A1(net196),
    .A2(_1164_),
    .B1(_1165_),
    .B2(\core_1.execute.sreg_priv_control.o_d[11] ),
    .X(_1189_));
 sky130_fd_sc_hd__and2_1 _4176_ (.A(_1184_),
    .B(_1189_),
    .X(_1190_));
 sky130_fd_sc_hd__clkbuf_1 _4177_ (.A(_1190_),
    .X(_0077_));
 sky130_fd_sc_hd__a22o_1 _4178_ (.A1(net197),
    .A2(_1164_),
    .B1(_1165_),
    .B2(\core_1.execute.sreg_priv_control.o_d[12] ),
    .X(_1191_));
 sky130_fd_sc_hd__and2_1 _4179_ (.A(_1184_),
    .B(_1191_),
    .X(_1192_));
 sky130_fd_sc_hd__clkbuf_1 _4180_ (.A(_1192_),
    .X(_0078_));
 sky130_fd_sc_hd__a22o_1 _4181_ (.A1(net198),
    .A2(_1164_),
    .B1(_1165_),
    .B2(\core_1.execute.sreg_priv_control.o_d[13] ),
    .X(_1193_));
 sky130_fd_sc_hd__and2_1 _4182_ (.A(_1184_),
    .B(_1193_),
    .X(_1194_));
 sky130_fd_sc_hd__clkbuf_1 _4183_ (.A(_1194_),
    .X(_0079_));
 sky130_fd_sc_hd__a22o_1 _4184_ (.A1(net199),
    .A2(_1164_),
    .B1(_1165_),
    .B2(\core_1.execute.sreg_priv_control.o_d[14] ),
    .X(_1195_));
 sky130_fd_sc_hd__and2_1 _4185_ (.A(_1184_),
    .B(_1195_),
    .X(_1196_));
 sky130_fd_sc_hd__clkbuf_1 _4186_ (.A(_1196_),
    .X(_0080_));
 sky130_fd_sc_hd__a22o_1 _4187_ (.A1(net200),
    .A2(_1164_),
    .B1(_1165_),
    .B2(\core_1.execute.sreg_priv_control.o_d[15] ),
    .X(_1197_));
 sky130_fd_sc_hd__and2_1 _4188_ (.A(_1184_),
    .B(_1197_),
    .X(_1198_));
 sky130_fd_sc_hd__clkbuf_1 _4189_ (.A(_1198_),
    .X(_0081_));
 sky130_fd_sc_hd__clkbuf_4 _4190_ (.A(\core_1.execute.alu_mul_div.cbit[3] ),
    .X(_1199_));
 sky130_fd_sc_hd__buf_4 _4191_ (.A(_1199_),
    .X(_1200_));
 sky130_fd_sc_hd__clkinv_2 _4192_ (.A(\core_1.execute.alu_mul_div.cbit[2] ),
    .Y(_1201_));
 sky130_fd_sc_hd__buf_4 _4193_ (.A(_1201_),
    .X(_1202_));
 sky130_fd_sc_hd__clkbuf_4 _4194_ (.A(\core_1.execute.alu_mul_div.cbit[0] ),
    .X(_1203_));
 sky130_fd_sc_hd__clkbuf_4 _4195_ (.A(\core_1.execute.alu_mul_div.cbit[1] ),
    .X(_1204_));
 sky130_fd_sc_hd__nand2_2 _4196_ (.A(_1203_),
    .B(_1204_),
    .Y(_1205_));
 sky130_fd_sc_hd__nor2_2 _4197_ (.A(_1202_),
    .B(_1205_),
    .Y(_1206_));
 sky130_fd_sc_hd__nand2_4 _4198_ (.A(_1200_),
    .B(_1206_),
    .Y(_1207_));
 sky130_fd_sc_hd__clkbuf_4 _4199_ (.A(_1207_),
    .X(_1208_));
 sky130_fd_sc_hd__nor2_1 _4200_ (.A(\core_1.execute.alu_mul_div.comp ),
    .B(_0735_),
    .Y(_1209_));
 sky130_fd_sc_hd__or4_2 _4201_ (.A(_0785_),
    .B(net71),
    .C(_0690_),
    .D(_1209_),
    .X(_1210_));
 sky130_fd_sc_hd__o21ba_1 _4202_ (.A1(_0735_),
    .A2(_1208_),
    .B1_N(_1210_),
    .X(_0082_));
 sky130_fd_sc_hd__inv_2 _4203_ (.A(_1026_),
    .Y(_1211_));
 sky130_fd_sc_hd__or4b_1 _4204_ (.A(net71),
    .B(_0739_),
    .C(_1211_),
    .D_N(net70),
    .X(_1212_));
 sky130_fd_sc_hd__buf_4 _4205_ (.A(_1212_),
    .X(_1213_));
 sky130_fd_sc_hd__buf_6 _4206_ (.A(_1213_),
    .X(_1214_));
 sky130_fd_sc_hd__mux2_1 _4207_ (.A0(net38),
    .A1(\core_1.fetch.out_buffer_data_instr[0] ),
    .S(_1214_),
    .X(_1215_));
 sky130_fd_sc_hd__clkbuf_1 _4208_ (.A(_1215_),
    .X(_0083_));
 sky130_fd_sc_hd__mux2_1 _4209_ (.A0(net49),
    .A1(\core_1.fetch.out_buffer_data_instr[1] ),
    .S(_1214_),
    .X(_1216_));
 sky130_fd_sc_hd__clkbuf_1 _4210_ (.A(_1216_),
    .X(_0084_));
 sky130_fd_sc_hd__mux2_1 _4211_ (.A0(net60),
    .A1(\core_1.fetch.out_buffer_data_instr[2] ),
    .S(_1214_),
    .X(_1217_));
 sky130_fd_sc_hd__clkbuf_1 _4212_ (.A(_1217_),
    .X(_0085_));
 sky130_fd_sc_hd__mux2_1 _4213_ (.A0(net63),
    .A1(\core_1.fetch.out_buffer_data_instr[3] ),
    .S(_1214_),
    .X(_1218_));
 sky130_fd_sc_hd__clkbuf_1 _4214_ (.A(_1218_),
    .X(_0086_));
 sky130_fd_sc_hd__mux2_1 _4215_ (.A0(net64),
    .A1(\core_1.fetch.out_buffer_data_instr[4] ),
    .S(_1214_),
    .X(_1219_));
 sky130_fd_sc_hd__clkbuf_1 _4216_ (.A(_1219_),
    .X(_0087_));
 sky130_fd_sc_hd__mux2_1 _4217_ (.A0(net65),
    .A1(\core_1.fetch.out_buffer_data_instr[5] ),
    .S(_1214_),
    .X(_1220_));
 sky130_fd_sc_hd__clkbuf_1 _4218_ (.A(_1220_),
    .X(_0088_));
 sky130_fd_sc_hd__mux2_1 _4219_ (.A0(net66),
    .A1(\core_1.fetch.out_buffer_data_instr[6] ),
    .S(_1214_),
    .X(_1221_));
 sky130_fd_sc_hd__clkbuf_1 _4220_ (.A(_1221_),
    .X(_0089_));
 sky130_fd_sc_hd__mux2_1 _4221_ (.A0(net67),
    .A1(\core_1.fetch.out_buffer_data_instr[7] ),
    .S(_1214_),
    .X(_1222_));
 sky130_fd_sc_hd__clkbuf_1 _4222_ (.A(_1222_),
    .X(_0090_));
 sky130_fd_sc_hd__mux2_1 _4223_ (.A0(net68),
    .A1(\core_1.fetch.out_buffer_data_instr[8] ),
    .S(_1214_),
    .X(_1223_));
 sky130_fd_sc_hd__clkbuf_1 _4224_ (.A(_1223_),
    .X(_0091_));
 sky130_fd_sc_hd__mux2_1 _4225_ (.A0(net69),
    .A1(\core_1.fetch.out_buffer_data_instr[9] ),
    .S(_1214_),
    .X(_1224_));
 sky130_fd_sc_hd__clkbuf_1 _4226_ (.A(_1224_),
    .X(_0092_));
 sky130_fd_sc_hd__clkbuf_8 _4227_ (.A(_1213_),
    .X(_1225_));
 sky130_fd_sc_hd__mux2_1 _4228_ (.A0(net39),
    .A1(\core_1.fetch.out_buffer_data_instr[10] ),
    .S(_1225_),
    .X(_1226_));
 sky130_fd_sc_hd__clkbuf_1 _4229_ (.A(_1226_),
    .X(_0093_));
 sky130_fd_sc_hd__mux2_1 _4230_ (.A0(net40),
    .A1(\core_1.fetch.out_buffer_data_instr[11] ),
    .S(_1225_),
    .X(_1227_));
 sky130_fd_sc_hd__clkbuf_1 _4231_ (.A(_1227_),
    .X(_0094_));
 sky130_fd_sc_hd__mux2_1 _4232_ (.A0(net41),
    .A1(\core_1.fetch.out_buffer_data_instr[12] ),
    .S(_1225_),
    .X(_1228_));
 sky130_fd_sc_hd__clkbuf_1 _4233_ (.A(_1228_),
    .X(_0095_));
 sky130_fd_sc_hd__mux2_1 _4234_ (.A0(net42),
    .A1(\core_1.fetch.out_buffer_data_instr[13] ),
    .S(_1225_),
    .X(_1229_));
 sky130_fd_sc_hd__clkbuf_1 _4235_ (.A(_1229_),
    .X(_0096_));
 sky130_fd_sc_hd__mux2_1 _4236_ (.A0(net43),
    .A1(\core_1.fetch.out_buffer_data_instr[14] ),
    .S(_1225_),
    .X(_1230_));
 sky130_fd_sc_hd__clkbuf_1 _4237_ (.A(_1230_),
    .X(_0097_));
 sky130_fd_sc_hd__mux2_1 _4238_ (.A0(net44),
    .A1(\core_1.fetch.out_buffer_data_instr[15] ),
    .S(_1225_),
    .X(_1231_));
 sky130_fd_sc_hd__clkbuf_1 _4239_ (.A(_1231_),
    .X(_0098_));
 sky130_fd_sc_hd__mux2_1 _4240_ (.A0(net45),
    .A1(\core_1.fetch.out_buffer_data_instr[16] ),
    .S(_1225_),
    .X(_1232_));
 sky130_fd_sc_hd__clkbuf_1 _4241_ (.A(_1232_),
    .X(_0099_));
 sky130_fd_sc_hd__mux2_1 _4242_ (.A0(net46),
    .A1(\core_1.fetch.out_buffer_data_instr[17] ),
    .S(_1225_),
    .X(_1233_));
 sky130_fd_sc_hd__clkbuf_1 _4243_ (.A(_1233_),
    .X(_0100_));
 sky130_fd_sc_hd__mux2_1 _4244_ (.A0(net47),
    .A1(\core_1.fetch.out_buffer_data_instr[18] ),
    .S(_1225_),
    .X(_1234_));
 sky130_fd_sc_hd__clkbuf_1 _4245_ (.A(_1234_),
    .X(_0101_));
 sky130_fd_sc_hd__mux2_1 _4246_ (.A0(net48),
    .A1(\core_1.fetch.out_buffer_data_instr[19] ),
    .S(_1225_),
    .X(_1235_));
 sky130_fd_sc_hd__clkbuf_1 _4247_ (.A(_1235_),
    .X(_0102_));
 sky130_fd_sc_hd__buf_4 _4248_ (.A(_1213_),
    .X(_1236_));
 sky130_fd_sc_hd__mux2_1 _4249_ (.A0(net50),
    .A1(\core_1.fetch.out_buffer_data_instr[20] ),
    .S(_1236_),
    .X(_1237_));
 sky130_fd_sc_hd__clkbuf_1 _4250_ (.A(_1237_),
    .X(_0103_));
 sky130_fd_sc_hd__mux2_1 _4251_ (.A0(net51),
    .A1(\core_1.fetch.out_buffer_data_instr[21] ),
    .S(_1236_),
    .X(_1238_));
 sky130_fd_sc_hd__clkbuf_1 _4252_ (.A(_1238_),
    .X(_0104_));
 sky130_fd_sc_hd__mux2_1 _4253_ (.A0(net52),
    .A1(\core_1.fetch.out_buffer_data_instr[22] ),
    .S(_1236_),
    .X(_1239_));
 sky130_fd_sc_hd__clkbuf_1 _4254_ (.A(_1239_),
    .X(_0105_));
 sky130_fd_sc_hd__mux2_1 _4255_ (.A0(net53),
    .A1(\core_1.fetch.out_buffer_data_instr[23] ),
    .S(_1236_),
    .X(_1240_));
 sky130_fd_sc_hd__clkbuf_1 _4256_ (.A(_1240_),
    .X(_0106_));
 sky130_fd_sc_hd__mux2_1 _4257_ (.A0(net54),
    .A1(\core_1.fetch.out_buffer_data_instr[24] ),
    .S(_1236_),
    .X(_1241_));
 sky130_fd_sc_hd__clkbuf_1 _4258_ (.A(_1241_),
    .X(_0107_));
 sky130_fd_sc_hd__mux2_1 _4259_ (.A0(net55),
    .A1(\core_1.fetch.out_buffer_data_instr[25] ),
    .S(_1236_),
    .X(_1242_));
 sky130_fd_sc_hd__clkbuf_1 _4260_ (.A(_1242_),
    .X(_0108_));
 sky130_fd_sc_hd__mux2_1 _4261_ (.A0(net56),
    .A1(\core_1.fetch.out_buffer_data_instr[26] ),
    .S(_1236_),
    .X(_1243_));
 sky130_fd_sc_hd__clkbuf_1 _4262_ (.A(_1243_),
    .X(_0109_));
 sky130_fd_sc_hd__mux2_1 _4263_ (.A0(net57),
    .A1(\core_1.fetch.out_buffer_data_instr[27] ),
    .S(_1236_),
    .X(_1244_));
 sky130_fd_sc_hd__clkbuf_1 _4264_ (.A(_1244_),
    .X(_0110_));
 sky130_fd_sc_hd__mux2_1 _4265_ (.A0(net58),
    .A1(\core_1.fetch.out_buffer_data_instr[28] ),
    .S(_1236_),
    .X(_1245_));
 sky130_fd_sc_hd__clkbuf_1 _4266_ (.A(_1245_),
    .X(_0111_));
 sky130_fd_sc_hd__mux2_1 _4267_ (.A0(net59),
    .A1(\core_1.fetch.out_buffer_data_instr[29] ),
    .S(_1236_),
    .X(_1246_));
 sky130_fd_sc_hd__clkbuf_1 _4268_ (.A(_1246_),
    .X(_0112_));
 sky130_fd_sc_hd__mux2_1 _4269_ (.A0(net61),
    .A1(\core_1.fetch.out_buffer_data_instr[30] ),
    .S(_1213_),
    .X(_1247_));
 sky130_fd_sc_hd__clkbuf_1 _4270_ (.A(_1247_),
    .X(_0113_));
 sky130_fd_sc_hd__mux2_1 _4271_ (.A0(net62),
    .A1(\core_1.fetch.out_buffer_data_instr[31] ),
    .S(_1213_),
    .X(_1248_));
 sky130_fd_sc_hd__clkbuf_1 _4272_ (.A(_1248_),
    .X(_0114_));
 sky130_fd_sc_hd__a21oi_1 _4273_ (.A1(net70),
    .A2(_1026_),
    .B1(_0666_),
    .Y(_1249_));
 sky130_fd_sc_hd__nor4_1 _4274_ (.A(_0785_),
    .B(_1122_),
    .C(_0739_),
    .D(_1249_),
    .Y(_0115_));
 sky130_fd_sc_hd__nor2_1 _4275_ (.A(_0811_),
    .B(_1121_),
    .Y(_1250_));
 sky130_fd_sc_hd__mux2_1 _4276_ (.A0(_1250_),
    .A1(net161),
    .S(_0784_),
    .X(_1251_));
 sky130_fd_sc_hd__clkbuf_1 _4277_ (.A(_1251_),
    .X(_0116_));
 sky130_fd_sc_hd__or3_1 _4278_ (.A(_0813_),
    .B(_1121_),
    .C(_0782_),
    .X(_1252_));
 sky130_fd_sc_hd__a21bo_1 _4279_ (.A1(net177),
    .A2(net168),
    .B1_N(_1252_),
    .X(_0117_));
 sky130_fd_sc_hd__or3b_1 _4280_ (.A(_1121_),
    .B(_0782_),
    .C_N(\core_1.fetch.prev_request_pc[2] ),
    .X(_1253_));
 sky130_fd_sc_hd__a21bo_1 _4281_ (.A1(net177),
    .A2(net169),
    .B1_N(_1253_),
    .X(_0118_));
 sky130_fd_sc_hd__and2_1 _4282_ (.A(\core_1.fetch.prev_request_pc[3] ),
    .B(_0662_),
    .X(_1254_));
 sky130_fd_sc_hd__mux2_1 _4283_ (.A0(_1254_),
    .A1(net170),
    .S(_0784_),
    .X(_1255_));
 sky130_fd_sc_hd__clkbuf_1 _4284_ (.A(_1255_),
    .X(_0119_));
 sky130_fd_sc_hd__or3_1 _4285_ (.A(_0822_),
    .B(_1121_),
    .C(_0782_),
    .X(_1256_));
 sky130_fd_sc_hd__a21bo_1 _4286_ (.A1(net177),
    .A2(net171),
    .B1_N(_1256_),
    .X(_0120_));
 sky130_fd_sc_hd__or3_1 _4287_ (.A(_0819_),
    .B(_1121_),
    .C(_0782_),
    .X(_1257_));
 sky130_fd_sc_hd__a21bo_1 _4288_ (.A1(net177),
    .A2(net172),
    .B1_N(_1257_),
    .X(_0121_));
 sky130_fd_sc_hd__nor2_1 _4289_ (.A(_0818_),
    .B(_1121_),
    .Y(_1258_));
 sky130_fd_sc_hd__mux2_1 _4290_ (.A0(_1258_),
    .A1(net173),
    .S(_0784_),
    .X(_1259_));
 sky130_fd_sc_hd__clkbuf_1 _4291_ (.A(_1259_),
    .X(_0122_));
 sky130_fd_sc_hd__nor2_1 _4292_ (.A(_0809_),
    .B(_1121_),
    .Y(_1260_));
 sky130_fd_sc_hd__mux2_1 _4293_ (.A0(_1260_),
    .A1(net174),
    .S(_0784_),
    .X(_1261_));
 sky130_fd_sc_hd__clkbuf_1 _4294_ (.A(_1261_),
    .X(_0123_));
 sky130_fd_sc_hd__nor2_4 _4295_ (.A(net71),
    .B(_0782_),
    .Y(_1262_));
 sky130_fd_sc_hd__a22o_1 _4296_ (.A1(net177),
    .A2(net175),
    .B1(_1262_),
    .B2(\core_1.fetch.prev_request_pc[8] ),
    .X(_0124_));
 sky130_fd_sc_hd__a22o_1 _4297_ (.A1(net177),
    .A2(net176),
    .B1(_1262_),
    .B2(\core_1.fetch.prev_request_pc[9] ),
    .X(_0125_));
 sky130_fd_sc_hd__a22o_1 _4298_ (.A1(net177),
    .A2(net162),
    .B1(_1262_),
    .B2(\core_1.fetch.prev_request_pc[10] ),
    .X(_0126_));
 sky130_fd_sc_hd__a22o_1 _4299_ (.A1(net177),
    .A2(net163),
    .B1(_1262_),
    .B2(\core_1.fetch.prev_request_pc[11] ),
    .X(_0127_));
 sky130_fd_sc_hd__a22o_1 _4300_ (.A1(_0784_),
    .A2(net164),
    .B1(_1262_),
    .B2(\core_1.fetch.prev_request_pc[12] ),
    .X(_0128_));
 sky130_fd_sc_hd__a22o_1 _4301_ (.A1(_0784_),
    .A2(net165),
    .B1(_1262_),
    .B2(\core_1.fetch.prev_request_pc[13] ),
    .X(_0129_));
 sky130_fd_sc_hd__a22o_1 _4302_ (.A1(_0784_),
    .A2(net166),
    .B1(_1262_),
    .B2(\core_1.fetch.prev_request_pc[14] ),
    .X(_0130_));
 sky130_fd_sc_hd__a22o_1 _4303_ (.A1(_0784_),
    .A2(net167),
    .B1(_1262_),
    .B2(\core_1.fetch.prev_request_pc[15] ),
    .X(_0131_));
 sky130_fd_sc_hd__mux2_1 _4304_ (.A0(\core_1.fetch.current_req_branch_pred ),
    .A1(\core_1.fetch.out_buffer_data_pred ),
    .S(_1213_),
    .X(_1263_));
 sky130_fd_sc_hd__clkbuf_1 _4305_ (.A(_1263_),
    .X(_0132_));
 sky130_fd_sc_hd__buf_4 _4306_ (.A(_1027_),
    .X(_1264_));
 sky130_fd_sc_hd__mux2_1 _4307_ (.A0(_0742_),
    .A1(\core_1.decode.i_instr_l[0] ),
    .S(_1264_),
    .X(_1265_));
 sky130_fd_sc_hd__clkbuf_1 _4308_ (.A(_1265_),
    .X(_0133_));
 sky130_fd_sc_hd__mux2_1 _4309_ (.A0(_0743_),
    .A1(\core_1.decode.i_instr_l[1] ),
    .S(_1264_),
    .X(_1266_));
 sky130_fd_sc_hd__clkbuf_1 _4310_ (.A(_1266_),
    .X(_0134_));
 sky130_fd_sc_hd__mux2_1 _4311_ (.A0(_0745_),
    .A1(\core_1.decode.i_instr_l[2] ),
    .S(_1264_),
    .X(_1267_));
 sky130_fd_sc_hd__clkbuf_1 _4312_ (.A(_1267_),
    .X(_0135_));
 sky130_fd_sc_hd__mux2_1 _4313_ (.A0(_0746_),
    .A1(\core_1.decode.i_instr_l[3] ),
    .S(_1264_),
    .X(_1268_));
 sky130_fd_sc_hd__clkbuf_1 _4314_ (.A(_1268_),
    .X(_0136_));
 sky130_fd_sc_hd__mux2_1 _4315_ (.A0(_0779_),
    .A1(\core_1.decode.i_instr_l[4] ),
    .S(_1264_),
    .X(_1269_));
 sky130_fd_sc_hd__clkbuf_1 _4316_ (.A(_1269_),
    .X(_0137_));
 sky130_fd_sc_hd__mux2_1 _4317_ (.A0(_0741_),
    .A1(\core_1.decode.i_instr_l[5] ),
    .S(_1264_),
    .X(_1270_));
 sky130_fd_sc_hd__clkbuf_1 _4318_ (.A(_1270_),
    .X(_0138_));
 sky130_fd_sc_hd__mux2_1 _4319_ (.A0(_0740_),
    .A1(\core_1.decode.i_instr_l[6] ),
    .S(_1264_),
    .X(_1271_));
 sky130_fd_sc_hd__clkbuf_1 _4320_ (.A(_1271_),
    .X(_0139_));
 sky130_fd_sc_hd__mux2_1 _4321_ (.A0(_0840_),
    .A1(\core_1.decode.i_instr_l[7] ),
    .S(_1264_),
    .X(_1272_));
 sky130_fd_sc_hd__clkbuf_1 _4322_ (.A(_1272_),
    .X(_0140_));
 sky130_fd_sc_hd__mux2_1 _4323_ (.A0(_0839_),
    .A1(\core_1.decode.i_instr_l[8] ),
    .S(_1264_),
    .X(_1273_));
 sky130_fd_sc_hd__clkbuf_1 _4324_ (.A(_1273_),
    .X(_0141_));
 sky130_fd_sc_hd__mux2_1 _4325_ (.A0(_0842_),
    .A1(\core_1.decode.i_instr_l[9] ),
    .S(_1264_),
    .X(_1274_));
 sky130_fd_sc_hd__clkbuf_1 _4326_ (.A(_1274_),
    .X(_0142_));
 sky130_fd_sc_hd__buf_4 _4327_ (.A(_1027_),
    .X(_1275_));
 sky130_fd_sc_hd__mux2_1 _4328_ (.A0(_0841_),
    .A1(\core_1.decode.i_instr_l[10] ),
    .S(_1275_),
    .X(_1276_));
 sky130_fd_sc_hd__clkbuf_1 _4329_ (.A(_1276_),
    .X(_0143_));
 sky130_fd_sc_hd__mux2_1 _4330_ (.A0(net40),
    .A1(\core_1.fetch.out_buffer_data_instr[11] ),
    .S(_0666_),
    .X(_1277_));
 sky130_fd_sc_hd__mux2_1 _4331_ (.A0(_1277_),
    .A1(\core_1.decode.i_instr_l[11] ),
    .S(_1275_),
    .X(_1278_));
 sky130_fd_sc_hd__clkbuf_1 _4332_ (.A(_1278_),
    .X(_0144_));
 sky130_fd_sc_hd__mux2_1 _4333_ (.A0(net41),
    .A1(\core_1.fetch.out_buffer_data_instr[12] ),
    .S(_0666_),
    .X(_1279_));
 sky130_fd_sc_hd__mux2_1 _4334_ (.A0(_1279_),
    .A1(\core_1.decode.i_instr_l[12] ),
    .S(_1275_),
    .X(_1280_));
 sky130_fd_sc_hd__clkbuf_1 _4335_ (.A(_1280_),
    .X(_0145_));
 sky130_fd_sc_hd__mux2_1 _4336_ (.A0(net42),
    .A1(\core_1.fetch.out_buffer_data_instr[13] ),
    .S(_0666_),
    .X(_1281_));
 sky130_fd_sc_hd__mux2_1 _4337_ (.A0(_1281_),
    .A1(\core_1.decode.i_instr_l[13] ),
    .S(_1275_),
    .X(_1282_));
 sky130_fd_sc_hd__clkbuf_1 _4338_ (.A(_1282_),
    .X(_0146_));
 sky130_fd_sc_hd__mux2_1 _4339_ (.A0(net43),
    .A1(\core_1.fetch.out_buffer_data_instr[14] ),
    .S(_0666_),
    .X(_1283_));
 sky130_fd_sc_hd__mux2_1 _4340_ (.A0(_1283_),
    .A1(\core_1.decode.i_instr_l[14] ),
    .S(_1275_),
    .X(_1284_));
 sky130_fd_sc_hd__clkbuf_1 _4341_ (.A(_1284_),
    .X(_0147_));
 sky130_fd_sc_hd__mux2_1 _4342_ (.A0(net44),
    .A1(\core_1.fetch.out_buffer_data_instr[15] ),
    .S(_0666_),
    .X(_1285_));
 sky130_fd_sc_hd__mux2_1 _4343_ (.A0(_1285_),
    .A1(\core_1.decode.i_instr_l[15] ),
    .S(_1275_),
    .X(_1286_));
 sky130_fd_sc_hd__clkbuf_1 _4344_ (.A(_1286_),
    .X(_0148_));
 sky130_fd_sc_hd__mux2_1 _4345_ (.A0(_0763_),
    .A1(\core_1.decode.i_imm_pass[0] ),
    .S(_1275_),
    .X(_1287_));
 sky130_fd_sc_hd__clkbuf_1 _4346_ (.A(_1287_),
    .X(_0149_));
 sky130_fd_sc_hd__mux2_1 _4347_ (.A0(_0751_),
    .A1(\core_1.decode.i_imm_pass[1] ),
    .S(_1275_),
    .X(_1288_));
 sky130_fd_sc_hd__clkbuf_1 _4348_ (.A(_1288_),
    .X(_0150_));
 sky130_fd_sc_hd__mux2_1 _4349_ (.A0(_0758_),
    .A1(\core_1.decode.i_imm_pass[2] ),
    .S(_1275_),
    .X(_1289_));
 sky130_fd_sc_hd__clkbuf_1 _4350_ (.A(_1289_),
    .X(_0151_));
 sky130_fd_sc_hd__mux2_1 _4351_ (.A0(_0754_),
    .A1(\core_1.decode.i_imm_pass[3] ),
    .S(_1275_),
    .X(_1290_));
 sky130_fd_sc_hd__clkbuf_1 _4352_ (.A(_1290_),
    .X(_0152_));
 sky130_fd_sc_hd__clkbuf_4 _4353_ (.A(_1027_),
    .X(_1291_));
 sky130_fd_sc_hd__mux2_1 _4354_ (.A0(_0759_),
    .A1(\core_1.decode.i_imm_pass[4] ),
    .S(_1291_),
    .X(_1292_));
 sky130_fd_sc_hd__clkbuf_1 _4355_ (.A(_1292_),
    .X(_0153_));
 sky130_fd_sc_hd__mux2_1 _4356_ (.A0(_0762_),
    .A1(\core_1.decode.i_imm_pass[5] ),
    .S(_1291_),
    .X(_1293_));
 sky130_fd_sc_hd__clkbuf_1 _4357_ (.A(_1293_),
    .X(_0154_));
 sky130_fd_sc_hd__mux2_1 _4358_ (.A0(_0769_),
    .A1(\core_1.decode.i_imm_pass[6] ),
    .S(_1291_),
    .X(_1294_));
 sky130_fd_sc_hd__clkbuf_1 _4359_ (.A(_1294_),
    .X(_0155_));
 sky130_fd_sc_hd__mux2_1 _4360_ (.A0(_0756_),
    .A1(\core_1.decode.i_imm_pass[7] ),
    .S(_1291_),
    .X(_1295_));
 sky130_fd_sc_hd__clkbuf_1 _4361_ (.A(_1295_),
    .X(_0156_));
 sky130_fd_sc_hd__mux2_1 _4362_ (.A0(_0749_),
    .A1(\core_1.decode.i_imm_pass[8] ),
    .S(_1291_),
    .X(_1296_));
 sky130_fd_sc_hd__clkbuf_1 _4363_ (.A(_1296_),
    .X(_0157_));
 sky130_fd_sc_hd__mux2_1 _4364_ (.A0(_0772_),
    .A1(\core_1.decode.i_imm_pass[9] ),
    .S(_1291_),
    .X(_1297_));
 sky130_fd_sc_hd__clkbuf_1 _4365_ (.A(_1297_),
    .X(_0158_));
 sky130_fd_sc_hd__mux2_1 _4366_ (.A0(_0750_),
    .A1(\core_1.decode.i_imm_pass[10] ),
    .S(_1291_),
    .X(_1298_));
 sky130_fd_sc_hd__clkbuf_1 _4367_ (.A(_1298_),
    .X(_0159_));
 sky130_fd_sc_hd__mux2_1 _4368_ (.A0(_0770_),
    .A1(\core_1.decode.i_imm_pass[11] ),
    .S(_1291_),
    .X(_1299_));
 sky130_fd_sc_hd__clkbuf_1 _4369_ (.A(_1299_),
    .X(_0160_));
 sky130_fd_sc_hd__mux2_1 _4370_ (.A0(_0765_),
    .A1(\core_1.decode.i_imm_pass[12] ),
    .S(_1291_),
    .X(_1300_));
 sky130_fd_sc_hd__clkbuf_1 _4371_ (.A(_1300_),
    .X(_0161_));
 sky130_fd_sc_hd__mux2_1 _4372_ (.A0(_0773_),
    .A1(\core_1.decode.i_imm_pass[13] ),
    .S(_1291_),
    .X(_1301_));
 sky130_fd_sc_hd__clkbuf_1 _4373_ (.A(_1301_),
    .X(_0162_));
 sky130_fd_sc_hd__mux2_1 _4374_ (.A0(_0760_),
    .A1(\core_1.decode.i_imm_pass[14] ),
    .S(_1027_),
    .X(_1302_));
 sky130_fd_sc_hd__clkbuf_1 _4375_ (.A(_1302_),
    .X(_0163_));
 sky130_fd_sc_hd__mux2_1 _4376_ (.A0(_0767_),
    .A1(\core_1.decode.i_imm_pass[15] ),
    .S(_1027_),
    .X(_1303_));
 sky130_fd_sc_hd__clkbuf_1 _4377_ (.A(_1303_),
    .X(_0164_));
 sky130_fd_sc_hd__nor2_1 _4378_ (.A(_1122_),
    .B(net70),
    .Y(_1304_));
 sky130_fd_sc_hd__a21o_1 _4379_ (.A1(\core_1.fetch.dbg_out ),
    .A2(_1304_),
    .B1(net177),
    .X(_0165_));
 sky130_fd_sc_hd__o211a_1 _4380_ (.A1(\core_1.fetch.flush_event_invalidate ),
    .A2(\core_1.fetch.dbg_out ),
    .B1(_1211_),
    .C1(_1304_),
    .X(_0166_));
 sky130_fd_sc_hd__and2_1 _4381_ (.A(_0850_),
    .B(_1262_),
    .X(_1305_));
 sky130_fd_sc_hd__clkbuf_1 _4382_ (.A(_1305_),
    .X(_0167_));
 sky130_fd_sc_hd__clkbuf_1 _4383_ (.A(_1122_),
    .X(_1306_));
 sky130_fd_sc_hd__clkbuf_1 _4384_ (.A(_1306_),
    .X(_0168_));
 sky130_fd_sc_hd__buf_6 _4385_ (.A(_0662_),
    .X(_1307_));
 sky130_fd_sc_hd__clkinv_2 _4386_ (.A(net37),
    .Y(_1308_));
 sky130_fd_sc_hd__clkbuf_4 _4387_ (.A(\core_1.ew_mem_access ),
    .X(_1309_));
 sky130_fd_sc_hd__clkbuf_8 _4388_ (.A(_1309_),
    .X(_1310_));
 sky130_fd_sc_hd__mux2_1 _4389_ (.A0(_1308_),
    .A1(_1310_),
    .S(\core_1.ew_submit ),
    .X(_1311_));
 sky130_fd_sc_hd__and3_1 _4390_ (.A(_1307_),
    .B(_0731_),
    .C(_1311_),
    .X(_1312_));
 sky130_fd_sc_hd__clkbuf_1 _4391_ (.A(_1312_),
    .X(_0169_));
 sky130_fd_sc_hd__mux2_2 _4392_ (.A0(\core_1.fetch.current_req_branch_pred ),
    .A1(\core_1.fetch.out_buffer_data_pred ),
    .S(_0666_),
    .X(_1313_));
 sky130_fd_sc_hd__mux2_1 _4393_ (.A0(\core_1.decode.i_jmp_pred_pass ),
    .A1(_1313_),
    .S(\core_1.fetch.submitable ),
    .X(_1314_));
 sky130_fd_sc_hd__clkbuf_1 _4394_ (.A(_1314_),
    .X(_0170_));
 sky130_fd_sc_hd__inv_4 _4395_ (.A(\core_1.dec_r_bus_imm ),
    .Y(_1315_));
 sky130_fd_sc_hd__o221a_4 _4396_ (.A1(net94),
    .A2(_0520_),
    .B1(_0531_),
    .B2(_0544_),
    .C1(_1315_),
    .X(_1316_));
 sky130_fd_sc_hd__a21oi_4 _4397_ (.A1(_1077_),
    .A2(net184),
    .B1(_1316_),
    .Y(_1317_));
 sky130_fd_sc_hd__or2_1 _4398_ (.A(\core_1.execute.alu_mul_div.div_cur[15] ),
    .B(_1317_),
    .X(_1318_));
 sky130_fd_sc_hd__and2_1 _4399_ (.A(\core_1.dec_r_bus_imm ),
    .B(net183),
    .X(_1319_));
 sky130_fd_sc_hd__buf_8 _4400_ (.A(_1315_),
    .X(_1320_));
 sky130_fd_sc_hd__o221a_2 _4401_ (.A1(net93),
    .A2(_0520_),
    .B1(_0548_),
    .B2(_0554_),
    .C1(_1320_),
    .X(_1321_));
 sky130_fd_sc_hd__or2_1 _4402_ (.A(_1319_),
    .B(_1321_),
    .X(_1322_));
 sky130_fd_sc_hd__buf_2 _4403_ (.A(_1322_),
    .X(_1323_));
 sky130_fd_sc_hd__inv_2 _4404_ (.A(_1323_),
    .Y(_1324_));
 sky130_fd_sc_hd__inv_2 _4405_ (.A(net182),
    .Y(_1325_));
 sky130_fd_sc_hd__mux2_4 _4406_ (.A0(_1325_),
    .A1(_0571_),
    .S(_1320_),
    .X(_1326_));
 sky130_fd_sc_hd__and2_1 _4407_ (.A(\core_1.execute.alu_mul_div.div_cur[13] ),
    .B(_1326_),
    .X(_1327_));
 sky130_fd_sc_hd__nand2_1 _4408_ (.A(_1076_),
    .B(net181),
    .Y(_1328_));
 sky130_fd_sc_hd__o21ai_4 _4409_ (.A1(_1076_),
    .A2(_0577_),
    .B1(_1328_),
    .Y(_1329_));
 sky130_fd_sc_hd__inv_2 _4410_ (.A(_1329_),
    .Y(_1330_));
 sky130_fd_sc_hd__and2_1 _4411_ (.A(\core_1.execute.alu_mul_div.div_cur[12] ),
    .B(_1330_),
    .X(_1331_));
 sky130_fd_sc_hd__nor2_1 _4412_ (.A(\core_1.execute.alu_mul_div.div_cur[12] ),
    .B(_1330_),
    .Y(_1332_));
 sky130_fd_sc_hd__nor2_1 _4413_ (.A(_1331_),
    .B(_1332_),
    .Y(_1333_));
 sky130_fd_sc_hd__o221a_4 _4414_ (.A1(net90),
    .A2(_0520_),
    .B1(_0581_),
    .B2(_0584_),
    .C1(_1320_),
    .X(_1334_));
 sky130_fd_sc_hd__a21oi_2 _4415_ (.A1(_1077_),
    .A2(net180),
    .B1(_1334_),
    .Y(_1335_));
 sky130_fd_sc_hd__or2_1 _4416_ (.A(\core_1.execute.alu_mul_div.div_cur[11] ),
    .B(_1335_),
    .X(_1336_));
 sky130_fd_sc_hd__and2_1 _4417_ (.A(\core_1.dec_r_bus_imm ),
    .B(net179),
    .X(_1337_));
 sky130_fd_sc_hd__o221a_2 _4418_ (.A1(net89),
    .A2(_0520_),
    .B1(_0589_),
    .B2(_0592_),
    .C1(_1320_),
    .X(_1338_));
 sky130_fd_sc_hd__or2_1 _4419_ (.A(_1337_),
    .B(_1338_),
    .X(_1339_));
 sky130_fd_sc_hd__clkbuf_4 _4420_ (.A(_1339_),
    .X(_1340_));
 sky130_fd_sc_hd__clkinv_2 _4421_ (.A(_1340_),
    .Y(_1341_));
 sky130_fd_sc_hd__nand2_1 _4422_ (.A(_1076_),
    .B(net193),
    .Y(_1342_));
 sky130_fd_sc_hd__o21ai_4 _4423_ (.A1(_1076_),
    .A2(_0600_),
    .B1(_1342_),
    .Y(_1343_));
 sky130_fd_sc_hd__and2b_1 _4424_ (.A_N(_1343_),
    .B(\core_1.execute.alu_mul_div.div_cur[9] ),
    .X(_1344_));
 sky130_fd_sc_hd__inv_2 _4425_ (.A(\core_1.execute.alu_mul_div.div_cur[8] ),
    .Y(_1345_));
 sky130_fd_sc_hd__mux2_1 _4426_ (.A0(net192),
    .A1(net208),
    .S(_1315_),
    .X(_1346_));
 sky130_fd_sc_hd__clkbuf_8 _4427_ (.A(_1346_),
    .X(_1347_));
 sky130_fd_sc_hd__nand2_1 _4428_ (.A(_1076_),
    .B(net191),
    .Y(_1348_));
 sky130_fd_sc_hd__o21a_4 _4429_ (.A1(_1077_),
    .A2(_0614_),
    .B1(_1348_),
    .X(_1349_));
 sky130_fd_sc_hd__or2_1 _4430_ (.A(\core_1.execute.alu_mul_div.div_cur[7] ),
    .B(_1349_),
    .X(_1350_));
 sky130_fd_sc_hd__mux2_4 _4431_ (.A0(net190),
    .A1(net206),
    .S(_1320_),
    .X(_1351_));
 sky130_fd_sc_hd__inv_2 _4432_ (.A(_1351_),
    .Y(_1352_));
 sky130_fd_sc_hd__and2_1 _4433_ (.A(\core_1.execute.alu_mul_div.div_cur[6] ),
    .B(_1352_),
    .X(_1353_));
 sky130_fd_sc_hd__nor2_1 _4434_ (.A(\core_1.execute.alu_mul_div.div_cur[6] ),
    .B(_1352_),
    .Y(_1354_));
 sky130_fd_sc_hd__nor2_1 _4435_ (.A(_1353_),
    .B(_1354_),
    .Y(_1355_));
 sky130_fd_sc_hd__nand2_1 _4436_ (.A(_1076_),
    .B(net189),
    .Y(_1356_));
 sky130_fd_sc_hd__o21a_4 _4437_ (.A1(_1076_),
    .A2(_0627_),
    .B1(_1356_),
    .X(_1357_));
 sky130_fd_sc_hd__or2_1 _4438_ (.A(\core_1.execute.alu_mul_div.div_cur[5] ),
    .B(_1357_),
    .X(_1358_));
 sky130_fd_sc_hd__inv_2 _4439_ (.A(\core_1.execute.alu_mul_div.div_cur[4] ),
    .Y(_1359_));
 sky130_fd_sc_hd__mux2_1 _4440_ (.A0(net188),
    .A1(net204),
    .S(_1315_),
    .X(_1360_));
 sky130_fd_sc_hd__buf_6 _4441_ (.A(_1360_),
    .X(_1361_));
 sky130_fd_sc_hd__nor2_1 _4442_ (.A(_1359_),
    .B(_1361_),
    .Y(_1362_));
 sky130_fd_sc_hd__inv_2 _4443_ (.A(net188),
    .Y(_1363_));
 sky130_fd_sc_hd__mux2_4 _4444_ (.A0(_1363_),
    .A1(_0633_),
    .S(_1320_),
    .X(_1364_));
 sky130_fd_sc_hd__nor2_1 _4445_ (.A(\core_1.execute.alu_mul_div.div_cur[4] ),
    .B(_1364_),
    .Y(_1365_));
 sky130_fd_sc_hd__nor2_1 _4446_ (.A(_1362_),
    .B(_1365_),
    .Y(_1366_));
 sky130_fd_sc_hd__or2_1 _4447_ (.A(_1320_),
    .B(net187),
    .X(_1367_));
 sky130_fd_sc_hd__o21ai_4 _4448_ (.A1(_1077_),
    .A2(net203),
    .B1(_1367_),
    .Y(_1368_));
 sky130_fd_sc_hd__buf_4 _4449_ (.A(_1368_),
    .X(_1369_));
 sky130_fd_sc_hd__or2_1 _4450_ (.A(\core_1.execute.alu_mul_div.div_cur[3] ),
    .B(_1369_),
    .X(_1370_));
 sky130_fd_sc_hd__mux2_1 _4451_ (.A0(net186),
    .A1(net202),
    .S(_1320_),
    .X(_1371_));
 sky130_fd_sc_hd__buf_6 _4452_ (.A(_1371_),
    .X(_1372_));
 sky130_fd_sc_hd__xnor2_1 _4453_ (.A(\core_1.execute.alu_mul_div.div_cur[2] ),
    .B(_1372_),
    .Y(_1373_));
 sky130_fd_sc_hd__nand2_4 _4454_ (.A(\core_1.dec_r_bus_imm ),
    .B(net185),
    .Y(_1374_));
 sky130_fd_sc_hd__o311ai_4 _4455_ (.A1(_0648_),
    .A2(_0649_),
    .A3(_0652_),
    .B1(_0653_),
    .C1(_1315_),
    .Y(_1375_));
 sky130_fd_sc_hd__a21o_1 _4456_ (.A1(_1374_),
    .A2(_1375_),
    .B1(\core_1.execute.alu_mul_div.div_cur[1] ),
    .X(_1376_));
 sky130_fd_sc_hd__nand2_8 _4457_ (.A(\core_1.dec_r_bus_imm ),
    .B(net178),
    .Y(_1377_));
 sky130_fd_sc_hd__o311ai_4 _4458_ (.A1(_0655_),
    .A2(_0656_),
    .A3(_0659_),
    .B1(_0660_),
    .C1(_1315_),
    .Y(_1378_));
 sky130_fd_sc_hd__a21o_1 _4459_ (.A1(_1377_),
    .A2(_1378_),
    .B1(\core_1.execute.alu_mul_div.div_cur[0] ),
    .X(_1379_));
 sky130_fd_sc_hd__and3_1 _4460_ (.A(\core_1.execute.alu_mul_div.div_cur[1] ),
    .B(_1374_),
    .C(_1375_),
    .X(_1380_));
 sky130_fd_sc_hd__a21o_1 _4461_ (.A1(_1376_),
    .A2(_1379_),
    .B1(_1380_),
    .X(_1381_));
 sky130_fd_sc_hd__and2_1 _4462_ (.A(\core_1.execute.alu_mul_div.div_cur[3] ),
    .B(_1369_),
    .X(_1382_));
 sky130_fd_sc_hd__mux2_2 _4463_ (.A0(_1050_),
    .A1(_0647_),
    .S(_1320_),
    .X(_1383_));
 sky130_fd_sc_hd__buf_6 _4464_ (.A(_1383_),
    .X(_1384_));
 sky130_fd_sc_hd__and2_1 _4465_ (.A(\core_1.execute.alu_mul_div.div_cur[2] ),
    .B(_1384_),
    .X(_1385_));
 sky130_fd_sc_hd__a211o_1 _4466_ (.A1(_1373_),
    .A2(_1381_),
    .B1(_1382_),
    .C1(_1385_),
    .X(_1386_));
 sky130_fd_sc_hd__and2_1 _4467_ (.A(\core_1.execute.alu_mul_div.div_cur[5] ),
    .B(_1357_),
    .X(_1387_));
 sky130_fd_sc_hd__a311o_1 _4468_ (.A1(_1366_),
    .A2(_1370_),
    .A3(_1386_),
    .B1(_1362_),
    .C1(_1387_),
    .X(_1388_));
 sky130_fd_sc_hd__and2_1 _4469_ (.A(\core_1.execute.alu_mul_div.div_cur[7] ),
    .B(_1349_),
    .X(_1389_));
 sky130_fd_sc_hd__a311o_1 _4470_ (.A1(_1355_),
    .A2(_1358_),
    .A3(_1388_),
    .B1(_1353_),
    .C1(_1389_),
    .X(_1390_));
 sky130_fd_sc_hd__xnor2_1 _4471_ (.A(\core_1.execute.alu_mul_div.div_cur[8] ),
    .B(_1347_),
    .Y(_1391_));
 sky130_fd_sc_hd__and3_1 _4472_ (.A(_1350_),
    .B(_1390_),
    .C(_1391_),
    .X(_1392_));
 sky130_fd_sc_hd__o21bai_2 _4473_ (.A1(_1345_),
    .A2(_1347_),
    .B1_N(_1392_),
    .Y(_1393_));
 sky130_fd_sc_hd__xnor2_1 _4474_ (.A(\core_1.execute.alu_mul_div.div_cur[10] ),
    .B(_1340_),
    .Y(_1394_));
 sky130_fd_sc_hd__or2b_1 _4475_ (.A(\core_1.execute.alu_mul_div.div_cur[9] ),
    .B_N(_1343_),
    .X(_1395_));
 sky130_fd_sc_hd__o211a_1 _4476_ (.A1(_1344_),
    .A2(_1393_),
    .B1(_1394_),
    .C1(_1395_),
    .X(_1396_));
 sky130_fd_sc_hd__a21o_1 _4477_ (.A1(\core_1.execute.alu_mul_div.div_cur[10] ),
    .A2(_1341_),
    .B1(_1396_),
    .X(_1397_));
 sky130_fd_sc_hd__nand2_1 _4478_ (.A(\core_1.execute.alu_mul_div.div_cur[11] ),
    .B(_1335_),
    .Y(_1398_));
 sky130_fd_sc_hd__a21bo_1 _4479_ (.A1(_1336_),
    .A2(_1397_),
    .B1_N(_1398_),
    .X(_1399_));
 sky130_fd_sc_hd__a21o_1 _4480_ (.A1(_1333_),
    .A2(_1399_),
    .B1(_1331_),
    .X(_1400_));
 sky130_fd_sc_hd__xnor2_1 _4481_ (.A(\core_1.execute.alu_mul_div.div_cur[14] ),
    .B(_1323_),
    .Y(_1401_));
 sky130_fd_sc_hd__or2_1 _4482_ (.A(\core_1.execute.alu_mul_div.div_cur[13] ),
    .B(_1326_),
    .X(_1402_));
 sky130_fd_sc_hd__o211a_1 _4483_ (.A1(_1327_),
    .A2(_1400_),
    .B1(_1401_),
    .C1(_1402_),
    .X(_1403_));
 sky130_fd_sc_hd__a21o_1 _4484_ (.A1(\core_1.execute.alu_mul_div.div_cur[14] ),
    .A2(_1324_),
    .B1(_1403_),
    .X(_1404_));
 sky130_fd_sc_hd__and2_1 _4485_ (.A(\core_1.execute.alu_mul_div.div_cur[15] ),
    .B(_1317_),
    .X(_1405_));
 sky130_fd_sc_hd__a21o_4 _4486_ (.A1(_1318_),
    .A2(_1404_),
    .B1(_1405_),
    .X(_1406_));
 sky130_fd_sc_hd__buf_2 _4487_ (.A(_0732_),
    .X(_1407_));
 sky130_fd_sc_hd__and2_1 _4488_ (.A(\core_1.execute.alu_mul_div.comp ),
    .B(_1407_),
    .X(_1408_));
 sky130_fd_sc_hd__o21a_2 _4489_ (.A1(_1208_),
    .A2(_1406_),
    .B1(_1408_),
    .X(_1409_));
 sky130_fd_sc_hd__clkbuf_4 _4490_ (.A(_1409_),
    .X(_1410_));
 sky130_fd_sc_hd__a21oi_2 _4491_ (.A1(_1318_),
    .A2(_1404_),
    .B1(_1405_),
    .Y(_1411_));
 sky130_fd_sc_hd__clkbuf_4 _4492_ (.A(_1411_),
    .X(_1412_));
 sky130_fd_sc_hd__o21ai_4 _4493_ (.A1(_1207_),
    .A2(_1406_),
    .B1(_1408_),
    .Y(_1413_));
 sky130_fd_sc_hd__clkbuf_4 _4494_ (.A(_1413_),
    .X(_1414_));
 sky130_fd_sc_hd__and2_2 _4495_ (.A(_1200_),
    .B(_1206_),
    .X(_1415_));
 sky130_fd_sc_hd__clkbuf_4 _4496_ (.A(_1415_),
    .X(_1416_));
 sky130_fd_sc_hd__and2_2 _4497_ (.A(_1377_),
    .B(_1378_),
    .X(_1417_));
 sky130_fd_sc_hd__buf_4 _4498_ (.A(_1417_),
    .X(_1418_));
 sky130_fd_sc_hd__clkbuf_8 _4499_ (.A(_1418_),
    .X(_1419_));
 sky130_fd_sc_hd__nand2_1 _4500_ (.A(\core_1.execute.alu_mul_div.div_cur[0] ),
    .B(_1419_),
    .Y(_1420_));
 sky130_fd_sc_hd__nand2_1 _4501_ (.A(_1379_),
    .B(_1420_),
    .Y(_1421_));
 sky130_fd_sc_hd__and2b_1 _4502_ (.A_N(_1380_),
    .B(_1376_),
    .X(_1422_));
 sky130_fd_sc_hd__xor2_1 _4503_ (.A(_1422_),
    .B(_1379_),
    .X(_1423_));
 sky130_fd_sc_hd__or2_1 _4504_ (.A(_1207_),
    .B(_1423_),
    .X(_1424_));
 sky130_fd_sc_hd__clkbuf_4 _4505_ (.A(_1406_),
    .X(_1425_));
 sky130_fd_sc_hd__o211a_1 _4506_ (.A1(_1416_),
    .A2(_1421_),
    .B1(_1424_),
    .C1(_1425_),
    .X(_1426_));
 sky130_fd_sc_hd__a211o_1 _4507_ (.A1(\core_1.execute.alu_mul_div.div_cur[0] ),
    .A2(_1412_),
    .B1(_1414_),
    .C1(_1426_),
    .X(_1427_));
 sky130_fd_sc_hd__buf_2 _4508_ (.A(_0733_),
    .X(_1428_));
 sky130_fd_sc_hd__clkbuf_4 _4509_ (.A(_1428_),
    .X(_1429_));
 sky130_fd_sc_hd__o211a_1 _4510_ (.A1(\core_1.execute.alu_mul_div.div_cur[1] ),
    .A2(_1410_),
    .B1(_1427_),
    .C1(_1429_),
    .X(_0171_));
 sky130_fd_sc_hd__and2_1 _4511_ (.A(_1373_),
    .B(_1381_),
    .X(_1430_));
 sky130_fd_sc_hd__nor2_1 _4512_ (.A(_1373_),
    .B(_1381_),
    .Y(_1431_));
 sky130_fd_sc_hd__nor2_1 _4513_ (.A(_1430_),
    .B(_1431_),
    .Y(_1432_));
 sky130_fd_sc_hd__mux2_1 _4514_ (.A0(_1423_),
    .A1(_1432_),
    .S(_1415_),
    .X(_1433_));
 sky130_fd_sc_hd__mux2_1 _4515_ (.A0(\core_1.execute.alu_mul_div.div_cur[1] ),
    .A1(_1433_),
    .S(_1406_),
    .X(_1434_));
 sky130_fd_sc_hd__or2_1 _4516_ (.A(_1413_),
    .B(_1434_),
    .X(_1435_));
 sky130_fd_sc_hd__o211a_1 _4517_ (.A1(\core_1.execute.alu_mul_div.div_cur[2] ),
    .A2(_1410_),
    .B1(_1435_),
    .C1(_1429_),
    .X(_0172_));
 sky130_fd_sc_hd__nor2_1 _4518_ (.A(\core_1.execute.alu_mul_div.div_cur[3] ),
    .B(_1369_),
    .Y(_1436_));
 sky130_fd_sc_hd__or4_1 _4519_ (.A(_1436_),
    .B(_1382_),
    .C(_1385_),
    .D(_1430_),
    .X(_1437_));
 sky130_fd_sc_hd__o22ai_1 _4520_ (.A1(_1436_),
    .A2(_1382_),
    .B1(_1385_),
    .B2(_1430_),
    .Y(_1438_));
 sky130_fd_sc_hd__nand2_1 _4521_ (.A(_1437_),
    .B(_1438_),
    .Y(_1439_));
 sky130_fd_sc_hd__or2_1 _4522_ (.A(_1415_),
    .B(_1432_),
    .X(_1440_));
 sky130_fd_sc_hd__o211a_1 _4523_ (.A1(_1208_),
    .A2(_1439_),
    .B1(_1440_),
    .C1(_1425_),
    .X(_1441_));
 sky130_fd_sc_hd__a211o_1 _4524_ (.A1(\core_1.execute.alu_mul_div.div_cur[2] ),
    .A2(_1412_),
    .B1(_1414_),
    .C1(_1441_),
    .X(_1442_));
 sky130_fd_sc_hd__o211a_1 _4525_ (.A1(\core_1.execute.alu_mul_div.div_cur[3] ),
    .A2(_1410_),
    .B1(_1442_),
    .C1(_1429_),
    .X(_0173_));
 sky130_fd_sc_hd__nand2_1 _4526_ (.A(_1370_),
    .B(_1386_),
    .Y(_1443_));
 sky130_fd_sc_hd__xnor2_1 _4527_ (.A(_1366_),
    .B(_1443_),
    .Y(_1444_));
 sky130_fd_sc_hd__or2_1 _4528_ (.A(_1207_),
    .B(_1444_),
    .X(_1445_));
 sky130_fd_sc_hd__o211a_1 _4529_ (.A1(_1416_),
    .A2(_1439_),
    .B1(_1445_),
    .C1(_1425_),
    .X(_1446_));
 sky130_fd_sc_hd__a211o_1 _4530_ (.A1(\core_1.execute.alu_mul_div.div_cur[3] ),
    .A2(_1412_),
    .B1(_1414_),
    .C1(_1446_),
    .X(_1447_));
 sky130_fd_sc_hd__o211a_1 _4531_ (.A1(\core_1.execute.alu_mul_div.div_cur[4] ),
    .A2(_1410_),
    .B1(_1447_),
    .C1(_1429_),
    .X(_0174_));
 sky130_fd_sc_hd__a31o_1 _4532_ (.A1(_1366_),
    .A2(_1370_),
    .A3(_1386_),
    .B1(_1362_),
    .X(_1448_));
 sky130_fd_sc_hd__and2b_1 _4533_ (.A_N(_1387_),
    .B(_1358_),
    .X(_1449_));
 sky130_fd_sc_hd__xor2_1 _4534_ (.A(_1448_),
    .B(_1449_),
    .X(_1450_));
 sky130_fd_sc_hd__or2_1 _4535_ (.A(_1415_),
    .B(_1444_),
    .X(_1451_));
 sky130_fd_sc_hd__o211a_1 _4536_ (.A1(_1208_),
    .A2(_1450_),
    .B1(_1451_),
    .C1(_1425_),
    .X(_1452_));
 sky130_fd_sc_hd__a211o_1 _4537_ (.A1(\core_1.execute.alu_mul_div.div_cur[4] ),
    .A2(_1412_),
    .B1(_1414_),
    .C1(_1452_),
    .X(_1453_));
 sky130_fd_sc_hd__o211a_1 _4538_ (.A1(\core_1.execute.alu_mul_div.div_cur[5] ),
    .A2(_1410_),
    .B1(_1453_),
    .C1(_1429_),
    .X(_0175_));
 sky130_fd_sc_hd__and3_1 _4539_ (.A(_1355_),
    .B(_1358_),
    .C(_1388_),
    .X(_1454_));
 sky130_fd_sc_hd__a21oi_1 _4540_ (.A1(_1358_),
    .A2(_1388_),
    .B1(_1355_),
    .Y(_1455_));
 sky130_fd_sc_hd__nor2_1 _4541_ (.A(_1454_),
    .B(_1455_),
    .Y(_1456_));
 sky130_fd_sc_hd__mux2_1 _4542_ (.A0(_1450_),
    .A1(_1456_),
    .S(_1415_),
    .X(_1457_));
 sky130_fd_sc_hd__mux2_1 _4543_ (.A0(\core_1.execute.alu_mul_div.div_cur[5] ),
    .A1(_1457_),
    .S(_1406_),
    .X(_1458_));
 sky130_fd_sc_hd__or2_1 _4544_ (.A(_1413_),
    .B(_1458_),
    .X(_1459_));
 sky130_fd_sc_hd__o211a_1 _4545_ (.A1(\core_1.execute.alu_mul_div.div_cur[6] ),
    .A2(_1410_),
    .B1(_1459_),
    .C1(_1429_),
    .X(_0176_));
 sky130_fd_sc_hd__or2_1 _4546_ (.A(_1353_),
    .B(_1454_),
    .X(_1460_));
 sky130_fd_sc_hd__nor2_1 _4547_ (.A(\core_1.execute.alu_mul_div.div_cur[7] ),
    .B(_1349_),
    .Y(_1461_));
 sky130_fd_sc_hd__nor2_1 _4548_ (.A(_1461_),
    .B(_1389_),
    .Y(_1462_));
 sky130_fd_sc_hd__xor2_1 _4549_ (.A(_1460_),
    .B(_1462_),
    .X(_1463_));
 sky130_fd_sc_hd__or2_1 _4550_ (.A(_1415_),
    .B(_1456_),
    .X(_1464_));
 sky130_fd_sc_hd__o211a_1 _4551_ (.A1(_1208_),
    .A2(_1463_),
    .B1(_1464_),
    .C1(_1425_),
    .X(_1465_));
 sky130_fd_sc_hd__a211o_1 _4552_ (.A1(\core_1.execute.alu_mul_div.div_cur[6] ),
    .A2(_1412_),
    .B1(_1414_),
    .C1(_1465_),
    .X(_1466_));
 sky130_fd_sc_hd__o211a_1 _4553_ (.A1(\core_1.execute.alu_mul_div.div_cur[7] ),
    .A2(_1410_),
    .B1(_1466_),
    .C1(_1429_),
    .X(_0177_));
 sky130_fd_sc_hd__a21oi_1 _4554_ (.A1(_1350_),
    .A2(_1390_),
    .B1(_1391_),
    .Y(_1467_));
 sky130_fd_sc_hd__nor2_1 _4555_ (.A(_1392_),
    .B(_1467_),
    .Y(_1468_));
 sky130_fd_sc_hd__or2_1 _4556_ (.A(_1207_),
    .B(_1468_),
    .X(_1469_));
 sky130_fd_sc_hd__o211a_1 _4557_ (.A1(_1416_),
    .A2(_1463_),
    .B1(_1469_),
    .C1(_1425_),
    .X(_1470_));
 sky130_fd_sc_hd__a211o_1 _4558_ (.A1(\core_1.execute.alu_mul_div.div_cur[7] ),
    .A2(_1412_),
    .B1(_1414_),
    .C1(_1470_),
    .X(_1471_));
 sky130_fd_sc_hd__o211a_1 _4559_ (.A1(\core_1.execute.alu_mul_div.div_cur[8] ),
    .A2(_1410_),
    .B1(_1471_),
    .C1(_1429_),
    .X(_0178_));
 sky130_fd_sc_hd__xor2_1 _4560_ (.A(\core_1.execute.alu_mul_div.div_cur[9] ),
    .B(_1343_),
    .X(_1472_));
 sky130_fd_sc_hd__xnor2_1 _4561_ (.A(_1393_),
    .B(_1472_),
    .Y(_1473_));
 sky130_fd_sc_hd__or2_1 _4562_ (.A(_1415_),
    .B(_1468_),
    .X(_1474_));
 sky130_fd_sc_hd__o211a_1 _4563_ (.A1(_1208_),
    .A2(_1473_),
    .B1(_1474_),
    .C1(_1425_),
    .X(_1475_));
 sky130_fd_sc_hd__a211o_1 _4564_ (.A1(\core_1.execute.alu_mul_div.div_cur[8] ),
    .A2(_1412_),
    .B1(_1414_),
    .C1(_1475_),
    .X(_1476_));
 sky130_fd_sc_hd__clkbuf_4 _4565_ (.A(_1428_),
    .X(_1477_));
 sky130_fd_sc_hd__o211a_1 _4566_ (.A1(\core_1.execute.alu_mul_div.div_cur[9] ),
    .A2(_1410_),
    .B1(_1476_),
    .C1(_1477_),
    .X(_0179_));
 sky130_fd_sc_hd__o21ai_1 _4567_ (.A1(_1344_),
    .A2(_1393_),
    .B1(_1395_),
    .Y(_1478_));
 sky130_fd_sc_hd__xnor2_1 _4568_ (.A(_1394_),
    .B(_1478_),
    .Y(_1479_));
 sky130_fd_sc_hd__or2_1 _4569_ (.A(_1207_),
    .B(_1479_),
    .X(_1480_));
 sky130_fd_sc_hd__o211a_1 _4570_ (.A1(_1416_),
    .A2(_1473_),
    .B1(_1480_),
    .C1(_1425_),
    .X(_1481_));
 sky130_fd_sc_hd__a211o_1 _4571_ (.A1(\core_1.execute.alu_mul_div.div_cur[9] ),
    .A2(_1412_),
    .B1(_1414_),
    .C1(_1481_),
    .X(_1482_));
 sky130_fd_sc_hd__o211a_1 _4572_ (.A1(\core_1.execute.alu_mul_div.div_cur[10] ),
    .A2(_1410_),
    .B1(_1482_),
    .C1(_1477_),
    .X(_0180_));
 sky130_fd_sc_hd__nand2_1 _4573_ (.A(_1398_),
    .B(_1336_),
    .Y(_1483_));
 sky130_fd_sc_hd__xor2_1 _4574_ (.A(_1397_),
    .B(_1483_),
    .X(_1484_));
 sky130_fd_sc_hd__nand2_1 _4575_ (.A(_1416_),
    .B(_1484_),
    .Y(_1485_));
 sky130_fd_sc_hd__o211a_1 _4576_ (.A1(_1416_),
    .A2(_1479_),
    .B1(_1485_),
    .C1(_1425_),
    .X(_1486_));
 sky130_fd_sc_hd__a211o_1 _4577_ (.A1(\core_1.execute.alu_mul_div.div_cur[10] ),
    .A2(_1412_),
    .B1(_1414_),
    .C1(_1486_),
    .X(_1487_));
 sky130_fd_sc_hd__o211a_1 _4578_ (.A1(\core_1.execute.alu_mul_div.div_cur[11] ),
    .A2(_1409_),
    .B1(_1487_),
    .C1(_1477_),
    .X(_0181_));
 sky130_fd_sc_hd__xor2_1 _4579_ (.A(_1333_),
    .B(_1399_),
    .X(_1488_));
 sky130_fd_sc_hd__nand2_1 _4580_ (.A(_1208_),
    .B(_1484_),
    .Y(_1489_));
 sky130_fd_sc_hd__o211a_1 _4581_ (.A1(_1208_),
    .A2(_1488_),
    .B1(_1489_),
    .C1(_1425_),
    .X(_1490_));
 sky130_fd_sc_hd__a211o_1 _4582_ (.A1(\core_1.execute.alu_mul_div.div_cur[11] ),
    .A2(_1412_),
    .B1(_1414_),
    .C1(_1490_),
    .X(_1491_));
 sky130_fd_sc_hd__o211a_1 _4583_ (.A1(\core_1.execute.alu_mul_div.div_cur[12] ),
    .A2(_1409_),
    .B1(_1491_),
    .C1(_1477_),
    .X(_0182_));
 sky130_fd_sc_hd__inv_2 _4584_ (.A(_1402_),
    .Y(_1492_));
 sky130_fd_sc_hd__nor2_1 _4585_ (.A(_1492_),
    .B(_1327_),
    .Y(_1493_));
 sky130_fd_sc_hd__xor2_1 _4586_ (.A(_1400_),
    .B(_1493_),
    .X(_1494_));
 sky130_fd_sc_hd__or2_1 _4587_ (.A(_1415_),
    .B(_1488_),
    .X(_1495_));
 sky130_fd_sc_hd__o211a_1 _4588_ (.A1(_1208_),
    .A2(_1494_),
    .B1(_1495_),
    .C1(_1406_),
    .X(_1496_));
 sky130_fd_sc_hd__a211o_1 _4589_ (.A1(\core_1.execute.alu_mul_div.div_cur[12] ),
    .A2(_1411_),
    .B1(_1413_),
    .C1(_1496_),
    .X(_1497_));
 sky130_fd_sc_hd__o211a_1 _4590_ (.A1(\core_1.execute.alu_mul_div.div_cur[13] ),
    .A2(_1409_),
    .B1(_1497_),
    .C1(_1477_),
    .X(_0183_));
 sky130_fd_sc_hd__o21a_1 _4591_ (.A1(_1327_),
    .A2(_1400_),
    .B1(_1402_),
    .X(_1498_));
 sky130_fd_sc_hd__nor2_1 _4592_ (.A(_1401_),
    .B(_1498_),
    .Y(_1499_));
 sky130_fd_sc_hd__nor2_1 _4593_ (.A(_1403_),
    .B(_1499_),
    .Y(_1500_));
 sky130_fd_sc_hd__or2_1 _4594_ (.A(_1207_),
    .B(_1500_),
    .X(_1501_));
 sky130_fd_sc_hd__o211a_1 _4595_ (.A1(_1416_),
    .A2(_1494_),
    .B1(_1501_),
    .C1(_1406_),
    .X(_1502_));
 sky130_fd_sc_hd__a211o_1 _4596_ (.A1(\core_1.execute.alu_mul_div.div_cur[13] ),
    .A2(_1411_),
    .B1(_1413_),
    .C1(_1502_),
    .X(_1503_));
 sky130_fd_sc_hd__o211a_1 _4597_ (.A1(\core_1.execute.alu_mul_div.div_cur[14] ),
    .A2(_1409_),
    .B1(_1503_),
    .C1(_1477_),
    .X(_0184_));
 sky130_fd_sc_hd__clkinv_2 _4598_ (.A(_1318_),
    .Y(_1504_));
 sky130_fd_sc_hd__or2_1 _4599_ (.A(_1504_),
    .B(_1405_),
    .X(_1505_));
 sky130_fd_sc_hd__xnor2_1 _4600_ (.A(_1404_),
    .B(_1505_),
    .Y(_1506_));
 sky130_fd_sc_hd__or2_1 _4601_ (.A(_1415_),
    .B(_1500_),
    .X(_1507_));
 sky130_fd_sc_hd__o211a_1 _4602_ (.A1(_1208_),
    .A2(_1506_),
    .B1(_1507_),
    .C1(_1406_),
    .X(_1508_));
 sky130_fd_sc_hd__a211o_1 _4603_ (.A1(\core_1.execute.alu_mul_div.div_cur[14] ),
    .A2(_1411_),
    .B1(_1413_),
    .C1(_1508_),
    .X(_1509_));
 sky130_fd_sc_hd__o211a_1 _4604_ (.A1(\core_1.execute.alu_mul_div.div_cur[15] ),
    .A2(_1409_),
    .B1(_1509_),
    .C1(_1477_),
    .X(_0185_));
 sky130_fd_sc_hd__and2_1 _4605_ (.A(\core_1.decode.o_submit ),
    .B(_1407_),
    .X(_1510_));
 sky130_fd_sc_hd__clkbuf_2 _4606_ (.A(_1510_),
    .X(_1511_));
 sky130_fd_sc_hd__or3_4 _4607_ (.A(_0705_),
    .B(_0709_),
    .C(\core_1.dec_l_reg_sel[0] ),
    .X(_1512_));
 sky130_fd_sc_hd__buf_6 _4608_ (.A(_1512_),
    .X(_1513_));
 sky130_fd_sc_hd__nor2_4 _4609_ (.A(_0701_),
    .B(_0721_),
    .Y(_1514_));
 sky130_fd_sc_hd__nor3b_4 _4610_ (.A(_0705_),
    .B(\core_1.dec_l_reg_sel[0] ),
    .C_N(_0709_),
    .Y(_1515_));
 sky130_fd_sc_hd__buf_4 _4611_ (.A(_1515_),
    .X(_1516_));
 sky130_fd_sc_hd__a22o_1 _4612_ (.A1(\core_1.execute.rf.reg_outputs[5][15] ),
    .A2(_1514_),
    .B1(_1516_),
    .B2(\core_1.execute.rf.reg_outputs[2][15] ),
    .X(_1517_));
 sky130_fd_sc_hd__nor2_4 _4613_ (.A(_0699_),
    .B(_0702_),
    .Y(_1518_));
 sky130_fd_sc_hd__buf_4 _4614_ (.A(_1518_),
    .X(_1519_));
 sky130_fd_sc_hd__o21a_1 _4615_ (.A1(\core_1.execute.rf.reg_outputs[4][15] ),
    .A2(_0701_),
    .B1(_0712_),
    .X(_1520_));
 sky130_fd_sc_hd__a31o_1 _4616_ (.A1(\core_1.execute.rf.reg_outputs[1][15] ),
    .A2(_0707_),
    .A3(_1519_),
    .B1(_1520_),
    .X(_1521_));
 sky130_fd_sc_hd__nor2_8 _4617_ (.A(_0706_),
    .B(_0704_),
    .Y(_1522_));
 sky130_fd_sc_hd__and3_4 _4618_ (.A(_0706_),
    .B(_0710_),
    .C(_0703_),
    .X(_1523_));
 sky130_fd_sc_hd__and3b_4 _4619_ (.A_N(\core_1.dec_l_reg_sel[0] ),
    .B(_0709_),
    .C(_0705_),
    .X(_1524_));
 sky130_fd_sc_hd__buf_4 _4620_ (.A(_1524_),
    .X(_1525_));
 sky130_fd_sc_hd__a22o_1 _4621_ (.A1(\core_1.execute.rf.reg_outputs[7][15] ),
    .A2(_1523_),
    .B1(_1525_),
    .B2(\core_1.execute.rf.reg_outputs[6][15] ),
    .X(_1526_));
 sky130_fd_sc_hd__a21o_1 _4622_ (.A1(\core_1.execute.rf.reg_outputs[3][15] ),
    .A2(_1522_),
    .B1(_1526_),
    .X(_1527_));
 sky130_fd_sc_hd__or3_2 _4623_ (.A(_1517_),
    .B(_1521_),
    .C(_1527_),
    .X(_1528_));
 sky130_fd_sc_hd__o21a_4 _4624_ (.A1(net94),
    .A2(_1513_),
    .B1(_1528_),
    .X(_1529_));
 sky130_fd_sc_hd__and2_1 _4625_ (.A(\core_1.execute.rf.reg_outputs[3][9] ),
    .B(_1522_),
    .X(_1530_));
 sky130_fd_sc_hd__a221o_1 _4626_ (.A1(\core_1.execute.rf.reg_outputs[5][9] ),
    .A2(_1514_),
    .B1(_1516_),
    .B2(\core_1.execute.rf.reg_outputs[2][9] ),
    .C1(_1530_),
    .X(_1531_));
 sky130_fd_sc_hd__or2_1 _4627_ (.A(\core_1.execute.rf.reg_outputs[4][9] ),
    .B(_0700_),
    .X(_1532_));
 sky130_fd_sc_hd__a32o_1 _4628_ (.A1(\core_1.execute.rf.reg_outputs[1][9] ),
    .A2(_0703_),
    .A3(_1519_),
    .B1(_1532_),
    .B2(_0712_),
    .X(_1533_));
 sky130_fd_sc_hd__a221o_1 _4629_ (.A1(\core_1.execute.rf.reg_outputs[7][9] ),
    .A2(_1523_),
    .B1(_1525_),
    .B2(\core_1.execute.rf.reg_outputs[6][9] ),
    .C1(_1533_),
    .X(_1534_));
 sky130_fd_sc_hd__o22a_4 _4630_ (.A1(net103),
    .A2(_1513_),
    .B1(_1531_),
    .B2(_1534_),
    .X(_1535_));
 sky130_fd_sc_hd__inv_2 _4631_ (.A(_1535_),
    .Y(_1536_));
 sky130_fd_sc_hd__a22o_1 _4632_ (.A1(\core_1.execute.rf.reg_outputs[3][10] ),
    .A2(_1522_),
    .B1(_1525_),
    .B2(\core_1.execute.rf.reg_outputs[6][10] ),
    .X(_1537_));
 sky130_fd_sc_hd__a21o_1 _4633_ (.A1(\core_1.execute.rf.reg_outputs[5][10] ),
    .A2(_1514_),
    .B1(_1537_),
    .X(_1538_));
 sky130_fd_sc_hd__o21a_1 _4634_ (.A1(\core_1.execute.rf.reg_outputs[4][10] ),
    .A2(_0701_),
    .B1(_0712_),
    .X(_1539_));
 sky130_fd_sc_hd__a32o_1 _4635_ (.A1(\core_1.execute.rf.reg_outputs[1][10] ),
    .A2(_0707_),
    .A3(_1519_),
    .B1(_1516_),
    .B2(\core_1.execute.rf.reg_outputs[2][10] ),
    .X(_1540_));
 sky130_fd_sc_hd__a211o_1 _4636_ (.A1(\core_1.execute.rf.reg_outputs[7][10] ),
    .A2(_1523_),
    .B1(_1539_),
    .C1(_1540_),
    .X(_1541_));
 sky130_fd_sc_hd__o22a_4 _4637_ (.A1(net89),
    .A2(_1513_),
    .B1(_1538_),
    .B2(_1541_),
    .X(_1542_));
 sky130_fd_sc_hd__buf_4 _4638_ (.A(_1542_),
    .X(_1543_));
 sky130_fd_sc_hd__nor2_1 _4639_ (.A(_1203_),
    .B(_1543_),
    .Y(_1544_));
 sky130_fd_sc_hd__a21o_1 _4640_ (.A1(_1203_),
    .A2(_1536_),
    .B1(_1544_),
    .X(_1545_));
 sky130_fd_sc_hd__clkinv_2 _4641_ (.A(_1545_),
    .Y(_1546_));
 sky130_fd_sc_hd__and2b_2 _4642_ (.A_N(\core_1.dec_l_reg_sel[1] ),
    .B(_0705_),
    .X(_1547_));
 sky130_fd_sc_hd__and2b_2 _4643_ (.A_N(_0705_),
    .B(\core_1.dec_l_reg_sel[1] ),
    .X(_1548_));
 sky130_fd_sc_hd__and3_1 _4644_ (.A(\core_1.execute.rf.reg_outputs[7][7] ),
    .B(_0706_),
    .C(_0710_),
    .X(_1549_));
 sky130_fd_sc_hd__a221o_1 _4645_ (.A1(\core_1.execute.rf.reg_outputs[5][7] ),
    .A2(_1547_),
    .B1(_1548_),
    .B2(\core_1.execute.rf.reg_outputs[3][7] ),
    .C1(_1549_),
    .X(_1550_));
 sky130_fd_sc_hd__a22o_1 _4646_ (.A1(\core_1.execute.rf.reg_outputs[6][7] ),
    .A2(_1525_),
    .B1(_1516_),
    .B2(\core_1.execute.rf.reg_outputs[2][7] ),
    .X(_1551_));
 sky130_fd_sc_hd__nor3b_4 _4647_ (.A(_0702_),
    .B(_0703_),
    .C_N(_0699_),
    .Y(_1552_));
 sky130_fd_sc_hd__nor3_4 _4648_ (.A(_0699_),
    .B(_0709_),
    .C(\core_1.dec_l_reg_sel[0] ),
    .Y(_1553_));
 sky130_fd_sc_hd__a221o_1 _4649_ (.A1(\core_1.execute.rf.reg_outputs[1][7] ),
    .A2(_1519_),
    .B1(_1552_),
    .B2(\core_1.execute.rf.reg_outputs[4][7] ),
    .C1(_1553_),
    .X(_1554_));
 sky130_fd_sc_hd__a211o_1 _4650_ (.A1(_0707_),
    .A2(_1550_),
    .B1(_1551_),
    .C1(_1554_),
    .X(_1555_));
 sky130_fd_sc_hd__o21a_4 _4651_ (.A1(net101),
    .A2(_1513_),
    .B1(_1555_),
    .X(_1556_));
 sky130_fd_sc_hd__buf_4 _4652_ (.A(_1556_),
    .X(_1557_));
 sky130_fd_sc_hd__and3_1 _4653_ (.A(\core_1.execute.rf.reg_outputs[1][8] ),
    .B(_0707_),
    .C(_1519_),
    .X(_1558_));
 sky130_fd_sc_hd__a221o_1 _4654_ (.A1(\core_1.execute.rf.reg_outputs[5][8] ),
    .A2(_1514_),
    .B1(_1516_),
    .B2(\core_1.execute.rf.reg_outputs[2][8] ),
    .C1(_1558_),
    .X(_1559_));
 sky130_fd_sc_hd__or2_1 _4655_ (.A(\core_1.execute.rf.reg_outputs[4][8] ),
    .B(_0700_),
    .X(_1560_));
 sky130_fd_sc_hd__a22o_1 _4656_ (.A1(\core_1.execute.rf.reg_outputs[6][8] ),
    .A2(_1525_),
    .B1(_1560_),
    .B2(_0712_),
    .X(_1561_));
 sky130_fd_sc_hd__a221o_1 _4657_ (.A1(\core_1.execute.rf.reg_outputs[7][8] ),
    .A2(_1523_),
    .B1(_1522_),
    .B2(\core_1.execute.rf.reg_outputs[3][8] ),
    .C1(_1561_),
    .X(_1562_));
 sky130_fd_sc_hd__o22a_4 _4658_ (.A1(net102),
    .A2(_1513_),
    .B1(_1559_),
    .B2(_1562_),
    .X(_1563_));
 sky130_fd_sc_hd__buf_4 _4659_ (.A(_1563_),
    .X(_1564_));
 sky130_fd_sc_hd__clkinv_2 _4660_ (.A(\core_1.execute.alu_mul_div.cbit[0] ),
    .Y(_1565_));
 sky130_fd_sc_hd__buf_4 _4661_ (.A(_1565_),
    .X(_1566_));
 sky130_fd_sc_hd__mux2_1 _4662_ (.A0(_1557_),
    .A1(_1564_),
    .S(_1566_),
    .X(_1567_));
 sky130_fd_sc_hd__mux2_1 _4663_ (.A0(_1546_),
    .A1(_1567_),
    .S(_1204_),
    .X(_1568_));
 sky130_fd_sc_hd__clkinv_2 _4664_ (.A(\core_1.execute.alu_mul_div.cbit[3] ),
    .Y(_1569_));
 sky130_fd_sc_hd__clkbuf_4 _4665_ (.A(\core_1.execute.alu_mul_div.cbit[2] ),
    .X(_1570_));
 sky130_fd_sc_hd__nand2_1 _4666_ (.A(_1569_),
    .B(_1570_),
    .Y(_1571_));
 sky130_fd_sc_hd__inv_2 _4667_ (.A(_1571_),
    .Y(_1572_));
 sky130_fd_sc_hd__a22o_1 _4668_ (.A1(\core_1.execute.rf.reg_outputs[5][12] ),
    .A2(_1514_),
    .B1(_1522_),
    .B2(\core_1.execute.rf.reg_outputs[3][12] ),
    .X(_1573_));
 sky130_fd_sc_hd__or2_1 _4669_ (.A(\core_1.execute.rf.reg_outputs[4][12] ),
    .B(_0701_),
    .X(_1574_));
 sky130_fd_sc_hd__buf_4 _4670_ (.A(_1519_),
    .X(_1575_));
 sky130_fd_sc_hd__and3_1 _4671_ (.A(\core_1.execute.rf.reg_outputs[1][12] ),
    .B(_0708_),
    .C(_1575_),
    .X(_1576_));
 sky130_fd_sc_hd__a221o_1 _4672_ (.A1(\core_1.execute.rf.reg_outputs[2][12] ),
    .A2(_1516_),
    .B1(_1574_),
    .B2(_0712_),
    .C1(_1576_),
    .X(_1577_));
 sky130_fd_sc_hd__a221o_1 _4673_ (.A1(\core_1.execute.rf.reg_outputs[7][12] ),
    .A2(_1523_),
    .B1(_1525_),
    .B2(\core_1.execute.rf.reg_outputs[6][12] ),
    .C1(_1577_),
    .X(_1578_));
 sky130_fd_sc_hd__o22a_4 _4674_ (.A1(net91),
    .A2(_1513_),
    .B1(_1573_),
    .B2(_1578_),
    .X(_1579_));
 sky130_fd_sc_hd__clkbuf_8 _4675_ (.A(_1579_),
    .X(_1580_));
 sky130_fd_sc_hd__a22o_1 _4676_ (.A1(\core_1.execute.rf.reg_outputs[7][11] ),
    .A2(_1523_),
    .B1(_1522_),
    .B2(\core_1.execute.rf.reg_outputs[3][11] ),
    .X(_1581_));
 sky130_fd_sc_hd__a21o_1 _4677_ (.A1(\core_1.execute.rf.reg_outputs[6][11] ),
    .A2(_1525_),
    .B1(_1581_),
    .X(_1582_));
 sky130_fd_sc_hd__a22o_1 _4678_ (.A1(\core_1.execute.rf.reg_outputs[5][11] ),
    .A2(_1514_),
    .B1(_1516_),
    .B2(\core_1.execute.rf.reg_outputs[2][11] ),
    .X(_1583_));
 sky130_fd_sc_hd__or2_1 _4679_ (.A(\core_1.execute.rf.reg_outputs[4][11] ),
    .B(_0701_),
    .X(_1584_));
 sky130_fd_sc_hd__a32o_1 _4680_ (.A1(\core_1.execute.rf.reg_outputs[1][11] ),
    .A2(_0707_),
    .A3(_1519_),
    .B1(_1584_),
    .B2(_0712_),
    .X(_1585_));
 sky130_fd_sc_hd__o32a_4 _4681_ (.A1(_1582_),
    .A2(_1583_),
    .A3(_1585_),
    .B1(_1513_),
    .B2(net90),
    .X(_1586_));
 sky130_fd_sc_hd__mux2_1 _4682_ (.A0(_1580_),
    .A1(_1586_),
    .S(_1203_),
    .X(_1587_));
 sky130_fd_sc_hd__a32o_1 _4683_ (.A1(\core_1.execute.rf.reg_outputs[1][14] ),
    .A2(_0708_),
    .A3(_1575_),
    .B1(_1525_),
    .B2(\core_1.execute.rf.reg_outputs[6][14] ),
    .X(_1588_));
 sky130_fd_sc_hd__a21o_1 _4684_ (.A1(\core_1.execute.rf.reg_outputs[7][14] ),
    .A2(_1523_),
    .B1(_1588_),
    .X(_1589_));
 sky130_fd_sc_hd__or2_1 _4685_ (.A(\core_1.execute.rf.reg_outputs[4][14] ),
    .B(_0701_),
    .X(_1590_));
 sky130_fd_sc_hd__a22o_1 _4686_ (.A1(\core_1.execute.rf.reg_outputs[3][14] ),
    .A2(_1522_),
    .B1(_1590_),
    .B2(_0712_),
    .X(_1591_));
 sky130_fd_sc_hd__a221o_1 _4687_ (.A1(\core_1.execute.rf.reg_outputs[5][14] ),
    .A2(_1514_),
    .B1(_1516_),
    .B2(\core_1.execute.rf.reg_outputs[2][14] ),
    .C1(_1591_),
    .X(_1592_));
 sky130_fd_sc_hd__o22a_4 _4688_ (.A1(net93),
    .A2(_1513_),
    .B1(_1589_),
    .B2(_1592_),
    .X(_1593_));
 sky130_fd_sc_hd__buf_4 _4689_ (.A(_1593_),
    .X(_1594_));
 sky130_fd_sc_hd__nor2_2 _4690_ (.A(_1203_),
    .B(_1204_),
    .Y(_1595_));
 sky130_fd_sc_hd__a22o_1 _4691_ (.A1(\core_1.execute.rf.reg_outputs[5][13] ),
    .A2(_1514_),
    .B1(_1525_),
    .B2(\core_1.execute.rf.reg_outputs[6][13] ),
    .X(_1596_));
 sky130_fd_sc_hd__o21a_1 _4692_ (.A1(\core_1.execute.rf.reg_outputs[4][13] ),
    .A2(_0701_),
    .B1(_0712_),
    .X(_1597_));
 sky130_fd_sc_hd__a32o_1 _4693_ (.A1(\core_1.execute.rf.reg_outputs[1][13] ),
    .A2(_0707_),
    .A3(_1519_),
    .B1(_1522_),
    .B2(\core_1.execute.rf.reg_outputs[3][13] ),
    .X(_1598_));
 sky130_fd_sc_hd__a211o_1 _4694_ (.A1(\core_1.execute.rf.reg_outputs[2][13] ),
    .A2(_1516_),
    .B1(_1597_),
    .C1(_1598_),
    .X(_1599_));
 sky130_fd_sc_hd__a211o_1 _4695_ (.A1(\core_1.execute.rf.reg_outputs[7][13] ),
    .A2(_1523_),
    .B1(_1596_),
    .C1(_1599_),
    .X(_1600_));
 sky130_fd_sc_hd__o21ai_4 _4696_ (.A1(net92),
    .A2(_1513_),
    .B1(_1600_),
    .Y(_1601_));
 sky130_fd_sc_hd__inv_2 _4697_ (.A(\core_1.execute.alu_mul_div.cbit[1] ),
    .Y(_1602_));
 sky130_fd_sc_hd__clkbuf_4 _4698_ (.A(_1602_),
    .X(_1603_));
 sky130_fd_sc_hd__nand2_2 _4699_ (.A(_1203_),
    .B(_1603_),
    .Y(_1604_));
 sky130_fd_sc_hd__nor2_1 _4700_ (.A(_1601_),
    .B(_1604_),
    .Y(_1605_));
 sky130_fd_sc_hd__a221o_1 _4701_ (.A1(_1204_),
    .A2(_1587_),
    .B1(_1594_),
    .B2(_1595_),
    .C1(_1605_),
    .X(_1606_));
 sky130_fd_sc_hd__nor2_2 _4702_ (.A(_1199_),
    .B(_1570_),
    .Y(_1607_));
 sky130_fd_sc_hd__buf_4 _4703_ (.A(_1569_),
    .X(_1608_));
 sky130_fd_sc_hd__and3b_1 _4704_ (.A_N(_0702_),
    .B(_0699_),
    .C(\core_1.execute.rf.reg_outputs[5][2] ),
    .X(_1609_));
 sky130_fd_sc_hd__and3b_1 _4705_ (.A_N(_0706_),
    .B(_0702_),
    .C(\core_1.execute.rf.reg_outputs[3][2] ),
    .X(_1610_));
 sky130_fd_sc_hd__and3_1 _4706_ (.A(\core_1.execute.rf.reg_outputs[7][2] ),
    .B(_0706_),
    .C(_0702_),
    .X(_1611_));
 sky130_fd_sc_hd__o31a_1 _4707_ (.A1(_1609_),
    .A2(_1610_),
    .A3(_1611_),
    .B1(_0703_),
    .X(_1612_));
 sky130_fd_sc_hd__a221o_1 _4708_ (.A1(\core_1.execute.rf.reg_outputs[1][2] ),
    .A2(_1518_),
    .B1(_1515_),
    .B2(\core_1.execute.rf.reg_outputs[2][2] ),
    .C1(_1553_),
    .X(_1613_));
 sky130_fd_sc_hd__a22o_1 _4709_ (.A1(\core_1.execute.rf.reg_outputs[6][2] ),
    .A2(_1524_),
    .B1(_1552_),
    .B2(\core_1.execute.rf.reg_outputs[4][2] ),
    .X(_1614_));
 sky130_fd_sc_hd__or3_4 _4710_ (.A(_1612_),
    .B(_1613_),
    .C(_1614_),
    .X(_1615_));
 sky130_fd_sc_hd__or2_2 _4711_ (.A(net96),
    .B(_1512_),
    .X(_1616_));
 sky130_fd_sc_hd__a21oi_1 _4712_ (.A1(_1615_),
    .A2(_1616_),
    .B1(\core_1.execute.alu_mul_div.cbit[0] ),
    .Y(_1617_));
 sky130_fd_sc_hd__or2_2 _4713_ (.A(net95),
    .B(_1512_),
    .X(_1618_));
 sky130_fd_sc_hd__a22o_1 _4714_ (.A1(\core_1.execute.rf.reg_outputs[6][1] ),
    .A2(_1524_),
    .B1(_1552_),
    .B2(\core_1.execute.rf.reg_outputs[4][1] ),
    .X(_1619_));
 sky130_fd_sc_hd__and3_1 _4715_ (.A(\core_1.execute.rf.reg_outputs[7][1] ),
    .B(_0699_),
    .C(_0709_),
    .X(_1620_));
 sky130_fd_sc_hd__and3b_1 _4716_ (.A_N(_0702_),
    .B(_0699_),
    .C(\core_1.execute.rf.reg_outputs[5][1] ),
    .X(_1621_));
 sky130_fd_sc_hd__and3b_1 _4717_ (.A_N(_0699_),
    .B(_0709_),
    .C(\core_1.execute.rf.reg_outputs[3][1] ),
    .X(_1622_));
 sky130_fd_sc_hd__o31a_1 _4718_ (.A1(_1620_),
    .A2(_1621_),
    .A3(_1622_),
    .B1(_0703_),
    .X(_1623_));
 sky130_fd_sc_hd__a221o_1 _4719_ (.A1(\core_1.execute.rf.reg_outputs[1][1] ),
    .A2(_1518_),
    .B1(_1515_),
    .B2(\core_1.execute.rf.reg_outputs[2][1] ),
    .C1(_1553_),
    .X(_1624_));
 sky130_fd_sc_hd__or3_4 _4720_ (.A(_1619_),
    .B(_1623_),
    .C(_1624_),
    .X(_1625_));
 sky130_fd_sc_hd__a21oi_1 _4721_ (.A1(_1618_),
    .A2(_1625_),
    .B1(_1565_),
    .Y(_1626_));
 sky130_fd_sc_hd__and3_1 _4722_ (.A(\core_1.execute.rf.reg_outputs[7][0] ),
    .B(_0705_),
    .C(\core_1.dec_l_reg_sel[1] ),
    .X(_1627_));
 sky130_fd_sc_hd__and3b_1 _4723_ (.A_N(_0709_),
    .B(_0705_),
    .C(\core_1.execute.rf.reg_outputs[5][0] ),
    .X(_1628_));
 sky130_fd_sc_hd__and3b_1 _4724_ (.A_N(_0705_),
    .B(_0709_),
    .C(\core_1.execute.rf.reg_outputs[3][0] ),
    .X(_1629_));
 sky130_fd_sc_hd__o31a_2 _4725_ (.A1(_1627_),
    .A2(_1628_),
    .A3(_1629_),
    .B1(_0703_),
    .X(_1630_));
 sky130_fd_sc_hd__or2b_1 _4726_ (.A(\core_1.execute.rf.reg_outputs[4][0] ),
    .B_N(_0699_),
    .X(_1631_));
 sky130_fd_sc_hd__a22o_2 _4727_ (.A1(\core_1.execute.rf.reg_outputs[1][0] ),
    .A2(_1518_),
    .B1(_1631_),
    .B2(_0712_),
    .X(_1632_));
 sky130_fd_sc_hd__a22o_2 _4728_ (.A1(\core_1.execute.rf.reg_outputs[6][0] ),
    .A2(_1524_),
    .B1(_1515_),
    .B2(\core_1.execute.rf.reg_outputs[2][0] ),
    .X(_1633_));
 sky130_fd_sc_hd__or2_2 _4729_ (.A(net88),
    .B(_1512_),
    .X(_1634_));
 sky130_fd_sc_hd__o31ai_4 _4730_ (.A1(_1630_),
    .A2(_1632_),
    .A3(_1633_),
    .B1(_1634_),
    .Y(_1635_));
 sky130_fd_sc_hd__nand2_2 _4731_ (.A(_1566_),
    .B(\core_1.execute.alu_mul_div.cbit[1] ),
    .Y(_1636_));
 sky130_fd_sc_hd__o32a_2 _4732_ (.A1(\core_1.execute.alu_mul_div.cbit[1] ),
    .A2(_1617_),
    .A3(_1626_),
    .B1(_1635_),
    .B2(_1636_),
    .X(_1637_));
 sky130_fd_sc_hd__and3_1 _4733_ (.A(\core_1.execute.rf.reg_outputs[7][3] ),
    .B(_0706_),
    .C(_0710_),
    .X(_1638_));
 sky130_fd_sc_hd__a221o_4 _4734_ (.A1(\core_1.execute.rf.reg_outputs[5][3] ),
    .A2(_1547_),
    .B1(_1548_),
    .B2(\core_1.execute.rf.reg_outputs[3][3] ),
    .C1(_1638_),
    .X(_1639_));
 sky130_fd_sc_hd__a22o_1 _4735_ (.A1(\core_1.execute.rf.reg_outputs[1][3] ),
    .A2(_1519_),
    .B1(_1515_),
    .B2(\core_1.execute.rf.reg_outputs[2][3] ),
    .X(_1640_));
 sky130_fd_sc_hd__a22o_1 _4736_ (.A1(\core_1.execute.rf.reg_outputs[6][3] ),
    .A2(_1524_),
    .B1(_1552_),
    .B2(\core_1.execute.rf.reg_outputs[4][3] ),
    .X(_1641_));
 sky130_fd_sc_hd__o21a_2 _4737_ (.A1(_1640_),
    .A2(_1641_),
    .B1(_1512_),
    .X(_1642_));
 sky130_fd_sc_hd__a221oi_4 _4738_ (.A1(net97),
    .A2(_1553_),
    .B1(_1639_),
    .B2(_0707_),
    .C1(_1642_),
    .Y(_1643_));
 sky130_fd_sc_hd__a22o_1 _4739_ (.A1(\core_1.execute.rf.reg_outputs[6][4] ),
    .A2(_1524_),
    .B1(_1515_),
    .B2(\core_1.execute.rf.reg_outputs[2][4] ),
    .X(_1644_));
 sky130_fd_sc_hd__a22o_1 _4740_ (.A1(\core_1.execute.rf.reg_outputs[1][4] ),
    .A2(_1518_),
    .B1(_1552_),
    .B2(\core_1.execute.rf.reg_outputs[4][4] ),
    .X(_1645_));
 sky130_fd_sc_hd__o21a_2 _4741_ (.A1(_1644_),
    .A2(_1645_),
    .B1(_1512_),
    .X(_1646_));
 sky130_fd_sc_hd__and3_1 _4742_ (.A(\core_1.execute.rf.reg_outputs[7][4] ),
    .B(_0699_),
    .C(_0702_),
    .X(_1647_));
 sky130_fd_sc_hd__a221o_1 _4743_ (.A1(\core_1.execute.rf.reg_outputs[5][4] ),
    .A2(_1547_),
    .B1(_1548_),
    .B2(\core_1.execute.rf.reg_outputs[3][4] ),
    .C1(_1647_),
    .X(_1648_));
 sky130_fd_sc_hd__and2_1 _4744_ (.A(_0707_),
    .B(_1648_),
    .X(_1649_));
 sky130_fd_sc_hd__a211oi_4 _4745_ (.A1(net98),
    .A2(_1553_),
    .B1(_1646_),
    .C1(_1649_),
    .Y(_1650_));
 sky130_fd_sc_hd__mux2_1 _4746_ (.A0(_1643_),
    .A1(_1650_),
    .S(_1566_),
    .X(_1651_));
 sky130_fd_sc_hd__a22o_1 _4747_ (.A1(\core_1.execute.rf.reg_outputs[1][6] ),
    .A2(_1519_),
    .B1(_1525_),
    .B2(\core_1.execute.rf.reg_outputs[6][6] ),
    .X(_1652_));
 sky130_fd_sc_hd__a221o_2 _4748_ (.A1(\core_1.execute.rf.reg_outputs[2][6] ),
    .A2(_1516_),
    .B1(_1552_),
    .B2(\core_1.execute.rf.reg_outputs[4][6] ),
    .C1(_1652_),
    .X(_1653_));
 sky130_fd_sc_hd__and3_1 _4749_ (.A(\core_1.execute.rf.reg_outputs[7][6] ),
    .B(_0706_),
    .C(_0702_),
    .X(_1654_));
 sky130_fd_sc_hd__a221o_1 _4750_ (.A1(\core_1.execute.rf.reg_outputs[5][6] ),
    .A2(_1547_),
    .B1(_1548_),
    .B2(\core_1.execute.rf.reg_outputs[3][6] ),
    .C1(_1654_),
    .X(_1655_));
 sky130_fd_sc_hd__a22o_1 _4751_ (.A1(net100),
    .A2(_1553_),
    .B1(_1655_),
    .B2(_0707_),
    .X(_1656_));
 sky130_fd_sc_hd__a21o_2 _4752_ (.A1(_1512_),
    .A2(_1653_),
    .B1(_1656_),
    .X(_1657_));
 sky130_fd_sc_hd__buf_4 _4753_ (.A(_1657_),
    .X(_1658_));
 sky130_fd_sc_hd__and3_1 _4754_ (.A(\core_1.execute.rf.reg_outputs[7][5] ),
    .B(_0705_),
    .C(\core_1.dec_l_reg_sel[1] ),
    .X(_1659_));
 sky130_fd_sc_hd__a221o_1 _4755_ (.A1(\core_1.execute.rf.reg_outputs[5][5] ),
    .A2(_1547_),
    .B1(_1548_),
    .B2(\core_1.execute.rf.reg_outputs[3][5] ),
    .C1(_1659_),
    .X(_1660_));
 sky130_fd_sc_hd__and2_1 _4756_ (.A(_0703_),
    .B(_1660_),
    .X(_1661_));
 sky130_fd_sc_hd__a221o_1 _4757_ (.A1(\core_1.execute.rf.reg_outputs[1][5] ),
    .A2(_1518_),
    .B1(_1552_),
    .B2(\core_1.execute.rf.reg_outputs[4][5] ),
    .C1(_1553_),
    .X(_1662_));
 sky130_fd_sc_hd__a22o_1 _4758_ (.A1(\core_1.execute.rf.reg_outputs[6][5] ),
    .A2(_1524_),
    .B1(_1515_),
    .B2(\core_1.execute.rf.reg_outputs[2][5] ),
    .X(_1663_));
 sky130_fd_sc_hd__o32a_4 _4759_ (.A1(_1661_),
    .A2(_1662_),
    .A3(_1663_),
    .B1(_1512_),
    .B2(net99),
    .X(_1664_));
 sky130_fd_sc_hd__buf_4 _4760_ (.A(_1664_),
    .X(_1665_));
 sky130_fd_sc_hd__mux2_1 _4761_ (.A0(_1658_),
    .A1(_1665_),
    .S(_1203_),
    .X(_1666_));
 sky130_fd_sc_hd__nor2_1 _4762_ (.A(\core_1.execute.alu_mul_div.cbit[1] ),
    .B(_1666_),
    .Y(_1667_));
 sky130_fd_sc_hd__a21o_1 _4763_ (.A1(\core_1.execute.alu_mul_div.cbit[1] ),
    .A2(_1651_),
    .B1(_1667_),
    .X(_1668_));
 sky130_fd_sc_hd__mux2_1 _4764_ (.A0(_1637_),
    .A1(_1668_),
    .S(_1202_),
    .X(_1669_));
 sky130_fd_sc_hd__nor2_1 _4765_ (.A(_1608_),
    .B(_1669_),
    .Y(_1670_));
 sky130_fd_sc_hd__a221o_2 _4766_ (.A1(_1568_),
    .A2(_1572_),
    .B1(_1606_),
    .B2(_1607_),
    .C1(_1670_),
    .X(_1671_));
 sky130_fd_sc_hd__a211o_1 _4767_ (.A1(_1416_),
    .A2(_1421_),
    .B1(_1671_),
    .C1(_1413_),
    .X(_1672_));
 sky130_fd_sc_hd__o211a_1 _4768_ (.A1(\core_1.execute.alu_mul_div.div_cur[0] ),
    .A2(_1409_),
    .B1(_1672_),
    .C1(_1428_),
    .X(_1673_));
 sky130_fd_sc_hd__a21o_1 _4769_ (.A1(_1511_),
    .A2(_1529_),
    .B1(_1673_),
    .X(_0186_));
 sky130_fd_sc_hd__a21o_1 _4770_ (.A1(\core_1.dec_jump_cond_code[4] ),
    .A2(_1047_),
    .B1(\core_1.dec_pc_inc ),
    .X(_1674_));
 sky130_fd_sc_hd__a31o_1 _4771_ (.A1(net211),
    .A2(_1029_),
    .A3(_1674_),
    .B1(net79),
    .X(_1675_));
 sky130_fd_sc_hd__inv_2 _4772_ (.A(_1047_),
    .Y(_1676_));
 sky130_fd_sc_hd__a21o_1 _4773_ (.A1(\core_1.dec_jump_cond_code[4] ),
    .A2(_1676_),
    .B1(_1058_),
    .X(_1677_));
 sky130_fd_sc_hd__nand2_1 _4774_ (.A(_0737_),
    .B(_1677_),
    .Y(_1678_));
 sky130_fd_sc_hd__clkbuf_4 _4775_ (.A(_1678_),
    .X(_1679_));
 sky130_fd_sc_hd__and2_1 _4776_ (.A(_0737_),
    .B(_1674_),
    .X(_1680_));
 sky130_fd_sc_hd__buf_4 _4777_ (.A(_1680_),
    .X(_1681_));
 sky130_fd_sc_hd__nand3_1 _4778_ (.A(net211),
    .B(net79),
    .C(_1681_),
    .Y(_1682_));
 sky130_fd_sc_hd__a31o_1 _4779_ (.A1(_1675_),
    .A2(_1679_),
    .A3(_1682_),
    .B1(_0670_),
    .X(_1683_));
 sky130_fd_sc_hd__nor2_1 _4780_ (.A(_1057_),
    .B(_1153_),
    .Y(_1684_));
 sky130_fd_sc_hd__inv_2 _4781_ (.A(\core_1.execute.alu_mul_div.i_mod ),
    .Y(_1685_));
 sky130_fd_sc_hd__clkbuf_4 _4782_ (.A(_1685_),
    .X(_1686_));
 sky130_fd_sc_hd__a21bo_1 _4783_ (.A1(\core_1.execute.alu_mul_div.div_res[1] ),
    .A2(_1686_),
    .B1_N(_1407_),
    .X(_1687_));
 sky130_fd_sc_hd__buf_2 _4784_ (.A(_0958_),
    .X(_1688_));
 sky130_fd_sc_hd__o21a_4 _4785_ (.A1(_1077_),
    .A2(_0639_),
    .B1(_1367_),
    .X(_1689_));
 sky130_fd_sc_hd__and2_1 _4786_ (.A(_1374_),
    .B(_1375_),
    .X(_1690_));
 sky130_fd_sc_hd__buf_4 _4787_ (.A(_1690_),
    .X(_1691_));
 sky130_fd_sc_hd__nand2_4 _4788_ (.A(_1377_),
    .B(_1378_),
    .Y(_1692_));
 sky130_fd_sc_hd__buf_4 _4789_ (.A(_1692_),
    .X(_1693_));
 sky130_fd_sc_hd__nor2_2 _4790_ (.A(_1691_),
    .B(_1693_),
    .Y(_1694_));
 sky130_fd_sc_hd__o21ai_4 _4791_ (.A1(net94),
    .A2(_1513_),
    .B1(_1528_),
    .Y(_1695_));
 sky130_fd_sc_hd__o21ai_4 _4792_ (.A1(_1077_),
    .A2(_0627_),
    .B1(_1356_),
    .Y(_1696_));
 sky130_fd_sc_hd__o21ai_2 _4793_ (.A1(_1077_),
    .A2(_0614_),
    .B1(_1348_),
    .Y(_1697_));
 sky130_fd_sc_hd__or4_2 _4794_ (.A(_1343_),
    .B(_1347_),
    .C(_1697_),
    .D(_1351_),
    .X(_1698_));
 sky130_fd_sc_hd__mux2_4 _4795_ (.A0(net182),
    .A1(net198),
    .S(_1320_),
    .X(_1699_));
 sky130_fd_sc_hd__a2111o_1 _4796_ (.A1(_1076_),
    .A2(net184),
    .B1(_1316_),
    .C1(_1319_),
    .D1(_1321_),
    .X(_1700_));
 sky130_fd_sc_hd__a2111o_1 _4797_ (.A1(_1076_),
    .A2(net180),
    .B1(_1334_),
    .C1(_1337_),
    .D1(_1338_),
    .X(_1701_));
 sky130_fd_sc_hd__or4_4 _4798_ (.A(_1699_),
    .B(_1329_),
    .C(_1700_),
    .D(_1701_),
    .X(_1702_));
 sky130_fd_sc_hd__or3_4 _4799_ (.A(_1696_),
    .B(_1698_),
    .C(_1702_),
    .X(_1703_));
 sky130_fd_sc_hd__nor2_1 _4800_ (.A(_1695_),
    .B(_1703_),
    .Y(_1704_));
 sky130_fd_sc_hd__nand2_2 _4801_ (.A(_1374_),
    .B(_1375_),
    .Y(_1705_));
 sky130_fd_sc_hd__buf_4 _4802_ (.A(_1705_),
    .X(_1706_));
 sky130_fd_sc_hd__nor2_1 _4803_ (.A(_1418_),
    .B(_1703_),
    .Y(_1707_));
 sky130_fd_sc_hd__nor3_2 _4804_ (.A(_1696_),
    .B(_1698_),
    .C(_1702_),
    .Y(_1708_));
 sky130_fd_sc_hd__nand2_2 _4805_ (.A(_1418_),
    .B(_1708_),
    .Y(_1709_));
 sky130_fd_sc_hd__o2bb2a_1 _4806_ (.A1_N(_1594_),
    .A2_N(_1707_),
    .B1(_1709_),
    .B2(_1601_),
    .X(_1710_));
 sky130_fd_sc_hd__o2bb2a_1 _4807_ (.A1_N(_1694_),
    .A2_N(_1704_),
    .B1(_1706_),
    .B2(_1710_),
    .X(_1711_));
 sky130_fd_sc_hd__buf_2 _4808_ (.A(_1707_),
    .X(_1712_));
 sky130_fd_sc_hd__nor2_2 _4809_ (.A(_1692_),
    .B(_1703_),
    .Y(_1713_));
 sky130_fd_sc_hd__a22oi_1 _4810_ (.A1(_1580_),
    .A2(_1712_),
    .B1(_1713_),
    .B2(_1586_),
    .Y(_1714_));
 sky130_fd_sc_hd__o2bb2a_1 _4811_ (.A1_N(_1543_),
    .A2_N(_1712_),
    .B1(_1709_),
    .B2(_1536_),
    .X(_1715_));
 sky130_fd_sc_hd__mux2_1 _4812_ (.A0(_1714_),
    .A1(_1715_),
    .S(_1691_),
    .X(_1716_));
 sky130_fd_sc_hd__mux2_1 _4813_ (.A0(_1711_),
    .A1(_1716_),
    .S(_1384_),
    .X(_1717_));
 sky130_fd_sc_hd__a22o_1 _4814_ (.A1(_1658_),
    .A2(_1712_),
    .B1(_1713_),
    .B2(_1665_),
    .X(_1718_));
 sky130_fd_sc_hd__clkinv_2 _4815_ (.A(_1718_),
    .Y(_1719_));
 sky130_fd_sc_hd__a22oi_1 _4816_ (.A1(_1564_),
    .A2(_1712_),
    .B1(_1713_),
    .B2(_1557_),
    .Y(_1720_));
 sky130_fd_sc_hd__mux2_1 _4817_ (.A0(_1719_),
    .A1(_1720_),
    .S(_1706_),
    .X(_1721_));
 sky130_fd_sc_hd__nor2_1 _4818_ (.A(_1689_),
    .B(_1384_),
    .Y(_1722_));
 sky130_fd_sc_hd__a221o_4 _4819_ (.A1(net97),
    .A2(_1553_),
    .B1(_1639_),
    .B2(_0708_),
    .C1(_1642_),
    .X(_1723_));
 sky130_fd_sc_hd__a211o_4 _4820_ (.A1(net98),
    .A2(_1553_),
    .B1(_1646_),
    .C1(_1649_),
    .X(_1724_));
 sky130_fd_sc_hd__mux2_1 _4821_ (.A0(_1723_),
    .A1(_1724_),
    .S(_1693_),
    .X(_1725_));
 sky130_fd_sc_hd__nor2_1 _4822_ (.A(_1691_),
    .B(_1725_),
    .Y(_1726_));
 sky130_fd_sc_hd__nand2_8 _4823_ (.A(_1615_),
    .B(_1616_),
    .Y(_1727_));
 sky130_fd_sc_hd__nor2_2 _4824_ (.A(_1705_),
    .B(_1417_),
    .Y(_1728_));
 sky130_fd_sc_hd__and4_1 _4825_ (.A(_1374_),
    .B(_1375_),
    .C(_1377_),
    .D(_1378_),
    .X(_1729_));
 sky130_fd_sc_hd__clkbuf_4 _4826_ (.A(_1729_),
    .X(_1730_));
 sky130_fd_sc_hd__nand2_4 _4827_ (.A(_1618_),
    .B(_1625_),
    .Y(_1731_));
 sky130_fd_sc_hd__a22o_1 _4828_ (.A1(_1727_),
    .A2(_1728_),
    .B1(_1730_),
    .B2(_1731_),
    .X(_1732_));
 sky130_fd_sc_hd__or3_1 _4829_ (.A(_1703_),
    .B(_1726_),
    .C(_1732_),
    .X(_1733_));
 sky130_fd_sc_hd__nor2_2 _4830_ (.A(_1689_),
    .B(_1372_),
    .Y(_1734_));
 sky130_fd_sc_hd__nor2_1 _4831_ (.A(\core_1.decode.oc_alu_mode[1] ),
    .B(_0988_),
    .Y(_1735_));
 sky130_fd_sc_hd__or2_2 _4832_ (.A(_1361_),
    .B(_1735_),
    .X(_1736_));
 sky130_fd_sc_hd__a221o_1 _4833_ (.A1(_1721_),
    .A2(_1722_),
    .B1(_1733_),
    .B2(_1734_),
    .C1(_1736_),
    .X(_1737_));
 sky130_fd_sc_hd__a21oi_1 _4834_ (.A1(_1689_),
    .A2(_1717_),
    .B1(_1737_),
    .Y(_1738_));
 sky130_fd_sc_hd__a21oi_2 _4835_ (.A1(\core_1.decode.oc_alu_mode[12] ),
    .A2(_1692_),
    .B1(_1690_),
    .Y(_1739_));
 sky130_fd_sc_hd__a21o_2 _4836_ (.A1(_0988_),
    .A2(_1728_),
    .B1(_1739_),
    .X(_1740_));
 sky130_fd_sc_hd__o31a_4 _4837_ (.A1(_1630_),
    .A2(_1632_),
    .A3(_1633_),
    .B1(_1634_),
    .X(_1741_));
 sky130_fd_sc_hd__inv_2 _4838_ (.A(\core_1.decode.oc_alu_mode[12] ),
    .Y(_1742_));
 sky130_fd_sc_hd__a311oi_2 _4839_ (.A1(_1368_),
    .A2(_1383_),
    .A3(_1730_),
    .B1(_1364_),
    .C1(_1742_),
    .Y(_1743_));
 sky130_fd_sc_hd__nor2_1 _4840_ (.A(_1742_),
    .B(_1357_),
    .Y(_1744_));
 sky130_fd_sc_hd__or4_4 _4841_ (.A(_1698_),
    .B(_1702_),
    .C(_1743_),
    .D(_1744_),
    .X(_1745_));
 sky130_fd_sc_hd__nor2_1 _4842_ (.A(_1742_),
    .B(_1529_),
    .Y(_1746_));
 sky130_fd_sc_hd__nor2_4 _4843_ (.A(_1745_),
    .B(_1746_),
    .Y(_1747_));
 sky130_fd_sc_hd__buf_2 _4844_ (.A(_1747_),
    .X(_1748_));
 sky130_fd_sc_hd__o21ai_1 _4845_ (.A1(_0988_),
    .A2(_1741_),
    .B1(_1748_),
    .Y(_1749_));
 sky130_fd_sc_hd__buf_2 _4846_ (.A(\core_1.decode.oc_alu_mode[12] ),
    .X(_1750_));
 sky130_fd_sc_hd__and2_4 _4847_ (.A(_1618_),
    .B(_1625_),
    .X(_1751_));
 sky130_fd_sc_hd__o21ai_1 _4848_ (.A1(_1750_),
    .A2(_1751_),
    .B1(_1747_),
    .Y(_1752_));
 sky130_fd_sc_hd__mux2_1 _4849_ (.A0(_1749_),
    .A1(_1752_),
    .S(_1419_),
    .X(_1753_));
 sky130_fd_sc_hd__nor2_1 _4850_ (.A(_1740_),
    .B(_1753_),
    .Y(_1754_));
 sky130_fd_sc_hd__and3_1 _4851_ (.A(_0988_),
    .B(_1730_),
    .C(_1734_),
    .X(_1755_));
 sky130_fd_sc_hd__xnor2_2 _4852_ (.A(_1361_),
    .B(_1755_),
    .Y(_1756_));
 sky130_fd_sc_hd__o211ai_4 _4853_ (.A1(_0988_),
    .A2(\core_1.decode.oc_alu_mode[13] ),
    .B1(_1357_),
    .C1(_1756_),
    .Y(_1757_));
 sky130_fd_sc_hd__nand2_1 _4854_ (.A(_1384_),
    .B(_1730_),
    .Y(_1758_));
 sky130_fd_sc_hd__nand2_1 _4855_ (.A(_1750_),
    .B(_1758_),
    .Y(_1759_));
 sky130_fd_sc_hd__xnor2_1 _4856_ (.A(_1369_),
    .B(_1759_),
    .Y(_1760_));
 sky130_fd_sc_hd__clkinv_2 _4857_ (.A(_1760_),
    .Y(_1761_));
 sky130_fd_sc_hd__nor2_4 _4858_ (.A(_1757_),
    .B(_1761_),
    .Y(_1762_));
 sky130_fd_sc_hd__nor2_4 _4859_ (.A(_1742_),
    .B(_1730_),
    .Y(_1763_));
 sky130_fd_sc_hd__xnor2_4 _4860_ (.A(_1372_),
    .B(_1763_),
    .Y(_1764_));
 sky130_fd_sc_hd__buf_2 _4861_ (.A(_1764_),
    .X(_1765_));
 sky130_fd_sc_hd__nand2_2 _4862_ (.A(\core_1.execute.alu_flag_reg.o_d[1] ),
    .B(\core_1.dec_alu_carry_en ),
    .Y(_1766_));
 sky130_fd_sc_hd__and2_1 _4863_ (.A(_1741_),
    .B(_1766_),
    .X(_1767_));
 sky130_fd_sc_hd__or2_1 _4864_ (.A(_1741_),
    .B(_1766_),
    .X(_1768_));
 sky130_fd_sc_hd__o211a_1 _4865_ (.A1(_1417_),
    .A2(_1767_),
    .B1(_1768_),
    .C1(_1751_),
    .X(_1769_));
 sky130_fd_sc_hd__a311o_1 _4866_ (.A1(_1377_),
    .A2(_1378_),
    .A3(_1768_),
    .B1(_1767_),
    .C1(_1751_),
    .X(_1770_));
 sky130_fd_sc_hd__or2b_1 _4867_ (.A(_1769_),
    .B_N(_1770_),
    .X(_1771_));
 sky130_fd_sc_hd__nand2_1 _4868_ (.A(_1706_),
    .B(_1771_),
    .Y(_1772_));
 sky130_fd_sc_hd__or2_1 _4869_ (.A(_1706_),
    .B(_1771_),
    .X(_1773_));
 sky130_fd_sc_hd__nor2_1 _4870_ (.A(_1705_),
    .B(_1751_),
    .Y(_1774_));
 sky130_fd_sc_hd__nor2_1 _4871_ (.A(_1690_),
    .B(_1731_),
    .Y(_1775_));
 sky130_fd_sc_hd__nor2_1 _4872_ (.A(_1774_),
    .B(_1775_),
    .Y(_1776_));
 sky130_fd_sc_hd__and3_1 _4873_ (.A(_1377_),
    .B(_1378_),
    .C(_1635_),
    .X(_1777_));
 sky130_fd_sc_hd__a21oi_1 _4874_ (.A1(_1377_),
    .A2(_1378_),
    .B1(_1635_),
    .Y(_1778_));
 sky130_fd_sc_hd__o21bai_2 _4875_ (.A1(_1766_),
    .A2(_1777_),
    .B1_N(_1778_),
    .Y(_1779_));
 sky130_fd_sc_hd__o21ai_1 _4876_ (.A1(_1776_),
    .A2(_1779_),
    .B1(\core_1.decode.oc_alu_mode[4] ),
    .Y(_1780_));
 sky130_fd_sc_hd__a21oi_1 _4877_ (.A1(_1776_),
    .A2(_1779_),
    .B1(_1780_),
    .Y(_1781_));
 sky130_fd_sc_hd__nand2_1 _4878_ (.A(_1690_),
    .B(_1731_),
    .Y(_1782_));
 sky130_fd_sc_hd__or4_1 _4879_ (.A(\core_1.decode.oc_alu_mode[9] ),
    .B(\core_1.decode.oc_alu_mode[13] ),
    .C(\core_1.decode.oc_alu_mode[3] ),
    .D(\core_1.decode.oc_alu_mode[2] ),
    .X(_1783_));
 sky130_fd_sc_hd__or4_1 _4880_ (.A(\core_1.decode.oc_alu_mode[1] ),
    .B(\core_1.decode.oc_alu_mode[6] ),
    .C(\core_1.decode.oc_alu_mode[7] ),
    .D(\core_1.decode.oc_alu_mode[12] ),
    .X(_1784_));
 sky130_fd_sc_hd__inv_4 _4881_ (.A(\core_1.decode.oc_alu_mode[4] ),
    .Y(_1785_));
 sky130_fd_sc_hd__inv_2 _4882_ (.A(\core_1.decode.oc_alu_mode[11] ),
    .Y(_1786_));
 sky130_fd_sc_hd__and4bb_4 _4883_ (.A_N(_1783_),
    .B_N(_1784_),
    .C(_1785_),
    .D(_1786_),
    .X(_1787_));
 sky130_fd_sc_hd__nor2_2 _4884_ (.A(\core_1.decode.oc_alu_mode[3] ),
    .B(_1787_),
    .Y(_1788_));
 sky130_fd_sc_hd__nor2_1 _4885_ (.A(_1731_),
    .B(_1788_),
    .Y(_1789_));
 sky130_fd_sc_hd__a221o_1 _4886_ (.A1(\core_1.decode.oc_alu_mode[7] ),
    .A2(_1705_),
    .B1(_1782_),
    .B2(\core_1.decode.oc_alu_mode[9] ),
    .C1(_1789_),
    .X(_1790_));
 sky130_fd_sc_hd__a221o_1 _4887_ (.A1(\core_1.decode.oc_alu_mode[2] ),
    .A2(_1775_),
    .B1(_1776_),
    .B2(\core_1.decode.oc_alu_mode[6] ),
    .C1(_1790_),
    .X(_1791_));
 sky130_fd_sc_hd__a311o_1 _4888_ (.A1(_0981_),
    .A2(_1772_),
    .A3(_1773_),
    .B1(_1781_),
    .C1(_1791_),
    .X(_1792_));
 sky130_fd_sc_hd__a31o_1 _4889_ (.A1(_1754_),
    .A2(_1762_),
    .A3(_1765_),
    .B1(_1792_),
    .X(_1793_));
 sky130_fd_sc_hd__nor2_1 _4890_ (.A(_1738_),
    .B(_1793_),
    .Y(_1794_));
 sky130_fd_sc_hd__nor2_1 _4891_ (.A(_1688_),
    .B(_1794_),
    .Y(_1795_));
 sky130_fd_sc_hd__a211o_1 _4892_ (.A1(_0959_),
    .A2(\core_1.execute.alu_mul_div.mul_res[1] ),
    .B1(_1795_),
    .C1(_0992_),
    .X(_1796_));
 sky130_fd_sc_hd__a22o_2 _4893_ (.A1(\core_1.execute.alu_mul_div.div_cur[1] ),
    .A2(_0964_),
    .B1(_1687_),
    .B2(_1796_),
    .X(_1797_));
 sky130_fd_sc_hd__inv_2 _4894_ (.A(\core_1.dec_sreg_irt ),
    .Y(_1798_));
 sky130_fd_sc_hd__buf_4 _4895_ (.A(_1798_),
    .X(_1799_));
 sky130_fd_sc_hd__and2_1 _4896_ (.A(_1799_),
    .B(_1153_),
    .X(_1800_));
 sky130_fd_sc_hd__buf_4 _4897_ (.A(_1800_),
    .X(_1801_));
 sky130_fd_sc_hd__and2_1 _4898_ (.A(\core_1.execute.sreg_irq_pc.o_d[1] ),
    .B(\core_1.dec_sreg_irt ),
    .X(_1802_));
 sky130_fd_sc_hd__a221o_1 _4899_ (.A1(_1684_),
    .A2(_1797_),
    .B1(_1801_),
    .B2(net201),
    .C1(_1802_),
    .X(_1803_));
 sky130_fd_sc_hd__and3_1 _4900_ (.A(_1029_),
    .B(_1677_),
    .C(_1803_),
    .X(_1804_));
 sky130_fd_sc_hd__o21a_1 _4901_ (.A1(_1683_),
    .A2(_1804_),
    .B1(_0999_),
    .X(_0187_));
 sky130_fd_sc_hd__or4_1 _4902_ (.A(_0785_),
    .B(net71),
    .C(_0690_),
    .D(_1209_),
    .X(_1805_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _4903_ (.A(_1805_),
    .X(_1806_));
 sky130_fd_sc_hd__nor2_1 _4904_ (.A(_0735_),
    .B(_1806_),
    .Y(_1807_));
 sky130_fd_sc_hd__nor2_1 _4905_ (.A(_1566_),
    .B(_1603_),
    .Y(_1808_));
 sky130_fd_sc_hd__nor2_1 _4906_ (.A(_1808_),
    .B(_1595_),
    .Y(_1809_));
 sky130_fd_sc_hd__a22o_1 _4907_ (.A1(_1204_),
    .A2(_1806_),
    .B1(_1807_),
    .B2(_1809_),
    .X(_0188_));
 sky130_fd_sc_hd__clkbuf_4 _4908_ (.A(_1570_),
    .X(_1810_));
 sky130_fd_sc_hd__nor2_1 _4909_ (.A(_1810_),
    .B(_1808_),
    .Y(_1811_));
 sky130_fd_sc_hd__or4_1 _4910_ (.A(_0735_),
    .B(_1210_),
    .C(_1206_),
    .D(_1811_),
    .X(_1812_));
 sky130_fd_sc_hd__a21bo_1 _4911_ (.A1(_1810_),
    .A2(_1806_),
    .B1_N(_1812_),
    .X(_0189_));
 sky130_fd_sc_hd__nor2_1 _4912_ (.A(_1200_),
    .B(_1206_),
    .Y(_1813_));
 sky130_fd_sc_hd__nor2_1 _4913_ (.A(_1416_),
    .B(_1813_),
    .Y(_1814_));
 sky130_fd_sc_hd__a22o_1 _4914_ (.A1(_1200_),
    .A2(_1806_),
    .B1(_1807_),
    .B2(_1814_),
    .X(_0190_));
 sky130_fd_sc_hd__mux2_1 _4915_ (.A0(\core_1.de_jmp_pred ),
    .A1(\core_1.decode.i_jmp_pred_pass ),
    .S(_0916_),
    .X(_1815_));
 sky130_fd_sc_hd__clkbuf_1 _4916_ (.A(_1815_),
    .X(_0191_));
 sky130_fd_sc_hd__mux2_1 _4917_ (.A0(\core_1.execute.sreg_data_page ),
    .A1(net104),
    .S(_0731_),
    .X(_1816_));
 sky130_fd_sc_hd__and2_1 _4918_ (.A(_1184_),
    .B(_1816_),
    .X(_1817_));
 sky130_fd_sc_hd__clkbuf_1 _4919_ (.A(_1817_),
    .X(_0192_));
 sky130_fd_sc_hd__buf_2 _4920_ (.A(_0729_),
    .X(_1818_));
 sky130_fd_sc_hd__clkbuf_2 _4921_ (.A(_0736_),
    .X(_1819_));
 sky130_fd_sc_hd__clkbuf_2 _4922_ (.A(_0692_),
    .X(_1820_));
 sky130_fd_sc_hd__or4_1 _4923_ (.A(net72),
    .B(_1818_),
    .C(_1819_),
    .D(_1820_),
    .X(_1821_));
 sky130_fd_sc_hd__o211a_1 _4924_ (.A1(\core_1.execute.mem_stage_pc[0] ),
    .A2(_1030_),
    .B1(_1821_),
    .C1(_0999_),
    .X(_0193_));
 sky130_fd_sc_hd__or4_1 _4925_ (.A(net79),
    .B(_1818_),
    .C(_1819_),
    .D(_1820_),
    .X(_1822_));
 sky130_fd_sc_hd__o211a_1 _4926_ (.A1(\core_1.execute.mem_stage_pc[1] ),
    .A2(_1030_),
    .B1(_1822_),
    .C1(_0999_),
    .X(_0194_));
 sky130_fd_sc_hd__or4_1 _4927_ (.A(net80),
    .B(_1818_),
    .C(_1819_),
    .D(_1820_),
    .X(_1823_));
 sky130_fd_sc_hd__o211a_1 _4928_ (.A1(\core_1.execute.mem_stage_pc[2] ),
    .A2(_1030_),
    .B1(_1823_),
    .C1(_0999_),
    .X(_0195_));
 sky130_fd_sc_hd__inv_2 _4929_ (.A(net81),
    .Y(_1824_));
 sky130_fd_sc_hd__buf_4 _4930_ (.A(_1029_),
    .X(_1825_));
 sky130_fd_sc_hd__nand2_1 _4931_ (.A(_1824_),
    .B(_1825_),
    .Y(_1826_));
 sky130_fd_sc_hd__o211a_1 _4932_ (.A1(\core_1.execute.mem_stage_pc[3] ),
    .A2(_1030_),
    .B1(_1826_),
    .C1(_0999_),
    .X(_0196_));
 sky130_fd_sc_hd__inv_2 _4933_ (.A(net82),
    .Y(_1827_));
 sky130_fd_sc_hd__o21ai_1 _4934_ (.A1(\core_1.execute.mem_stage_pc[4] ),
    .A2(_1825_),
    .B1(_1068_),
    .Y(_1828_));
 sky130_fd_sc_hd__a21oi_1 _4935_ (.A1(_1827_),
    .A2(_1071_),
    .B1(_1828_),
    .Y(_0197_));
 sky130_fd_sc_hd__or4_1 _4936_ (.A(net83),
    .B(_1818_),
    .C(_1819_),
    .D(_1820_),
    .X(_1829_));
 sky130_fd_sc_hd__o211a_1 _4937_ (.A1(\core_1.execute.mem_stage_pc[5] ),
    .A2(_1030_),
    .B1(_1829_),
    .C1(_0999_),
    .X(_0198_));
 sky130_fd_sc_hd__inv_2 _4938_ (.A(net84),
    .Y(_1830_));
 sky130_fd_sc_hd__nand2_1 _4939_ (.A(_1830_),
    .B(_1825_),
    .Y(_1831_));
 sky130_fd_sc_hd__o211a_1 _4940_ (.A1(\core_1.execute.mem_stage_pc[6] ),
    .A2(_1030_),
    .B1(_1831_),
    .C1(_0999_),
    .X(_0199_));
 sky130_fd_sc_hd__inv_2 _4941_ (.A(net85),
    .Y(_1832_));
 sky130_fd_sc_hd__nand2_1 _4942_ (.A(_1832_),
    .B(_1825_),
    .Y(_1833_));
 sky130_fd_sc_hd__clkbuf_4 _4943_ (.A(_1307_),
    .X(_1834_));
 sky130_fd_sc_hd__o211a_1 _4944_ (.A1(\core_1.execute.mem_stage_pc[7] ),
    .A2(_1030_),
    .B1(_1833_),
    .C1(_1834_),
    .X(_0200_));
 sky130_fd_sc_hd__or4_1 _4945_ (.A(net86),
    .B(_1818_),
    .C(_1819_),
    .D(_1820_),
    .X(_1835_));
 sky130_fd_sc_hd__o211a_1 _4946_ (.A1(\core_1.execute.mem_stage_pc[8] ),
    .A2(_1030_),
    .B1(_1835_),
    .C1(_1834_),
    .X(_0201_));
 sky130_fd_sc_hd__or4_1 _4947_ (.A(net87),
    .B(_1818_),
    .C(_1819_),
    .D(_1820_),
    .X(_1836_));
 sky130_fd_sc_hd__o211a_1 _4948_ (.A1(\core_1.execute.mem_stage_pc[9] ),
    .A2(_1030_),
    .B1(_1836_),
    .C1(_1834_),
    .X(_0202_));
 sky130_fd_sc_hd__or4_1 _4949_ (.A(net73),
    .B(_1818_),
    .C(_1819_),
    .D(_1820_),
    .X(_1837_));
 sky130_fd_sc_hd__o211a_1 _4950_ (.A1(\core_1.execute.mem_stage_pc[10] ),
    .A2(_1825_),
    .B1(_1837_),
    .C1(_1834_),
    .X(_0203_));
 sky130_fd_sc_hd__or4_1 _4951_ (.A(net74),
    .B(_1818_),
    .C(_1819_),
    .D(_1820_),
    .X(_1838_));
 sky130_fd_sc_hd__o211a_1 _4952_ (.A1(\core_1.execute.mem_stage_pc[11] ),
    .A2(_1825_),
    .B1(_1838_),
    .C1(_1834_),
    .X(_0204_));
 sky130_fd_sc_hd__or4_1 _4953_ (.A(net75),
    .B(_1818_),
    .C(_1819_),
    .D(_1820_),
    .X(_1839_));
 sky130_fd_sc_hd__o211a_1 _4954_ (.A1(\core_1.execute.mem_stage_pc[12] ),
    .A2(_1825_),
    .B1(_1839_),
    .C1(_1834_),
    .X(_0205_));
 sky130_fd_sc_hd__or4_1 _4955_ (.A(net76),
    .B(_1818_),
    .C(_1819_),
    .D(_1820_),
    .X(_1840_));
 sky130_fd_sc_hd__o211a_1 _4956_ (.A1(\core_1.execute.mem_stage_pc[13] ),
    .A2(_1825_),
    .B1(_1840_),
    .C1(_1834_),
    .X(_0206_));
 sky130_fd_sc_hd__or4_1 _4957_ (.A(net77),
    .B(_0729_),
    .C(_0736_),
    .D(_0692_),
    .X(_1841_));
 sky130_fd_sc_hd__o211a_1 _4958_ (.A1(\core_1.execute.mem_stage_pc[14] ),
    .A2(_1825_),
    .B1(_1841_),
    .C1(_1834_),
    .X(_0207_));
 sky130_fd_sc_hd__or4_1 _4959_ (.A(net78),
    .B(_0729_),
    .C(_0736_),
    .D(_0692_),
    .X(_1842_));
 sky130_fd_sc_hd__o211a_1 _4960_ (.A1(\core_1.execute.mem_stage_pc[15] ),
    .A2(_1825_),
    .B1(_1842_),
    .C1(_1834_),
    .X(_0208_));
 sky130_fd_sc_hd__nor2_1 _4961_ (.A(_1128_),
    .B(_0685_),
    .Y(_0209_));
 sky130_fd_sc_hd__nor2_1 _4962_ (.A(_1128_),
    .B(_0683_),
    .Y(_0210_));
 sky130_fd_sc_hd__nor2_1 _4963_ (.A(_1128_),
    .B(_0672_),
    .Y(_0211_));
 sky130_fd_sc_hd__nor2_1 _4964_ (.A(_1128_),
    .B(_0674_),
    .Y(_0212_));
 sky130_fd_sc_hd__nor2_1 _4965_ (.A(_1128_),
    .B(_0678_),
    .Y(_0213_));
 sky130_fd_sc_hd__nor2_1 _4966_ (.A(_1128_),
    .B(_0681_),
    .Y(_0214_));
 sky130_fd_sc_hd__nor2_1 _4967_ (.A(_1122_),
    .B(_0677_),
    .Y(_0215_));
 sky130_fd_sc_hd__nor2_1 _4968_ (.A(_1122_),
    .B(_0673_),
    .Y(_0216_));
 sky130_fd_sc_hd__and3_1 _4969_ (.A(\core_1.execute.trap_flag ),
    .B(_0998_),
    .C(_1071_),
    .X(_1843_));
 sky130_fd_sc_hd__clkbuf_1 _4970_ (.A(_1843_),
    .X(_0217_));
 sky130_fd_sc_hd__and3_1 _4971_ (.A(\core_1.dec_sys ),
    .B(_0998_),
    .C(_1071_),
    .X(_1844_));
 sky130_fd_sc_hd__clkbuf_1 _4972_ (.A(_1844_),
    .X(_0218_));
 sky130_fd_sc_hd__nand2_4 _4973_ (.A(_0662_),
    .B(_1029_),
    .Y(_1845_));
 sky130_fd_sc_hd__buf_6 _4974_ (.A(_1845_),
    .X(_1846_));
 sky130_fd_sc_hd__mux2_1 _4975_ (.A0(\core_1.dec_mem_we ),
    .A1(net159),
    .S(_1846_),
    .X(_1847_));
 sky130_fd_sc_hd__clkbuf_1 _4976_ (.A(_1847_),
    .X(_0219_));
 sky130_fd_sc_hd__a2111o_2 _4977_ (.A1(\core_1.execute.rf.reg_outputs[1][0] ),
    .A2(_1575_),
    .B1(_1627_),
    .C1(_1628_),
    .D1(_1629_),
    .X(_1848_));
 sky130_fd_sc_hd__a21o_2 _4978_ (.A1(_1077_),
    .A2(net184),
    .B1(_1316_),
    .X(_1849_));
 sky130_fd_sc_hd__nor2_1 _4979_ (.A(_1849_),
    .B(_1529_),
    .Y(_1850_));
 sky130_fd_sc_hd__nor2_1 _4980_ (.A(_1317_),
    .B(_1695_),
    .Y(_1851_));
 sky130_fd_sc_hd__nor2_4 _4981_ (.A(_1850_),
    .B(_1851_),
    .Y(_1852_));
 sky130_fd_sc_hd__o21a_1 _4982_ (.A1(_1324_),
    .A2(_1594_),
    .B1(_1852_),
    .X(_1853_));
 sky130_fd_sc_hd__clkinv_4 _4983_ (.A(_1601_),
    .Y(_1854_));
 sky130_fd_sc_hd__and2_1 _4984_ (.A(_1323_),
    .B(_1594_),
    .X(_1855_));
 sky130_fd_sc_hd__nor2_1 _4985_ (.A(_1323_),
    .B(_1594_),
    .Y(_1856_));
 sky130_fd_sc_hd__nor2_2 _4986_ (.A(_1855_),
    .B(_1856_),
    .Y(_1857_));
 sky130_fd_sc_hd__or3_1 _4987_ (.A(_1326_),
    .B(_1854_),
    .C(_1857_),
    .X(_1858_));
 sky130_fd_sc_hd__nand2_1 _4988_ (.A(_1326_),
    .B(_1601_),
    .Y(_1859_));
 sky130_fd_sc_hd__inv_2 _4989_ (.A(_1859_),
    .Y(_1860_));
 sky130_fd_sc_hd__nor2_1 _4990_ (.A(_1326_),
    .B(_1601_),
    .Y(_1861_));
 sky130_fd_sc_hd__nor2_2 _4991_ (.A(_1860_),
    .B(_1861_),
    .Y(_1862_));
 sky130_fd_sc_hd__o21a_1 _4992_ (.A1(_1330_),
    .A2(_1580_),
    .B1(_1862_),
    .X(_1863_));
 sky130_fd_sc_hd__or3_1 _4993_ (.A(_1330_),
    .B(_1580_),
    .C(_1862_),
    .X(_1864_));
 sky130_fd_sc_hd__and2b_1 _4994_ (.A_N(_1863_),
    .B(_1864_),
    .X(_1865_));
 sky130_fd_sc_hd__a21o_2 _4995_ (.A1(_1077_),
    .A2(net180),
    .B1(_1334_),
    .X(_1866_));
 sky130_fd_sc_hd__or2_1 _4996_ (.A(_1866_),
    .B(_1586_),
    .X(_1867_));
 sky130_fd_sc_hd__inv_2 _4997_ (.A(_1867_),
    .Y(_1868_));
 sky130_fd_sc_hd__and2_1 _4998_ (.A(_1866_),
    .B(_1586_),
    .X(_1869_));
 sky130_fd_sc_hd__nor2_2 _4999_ (.A(_1868_),
    .B(_1869_),
    .Y(_1870_));
 sky130_fd_sc_hd__o21a_1 _5000_ (.A1(_1341_),
    .A2(_1543_),
    .B1(_1870_),
    .X(_1871_));
 sky130_fd_sc_hd__nor3_1 _5001_ (.A(_1341_),
    .B(_1543_),
    .C(_1870_),
    .Y(_1872_));
 sky130_fd_sc_hd__nor2_1 _5002_ (.A(_1871_),
    .B(_1872_),
    .Y(_1873_));
 sky130_fd_sc_hd__inv_2 _5003_ (.A(_1564_),
    .Y(_1874_));
 sky130_fd_sc_hd__nor2_2 _5004_ (.A(_1343_),
    .B(_1535_),
    .Y(_1875_));
 sky130_fd_sc_hd__and2_1 _5005_ (.A(_1343_),
    .B(_1535_),
    .X(_1876_));
 sky130_fd_sc_hd__or2_1 _5006_ (.A(_1875_),
    .B(_1876_),
    .X(_1877_));
 sky130_fd_sc_hd__a21oi_1 _5007_ (.A1(_1347_),
    .A2(_1874_),
    .B1(_1877_),
    .Y(_1878_));
 sky130_fd_sc_hd__and3_1 _5008_ (.A(_1347_),
    .B(_1874_),
    .C(_1877_),
    .X(_1879_));
 sky130_fd_sc_hd__or2_1 _5009_ (.A(_1878_),
    .B(_1879_),
    .X(_1880_));
 sky130_fd_sc_hd__and2_2 _5010_ (.A(_1697_),
    .B(_1556_),
    .X(_1881_));
 sky130_fd_sc_hd__nor2_1 _5011_ (.A(_1697_),
    .B(_1556_),
    .Y(_1882_));
 sky130_fd_sc_hd__nor2_1 _5012_ (.A(_1881_),
    .B(_1882_),
    .Y(_1883_));
 sky130_fd_sc_hd__o21a_1 _5013_ (.A1(_1352_),
    .A2(_1658_),
    .B1(_1883_),
    .X(_1884_));
 sky130_fd_sc_hd__inv_2 _5014_ (.A(_1658_),
    .Y(_1885_));
 sky130_fd_sc_hd__o211a_1 _5015_ (.A1(_1881_),
    .A2(_1882_),
    .B1(_1351_),
    .C1(_1885_),
    .X(_1886_));
 sky130_fd_sc_hd__nor2_1 _5016_ (.A(_1884_),
    .B(_1886_),
    .Y(_1887_));
 sky130_fd_sc_hd__nand2_1 _5017_ (.A(_1351_),
    .B(_1658_),
    .Y(_1888_));
 sky130_fd_sc_hd__or2_1 _5018_ (.A(_1351_),
    .B(_1657_),
    .X(_1889_));
 sky130_fd_sc_hd__and2_1 _5019_ (.A(_1888_),
    .B(_1889_),
    .X(_1890_));
 sky130_fd_sc_hd__nor2_1 _5020_ (.A(_1665_),
    .B(_1890_),
    .Y(_1891_));
 sky130_fd_sc_hd__o21a_1 _5021_ (.A1(_1357_),
    .A2(_1665_),
    .B1(_1890_),
    .X(_1892_));
 sky130_fd_sc_hd__a21oi_2 _5022_ (.A1(_1696_),
    .A2(_1891_),
    .B1(_1892_),
    .Y(_1893_));
 sky130_fd_sc_hd__xnor2_2 _5023_ (.A(_1357_),
    .B(_1664_),
    .Y(_1894_));
 sky130_fd_sc_hd__o21ai_1 _5024_ (.A1(_1364_),
    .A2(_1724_),
    .B1(_1894_),
    .Y(_1895_));
 sky130_fd_sc_hd__or3_1 _5025_ (.A(_1364_),
    .B(_1724_),
    .C(_1894_),
    .X(_1896_));
 sky130_fd_sc_hd__and2_1 _5026_ (.A(_1895_),
    .B(_1896_),
    .X(_1897_));
 sky130_fd_sc_hd__nand2_1 _5027_ (.A(_1372_),
    .B(_1727_),
    .Y(_1898_));
 sky130_fd_sc_hd__a21o_1 _5028_ (.A1(_1690_),
    .A2(_1770_),
    .B1(_1769_),
    .X(_1899_));
 sky130_fd_sc_hd__nor2_1 _5029_ (.A(_1372_),
    .B(_1727_),
    .Y(_1900_));
 sky130_fd_sc_hd__nor2_1 _5030_ (.A(_1368_),
    .B(_1643_),
    .Y(_1901_));
 sky130_fd_sc_hd__nand2_1 _5031_ (.A(_1368_),
    .B(_1643_),
    .Y(_1902_));
 sky130_fd_sc_hd__and2b_1 _5032_ (.A_N(_1901_),
    .B(_1902_),
    .X(_1903_));
 sky130_fd_sc_hd__a211o_1 _5033_ (.A1(_1898_),
    .A2(_1899_),
    .B1(_1900_),
    .C1(_1903_),
    .X(_1904_));
 sky130_fd_sc_hd__xnor2_4 _5034_ (.A(_1361_),
    .B(_1650_),
    .Y(_1905_));
 sky130_fd_sc_hd__nand2_1 _5035_ (.A(_1689_),
    .B(_1643_),
    .Y(_1906_));
 sky130_fd_sc_hd__nand2_1 _5036_ (.A(_1905_),
    .B(_1906_),
    .Y(_1907_));
 sky130_fd_sc_hd__or2_1 _5037_ (.A(_1905_),
    .B(_1906_),
    .X(_1908_));
 sky130_fd_sc_hd__and2_1 _5038_ (.A(_1907_),
    .B(_1908_),
    .X(_1909_));
 sky130_fd_sc_hd__a21boi_1 _5039_ (.A1(_1895_),
    .A2(_1907_),
    .B1_N(_1896_),
    .Y(_1910_));
 sky130_fd_sc_hd__a31o_2 _5040_ (.A1(_1897_),
    .A2(_1904_),
    .A3(_1909_),
    .B1(_1910_),
    .X(_1911_));
 sky130_fd_sc_hd__o21ba_1 _5041_ (.A1(_1884_),
    .A2(_1892_),
    .B1_N(_1886_),
    .X(_1912_));
 sky130_fd_sc_hd__a31oi_4 _5042_ (.A1(_1887_),
    .A2(_1893_),
    .A3(_1911_),
    .B1(_1912_),
    .Y(_1913_));
 sky130_fd_sc_hd__nand2_2 _5043_ (.A(_1347_),
    .B(_1564_),
    .Y(_1914_));
 sky130_fd_sc_hd__or2_1 _5044_ (.A(_1347_),
    .B(_1563_),
    .X(_1915_));
 sky130_fd_sc_hd__and2_2 _5045_ (.A(_1914_),
    .B(_1915_),
    .X(_1916_));
 sky130_fd_sc_hd__o21ai_2 _5046_ (.A1(_1349_),
    .A2(_1557_),
    .B1(_1916_),
    .Y(_1917_));
 sky130_fd_sc_hd__or3_1 _5047_ (.A(_1349_),
    .B(_1556_),
    .C(_1916_),
    .X(_1918_));
 sky130_fd_sc_hd__nand2_1 _5048_ (.A(_1917_),
    .B(_1918_),
    .Y(_1919_));
 sky130_fd_sc_hd__o21ba_1 _5049_ (.A1(_1879_),
    .A2(_1917_),
    .B1_N(_1878_),
    .X(_1920_));
 sky130_fd_sc_hd__o31ai_4 _5050_ (.A1(_1880_),
    .A2(_1913_),
    .A3(_1919_),
    .B1(_1920_),
    .Y(_1921_));
 sky130_fd_sc_hd__and2_1 _5051_ (.A(_1340_),
    .B(_1542_),
    .X(_1922_));
 sky130_fd_sc_hd__nor2_1 _5052_ (.A(_1340_),
    .B(_1543_),
    .Y(_1923_));
 sky130_fd_sc_hd__or2_2 _5053_ (.A(_1922_),
    .B(_1923_),
    .X(_1924_));
 sky130_fd_sc_hd__a21oi_1 _5054_ (.A1(_1343_),
    .A2(_1536_),
    .B1(_1924_),
    .Y(_1925_));
 sky130_fd_sc_hd__and3_1 _5055_ (.A(_1343_),
    .B(_1536_),
    .C(_1924_),
    .X(_1926_));
 sky130_fd_sc_hd__nor2_1 _5056_ (.A(_1925_),
    .B(_1926_),
    .Y(_1927_));
 sky130_fd_sc_hd__o21ba_1 _5057_ (.A1(_1871_),
    .A2(_1925_),
    .B1_N(_1872_),
    .X(_1928_));
 sky130_fd_sc_hd__a31o_1 _5058_ (.A1(_1873_),
    .A2(_1921_),
    .A3(_1927_),
    .B1(_1928_),
    .X(_1929_));
 sky130_fd_sc_hd__and2_2 _5059_ (.A(_1329_),
    .B(_1579_),
    .X(_1930_));
 sky130_fd_sc_hd__nor2_1 _5060_ (.A(_1329_),
    .B(_1580_),
    .Y(_1931_));
 sky130_fd_sc_hd__nor2_2 _5061_ (.A(_1930_),
    .B(_1931_),
    .Y(_1932_));
 sky130_fd_sc_hd__nor2_1 _5062_ (.A(_1586_),
    .B(_1932_),
    .Y(_1933_));
 sky130_fd_sc_hd__o21a_1 _5063_ (.A1(_1335_),
    .A2(_1586_),
    .B1(_1932_),
    .X(_1934_));
 sky130_fd_sc_hd__a21oi_2 _5064_ (.A1(_1866_),
    .A2(_1933_),
    .B1(_1934_),
    .Y(_1935_));
 sky130_fd_sc_hd__a21o_1 _5065_ (.A1(_1864_),
    .A2(_1934_),
    .B1(_1863_),
    .X(_1936_));
 sky130_fd_sc_hd__a31o_1 _5066_ (.A1(_1865_),
    .A2(_1929_),
    .A3(_1935_),
    .B1(_1936_),
    .X(_1937_));
 sky130_fd_sc_hd__o21ai_1 _5067_ (.A1(_1326_),
    .A2(_1854_),
    .B1(_1857_),
    .Y(_1938_));
 sky130_fd_sc_hd__a21bo_1 _5068_ (.A1(_1858_),
    .A2(_1937_),
    .B1_N(_1938_),
    .X(_1939_));
 sky130_fd_sc_hd__nor3_1 _5069_ (.A(_1324_),
    .B(_1594_),
    .C(_1852_),
    .Y(_1940_));
 sky130_fd_sc_hd__a21oi_1 _5070_ (.A1(_1849_),
    .A2(_1695_),
    .B1(_1940_),
    .Y(_1941_));
 sky130_fd_sc_hd__o21ai_1 _5071_ (.A1(_1853_),
    .A2(_1939_),
    .B1(_1941_),
    .Y(_1942_));
 sky130_fd_sc_hd__or2_1 _5072_ (.A(_1869_),
    .B(_1922_),
    .X(_1943_));
 sky130_fd_sc_hd__inv_2 _5073_ (.A(_1876_),
    .Y(_1944_));
 sky130_fd_sc_hd__nand2_1 _5074_ (.A(_1384_),
    .B(_1727_),
    .Y(_1945_));
 sky130_fd_sc_hd__nor2_1 _5075_ (.A(_1383_),
    .B(_1727_),
    .Y(_1946_));
 sky130_fd_sc_hd__a211o_1 _5076_ (.A1(_1782_),
    .A2(_1779_),
    .B1(_1946_),
    .C1(_1775_),
    .X(_1947_));
 sky130_fd_sc_hd__a31o_1 _5077_ (.A1(_1902_),
    .A2(_1945_),
    .A3(_1947_),
    .B1(_1901_),
    .X(_1948_));
 sky130_fd_sc_hd__and2_1 _5078_ (.A(_1894_),
    .B(_1905_),
    .X(_1949_));
 sky130_fd_sc_hd__and4_1 _5079_ (.A(_1883_),
    .B(_1890_),
    .C(_1948_),
    .D(_1949_),
    .X(_1950_));
 sky130_fd_sc_hd__nor2_1 _5080_ (.A(_1352_),
    .B(_1885_),
    .Y(_1951_));
 sky130_fd_sc_hd__and2_1 _5081_ (.A(_1696_),
    .B(_1664_),
    .X(_1952_));
 sky130_fd_sc_hd__nor2_1 _5082_ (.A(_1364_),
    .B(_1650_),
    .Y(_1953_));
 sky130_fd_sc_hd__or2_1 _5083_ (.A(_1696_),
    .B(_1664_),
    .X(_1954_));
 sky130_fd_sc_hd__o21a_1 _5084_ (.A1(_1952_),
    .A2(_1953_),
    .B1(_1954_),
    .X(_1955_));
 sky130_fd_sc_hd__or2_1 _5085_ (.A(_1697_),
    .B(_1556_),
    .X(_1956_));
 sky130_fd_sc_hd__o211a_1 _5086_ (.A1(_1951_),
    .A2(_1955_),
    .B1(_1889_),
    .C1(_1956_),
    .X(_1957_));
 sky130_fd_sc_hd__o31ai_4 _5087_ (.A1(_1881_),
    .A2(_1950_),
    .A3(_1957_),
    .B1(_1916_),
    .Y(_1958_));
 sky130_fd_sc_hd__a311oi_4 _5088_ (.A1(_1944_),
    .A2(_1914_),
    .A3(_1958_),
    .B1(_1924_),
    .C1(_1875_),
    .Y(_1959_));
 sky130_fd_sc_hd__o211a_1 _5089_ (.A1(_1943_),
    .A2(_1959_),
    .B1(_1867_),
    .C1(_1932_),
    .X(_1960_));
 sky130_fd_sc_hd__o311a_2 _5090_ (.A1(_1861_),
    .A2(_1930_),
    .A3(_1960_),
    .B1(_1859_),
    .C1(_1857_),
    .X(_1961_));
 sky130_fd_sc_hd__nand2_1 _5091_ (.A(_1317_),
    .B(_1695_),
    .Y(_1962_));
 sky130_fd_sc_hd__o311a_1 _5092_ (.A1(_1851_),
    .A2(_1855_),
    .A3(_1961_),
    .B1(_1962_),
    .C1(_0966_),
    .X(_1963_));
 sky130_fd_sc_hd__xnor2_1 _5093_ (.A(_1696_),
    .B(_1743_),
    .Y(_1964_));
 sky130_fd_sc_hd__or2_1 _5094_ (.A(\core_1.decode.oc_alu_mode[12] ),
    .B(_1658_),
    .X(_1965_));
 sky130_fd_sc_hd__nand2_1 _5095_ (.A(_1748_),
    .B(_1965_),
    .Y(_1966_));
 sky130_fd_sc_hd__o21a_1 _5096_ (.A1(\core_1.decode.oc_alu_mode[12] ),
    .A2(_1665_),
    .B1(_1747_),
    .X(_1967_));
 sky130_fd_sc_hd__nor2_1 _5097_ (.A(_1418_),
    .B(_1967_),
    .Y(_1968_));
 sky130_fd_sc_hd__a21o_1 _5098_ (.A1(_1418_),
    .A2(_1966_),
    .B1(_1968_),
    .X(_1969_));
 sky130_fd_sc_hd__o21ai_1 _5099_ (.A1(_1750_),
    .A2(_1564_),
    .B1(_1747_),
    .Y(_1970_));
 sky130_fd_sc_hd__nor2_1 _5100_ (.A(\core_1.decode.oc_alu_mode[12] ),
    .B(_1557_),
    .Y(_1971_));
 sky130_fd_sc_hd__or4_1 _5101_ (.A(_1417_),
    .B(_1745_),
    .C(_1746_),
    .D(_1971_),
    .X(_1972_));
 sky130_fd_sc_hd__o21a_1 _5102_ (.A1(_1692_),
    .A2(_1970_),
    .B1(_1972_),
    .X(_1973_));
 sky130_fd_sc_hd__clkinv_2 _5103_ (.A(_1727_),
    .Y(_1974_));
 sky130_fd_sc_hd__o21ai_1 _5104_ (.A1(_1750_),
    .A2(_1974_),
    .B1(_1747_),
    .Y(_1975_));
 sky130_fd_sc_hd__mux2_1 _5105_ (.A0(_1752_),
    .A1(_1975_),
    .S(_1418_),
    .X(_1976_));
 sky130_fd_sc_hd__nand2_1 _5106_ (.A(_1742_),
    .B(_1643_),
    .Y(_1977_));
 sky130_fd_sc_hd__nand2_1 _5107_ (.A(_1748_),
    .B(_1977_),
    .Y(_1978_));
 sky130_fd_sc_hd__o21a_1 _5108_ (.A1(\core_1.decode.oc_alu_mode[12] ),
    .A2(_1724_),
    .B1(_1747_),
    .X(_1979_));
 sky130_fd_sc_hd__nor2_1 _5109_ (.A(_1692_),
    .B(_1979_),
    .Y(_1980_));
 sky130_fd_sc_hd__a21o_1 _5110_ (.A1(_1692_),
    .A2(_1978_),
    .B1(_1980_),
    .X(_1981_));
 sky130_fd_sc_hd__a21oi_4 _5111_ (.A1(_0988_),
    .A2(_1728_),
    .B1(_1739_),
    .Y(_1982_));
 sky130_fd_sc_hd__xnor2_4 _5112_ (.A(_1384_),
    .B(_1763_),
    .Y(_1983_));
 sky130_fd_sc_hd__mux4_1 _5113_ (.A0(_1969_),
    .A1(_1973_),
    .A2(_1976_),
    .A3(_1981_),
    .S0(_1982_),
    .S1(_1983_),
    .X(_1984_));
 sky130_fd_sc_hd__nand2_1 _5114_ (.A(_1761_),
    .B(_1984_),
    .Y(_1985_));
 sky130_fd_sc_hd__o21ai_1 _5115_ (.A1(_1750_),
    .A2(_1535_),
    .B1(_1747_),
    .Y(_1986_));
 sky130_fd_sc_hd__o21ai_1 _5116_ (.A1(_1750_),
    .A2(_1543_),
    .B1(_1747_),
    .Y(_1987_));
 sky130_fd_sc_hd__mux2_1 _5117_ (.A0(_1986_),
    .A1(_1987_),
    .S(_1418_),
    .X(_1988_));
 sky130_fd_sc_hd__o21ai_1 _5118_ (.A1(_1750_),
    .A2(_1586_),
    .B1(_1747_),
    .Y(_1989_));
 sky130_fd_sc_hd__o21ai_1 _5119_ (.A1(_1750_),
    .A2(_1580_),
    .B1(_1747_),
    .Y(_1990_));
 sky130_fd_sc_hd__mux2_1 _5120_ (.A0(_1989_),
    .A1(_1990_),
    .S(_1418_),
    .X(_1991_));
 sky130_fd_sc_hd__mux2_1 _5121_ (.A0(_1988_),
    .A1(_1991_),
    .S(_1982_),
    .X(_1992_));
 sky130_fd_sc_hd__o21ai_1 _5122_ (.A1(_1750_),
    .A2(_1854_),
    .B1(_1748_),
    .Y(_1993_));
 sky130_fd_sc_hd__o21ai_1 _5123_ (.A1(_1750_),
    .A2(_1593_),
    .B1(_1748_),
    .Y(_1994_));
 sky130_fd_sc_hd__mux2_1 _5124_ (.A0(_1993_),
    .A1(_1994_),
    .S(_1418_),
    .X(_1995_));
 sky130_fd_sc_hd__nor2_1 _5125_ (.A(_1695_),
    .B(_1745_),
    .Y(_1996_));
 sky130_fd_sc_hd__a21oi_1 _5126_ (.A1(_1692_),
    .A2(_1996_),
    .B1(_1740_),
    .Y(_1997_));
 sky130_fd_sc_hd__a211o_1 _5127_ (.A1(_1740_),
    .A2(_1995_),
    .B1(_1997_),
    .C1(_1983_),
    .X(_1998_));
 sky130_fd_sc_hd__buf_2 _5128_ (.A(_1760_),
    .X(_1999_));
 sky130_fd_sc_hd__o211ai_1 _5129_ (.A1(_1764_),
    .A2(_1992_),
    .B1(_1998_),
    .C1(_1999_),
    .Y(_2000_));
 sky130_fd_sc_hd__nor2_1 _5130_ (.A(_1758_),
    .B(_1749_),
    .Y(_2001_));
 sky130_fd_sc_hd__and3b_1 _5131_ (.A_N(_1756_),
    .B(_1999_),
    .C(_2001_),
    .X(_2002_));
 sky130_fd_sc_hd__a31o_1 _5132_ (.A1(_1756_),
    .A2(_1985_),
    .A3(_2000_),
    .B1(_2002_),
    .X(_2003_));
 sky130_fd_sc_hd__and3_1 _5133_ (.A(\core_1.decode.oc_alu_mode[13] ),
    .B(_1964_),
    .C(_2003_),
    .X(_2004_));
 sky130_fd_sc_hd__a211o_2 _5134_ (.A1(_0981_),
    .A2(_1942_),
    .B1(_1963_),
    .C1(_2004_),
    .X(_2005_));
 sky130_fd_sc_hd__nor2_1 _5135_ (.A(_1849_),
    .B(_2005_),
    .Y(_2006_));
 sky130_fd_sc_hd__xnor2_1 _5136_ (.A(_1848_),
    .B(_2006_),
    .Y(_2007_));
 sky130_fd_sc_hd__and2_1 _5137_ (.A(_0662_),
    .B(_1029_),
    .X(_2008_));
 sky130_fd_sc_hd__buf_6 _5138_ (.A(_2008_),
    .X(_2009_));
 sky130_fd_sc_hd__mux2_1 _5139_ (.A0(\core_1.ew_addr_high[0] ),
    .A1(_2007_),
    .S(_2009_),
    .X(_2010_));
 sky130_fd_sc_hd__clkbuf_1 _5140_ (.A(_2010_),
    .X(_0220_));
 sky130_fd_sc_hd__o21ba_1 _5141_ (.A1(_1849_),
    .A2(_1848_),
    .B1_N(_2005_),
    .X(_2011_));
 sky130_fd_sc_hd__and2_1 _5142_ (.A(\core_1.execute.rf.reg_outputs[1][1] ),
    .B(_1575_),
    .X(_2012_));
 sky130_fd_sc_hd__or3_1 _5143_ (.A(_1620_),
    .B(_1621_),
    .C(_1622_),
    .X(_2013_));
 sky130_fd_sc_hd__or3_2 _5144_ (.A(_2012_),
    .B(_2013_),
    .C(_1848_),
    .X(_2014_));
 sky130_fd_sc_hd__o21ai_1 _5145_ (.A1(_2012_),
    .A2(_2013_),
    .B1(_1848_),
    .Y(_2015_));
 sky130_fd_sc_hd__nand2_1 _5146_ (.A(_2014_),
    .B(_2015_),
    .Y(_2016_));
 sky130_fd_sc_hd__xnor2_1 _5147_ (.A(_2011_),
    .B(_2016_),
    .Y(_2017_));
 sky130_fd_sc_hd__mux2_1 _5148_ (.A0(net132),
    .A1(_2017_),
    .S(_2009_),
    .X(_2018_));
 sky130_fd_sc_hd__clkbuf_1 _5149_ (.A(_2018_),
    .X(_0221_));
 sky130_fd_sc_hd__clkinv_2 _5150_ (.A(_2014_),
    .Y(_2019_));
 sky130_fd_sc_hd__or2_1 _5151_ (.A(_1317_),
    .B(_2005_),
    .X(_2020_));
 sky130_fd_sc_hd__clkbuf_2 _5152_ (.A(_2020_),
    .X(_2021_));
 sky130_fd_sc_hd__a2bb2o_1 _5153_ (.A1_N(_2005_),
    .A2_N(_2019_),
    .B1(_2015_),
    .B2(_2021_),
    .X(_2022_));
 sky130_fd_sc_hd__a211o_1 _5154_ (.A1(\core_1.execute.rf.reg_outputs[1][2] ),
    .A2(_1575_),
    .B1(_1609_),
    .C1(_1611_),
    .X(_2023_));
 sky130_fd_sc_hd__or2_4 _5155_ (.A(_1610_),
    .B(_2023_),
    .X(_2024_));
 sky130_fd_sc_hd__nor2_1 _5156_ (.A(_2022_),
    .B(_2024_),
    .Y(_2025_));
 sky130_fd_sc_hd__and2_1 _5157_ (.A(_0662_),
    .B(_1071_),
    .X(_2026_));
 sky130_fd_sc_hd__buf_2 _5158_ (.A(_2026_),
    .X(_0228_));
 sky130_fd_sc_hd__a21bo_1 _5159_ (.A1(_2022_),
    .A2(_2024_),
    .B1_N(_0228_),
    .X(_2027_));
 sky130_fd_sc_hd__o22a_1 _5160_ (.A1(net133),
    .A2(_2009_),
    .B1(_2025_),
    .B2(_2027_),
    .X(_0222_));
 sky130_fd_sc_hd__nand3b_1 _5161_ (.A_N(_2015_),
    .B(_2024_),
    .C(_2005_),
    .Y(_2028_));
 sky130_fd_sc_hd__o31a_1 _5162_ (.A1(_2021_),
    .A2(_2014_),
    .A3(_2024_),
    .B1(_2028_),
    .X(_2029_));
 sky130_fd_sc_hd__a21oi_2 _5163_ (.A1(\core_1.execute.rf.reg_outputs[1][3] ),
    .A2(_1575_),
    .B1(_1639_),
    .Y(_2030_));
 sky130_fd_sc_hd__xor2_1 _5164_ (.A(_2029_),
    .B(_2030_),
    .X(_2031_));
 sky130_fd_sc_hd__mux2_1 _5165_ (.A0(net134),
    .A1(_2031_),
    .S(_2009_),
    .X(_2032_));
 sky130_fd_sc_hd__clkbuf_1 _5166_ (.A(_2032_),
    .X(_0223_));
 sky130_fd_sc_hd__a21o_1 _5167_ (.A1(\core_1.execute.rf.reg_outputs[1][4] ),
    .A2(_1575_),
    .B1(_1648_),
    .X(_2033_));
 sky130_fd_sc_hd__or2_1 _5168_ (.A(_2028_),
    .B(_2030_),
    .X(_2034_));
 sky130_fd_sc_hd__or4b_1 _5169_ (.A(_2021_),
    .B(_2014_),
    .C(_2024_),
    .D_N(_2030_),
    .X(_2035_));
 sky130_fd_sc_hd__nand2_1 _5170_ (.A(_2034_),
    .B(_2035_),
    .Y(_2036_));
 sky130_fd_sc_hd__xor2_1 _5171_ (.A(_2033_),
    .B(_2036_),
    .X(_2037_));
 sky130_fd_sc_hd__mux2_1 _5172_ (.A0(net135),
    .A1(_2037_),
    .S(_2009_),
    .X(_2038_));
 sky130_fd_sc_hd__clkbuf_1 _5173_ (.A(_2038_),
    .X(_0224_));
 sky130_fd_sc_hd__a21o_1 _5174_ (.A1(\core_1.execute.rf.reg_outputs[1][5] ),
    .A2(_1575_),
    .B1(_1660_),
    .X(_2039_));
 sky130_fd_sc_hd__mux2_1 _5175_ (.A0(_2035_),
    .A1(_2034_),
    .S(_2033_),
    .X(_2040_));
 sky130_fd_sc_hd__xnor2_1 _5176_ (.A(_2039_),
    .B(_2040_),
    .Y(_2041_));
 sky130_fd_sc_hd__mux2_1 _5177_ (.A0(net136),
    .A1(_2041_),
    .S(_2009_),
    .X(_2042_));
 sky130_fd_sc_hd__clkbuf_1 _5178_ (.A(_2042_),
    .X(_0225_));
 sky130_fd_sc_hd__a21o_1 _5179_ (.A1(\core_1.execute.rf.reg_outputs[1][6] ),
    .A2(_1575_),
    .B1(_1655_),
    .X(_2043_));
 sky130_fd_sc_hd__xor2_1 _5180_ (.A(_2021_),
    .B(_2039_),
    .X(_2044_));
 sky130_fd_sc_hd__or2_1 _5181_ (.A(_2040_),
    .B(_2044_),
    .X(_2045_));
 sky130_fd_sc_hd__xnor2_1 _5182_ (.A(_2043_),
    .B(_2045_),
    .Y(_2046_));
 sky130_fd_sc_hd__mux2_1 _5183_ (.A0(net137),
    .A1(_2046_),
    .S(_2009_),
    .X(_2047_));
 sky130_fd_sc_hd__clkbuf_1 _5184_ (.A(_2047_),
    .X(_0226_));
 sky130_fd_sc_hd__a21oi_2 _5185_ (.A1(\core_1.execute.rf.reg_outputs[1][7] ),
    .A2(_1575_),
    .B1(_1550_),
    .Y(_2048_));
 sky130_fd_sc_hd__xor2_1 _5186_ (.A(_2021_),
    .B(_2043_),
    .X(_2049_));
 sky130_fd_sc_hd__or4_1 _5187_ (.A(_2040_),
    .B(_2044_),
    .C(_2048_),
    .D(_2049_),
    .X(_2050_));
 sky130_fd_sc_hd__o31ai_1 _5188_ (.A1(_2040_),
    .A2(_2044_),
    .A3(_2049_),
    .B1(_2048_),
    .Y(_2051_));
 sky130_fd_sc_hd__and2_1 _5189_ (.A(net138),
    .B(_1846_),
    .X(_2052_));
 sky130_fd_sc_hd__a31o_1 _5190_ (.A1(_2009_),
    .A2(_2050_),
    .A3(_2051_),
    .B1(_2052_),
    .X(_0227_));
 sky130_fd_sc_hd__or2_2 _5191_ (.A(\core_1.execute.sreg_irq_pc.o_d[0] ),
    .B(_1798_),
    .X(_2053_));
 sky130_fd_sc_hd__inv_2 _5192_ (.A(\core_1.dec_sreg_jal_over ),
    .Y(_2054_));
 sky130_fd_sc_hd__or2_1 _5193_ (.A(net211),
    .B(_2054_),
    .X(_2055_));
 sky130_fd_sc_hd__and4_1 _5194_ (.A(net185),
    .B(net178),
    .C(_1053_),
    .D(_1054_),
    .X(_2056_));
 sky130_fd_sc_hd__and2_4 _5195_ (.A(_1052_),
    .B(_2056_),
    .X(_2057_));
 sky130_fd_sc_hd__and3_1 _5196_ (.A(net211),
    .B(_1052_),
    .C(_1056_),
    .X(_2058_));
 sky130_fd_sc_hd__and3b_1 _5197_ (.A_N(net187),
    .B(net186),
    .C(_1051_),
    .X(_2059_));
 sky130_fd_sc_hd__and4b_1 _5198_ (.A_N(net178),
    .B(_1053_),
    .C(_1054_),
    .D(net185),
    .X(_2060_));
 sky130_fd_sc_hd__and3_1 _5199_ (.A(\core_1.execute.sreg_scratch.o_d[0] ),
    .B(_2059_),
    .C(_2060_),
    .X(_2061_));
 sky130_fd_sc_hd__and3_1 _5200_ (.A(\core_1.execute.sreg_irq_flags.o_d[0] ),
    .B(_1160_),
    .C(_2059_),
    .X(_2062_));
 sky130_fd_sc_hd__a2111o_1 _5201_ (.A1(\core_1.execute.sreg_irq_pc.o_d[0] ),
    .A2(_2057_),
    .B1(_2058_),
    .C1(_2061_),
    .D1(_2062_),
    .X(_2063_));
 sky130_fd_sc_hd__and3_1 _5202_ (.A(net187),
    .B(net186),
    .C(_1051_),
    .X(_2064_));
 sky130_fd_sc_hd__and2_2 _5203_ (.A(_1160_),
    .B(_2064_),
    .X(_2065_));
 sky130_fd_sc_hd__buf_2 _5204_ (.A(_2059_),
    .X(_2066_));
 sky130_fd_sc_hd__a21o_1 _5205_ (.A1(_2066_),
    .A2(_2056_),
    .B1(\core_1.dec_sreg_jal_over ),
    .X(_2067_));
 sky130_fd_sc_hd__and4_1 _5206_ (.A(net187),
    .B(_1050_),
    .C(_1051_),
    .D(_1055_),
    .X(_2068_));
 sky130_fd_sc_hd__and3_1 _5207_ (.A(\core_1.execute.alu_flag_reg.o_d[0] ),
    .B(_1056_),
    .C(_2066_),
    .X(_2069_));
 sky130_fd_sc_hd__a2111o_1 _5208_ (.A1(\core_1.execute.pc_high_buff_out[0] ),
    .A2(_2065_),
    .B1(_2067_),
    .C1(_2068_),
    .D1(_2069_),
    .X(_2070_));
 sky130_fd_sc_hd__and4_2 _5209_ (.A(net187),
    .B(_1050_),
    .C(_1051_),
    .D(_1159_),
    .X(_2071_));
 sky130_fd_sc_hd__and3_1 _5210_ (.A(net106),
    .B(_1052_),
    .C(_2060_),
    .X(_2072_));
 sky130_fd_sc_hd__and3_1 _5211_ (.A(\core_1.execute.pc_high_out[0] ),
    .B(_1056_),
    .C(_2064_),
    .X(_2073_));
 sky130_fd_sc_hd__and3_1 _5212_ (.A(\core_1.execute.sreg_priv_control.o_d[0] ),
    .B(_1052_),
    .C(_1160_),
    .X(_2074_));
 sky130_fd_sc_hd__a2111o_1 _5213_ (.A1(net1),
    .A2(_2071_),
    .B1(_2072_),
    .C1(_2073_),
    .D1(_2074_),
    .X(_2075_));
 sky130_fd_sc_hd__or3_1 _5214_ (.A(_2063_),
    .B(_2070_),
    .C(_2075_),
    .X(_2076_));
 sky130_fd_sc_hd__a21o_1 _5215_ (.A1(_2055_),
    .A2(_2076_),
    .B1(\core_1.dec_sreg_irt ),
    .X(_2077_));
 sky130_fd_sc_hd__nand2_1 _5216_ (.A(_2053_),
    .B(_2077_),
    .Y(_2078_));
 sky130_fd_sc_hd__xnor2_1 _5217_ (.A(\core_1.dec_sreg_jal_over ),
    .B(_2078_),
    .Y(_2079_));
 sky130_fd_sc_hd__a21o_1 _5218_ (.A1(\core_1.execute.alu_mul_div.div_res[0] ),
    .A2(_0992_),
    .B1(\core_1.execute.alu_mul_div.i_mod ),
    .X(_2080_));
 sky130_fd_sc_hd__inv_2 _5219_ (.A(_0958_),
    .Y(_2081_));
 sky130_fd_sc_hd__o2bb2a_1 _5220_ (.A1_N(_1535_),
    .A2_N(_1712_),
    .B1(_1709_),
    .B2(_1874_),
    .X(_2082_));
 sky130_fd_sc_hd__nand2_1 _5221_ (.A(_1692_),
    .B(_1586_),
    .Y(_2083_));
 sky130_fd_sc_hd__o2bb2a_1 _5222_ (.A1_N(_1543_),
    .A2_N(_1713_),
    .B1(_2083_),
    .B2(_1703_),
    .X(_2084_));
 sky130_fd_sc_hd__a22oi_2 _5223_ (.A1(_1854_),
    .A2(_1712_),
    .B1(_1713_),
    .B2(_1580_),
    .Y(_2085_));
 sky130_fd_sc_hd__a22oi_2 _5224_ (.A1(_1529_),
    .A2(_1712_),
    .B1(_1713_),
    .B2(_1594_),
    .Y(_2086_));
 sky130_fd_sc_hd__buf_4 _5225_ (.A(_1372_),
    .X(_2087_));
 sky130_fd_sc_hd__mux4_2 _5226_ (.A0(_2082_),
    .A1(_2084_),
    .A2(_2085_),
    .A3(_2086_),
    .S0(_1706_),
    .S1(_2087_),
    .X(_2088_));
 sky130_fd_sc_hd__or2_1 _5227_ (.A(_1757_),
    .B(_1761_),
    .X(_2089_));
 sky130_fd_sc_hd__or2_1 _5228_ (.A(_1778_),
    .B(_1777_),
    .X(_2090_));
 sky130_fd_sc_hd__nor2_1 _5229_ (.A(_1766_),
    .B(_2090_),
    .Y(_2091_));
 sky130_fd_sc_hd__a22o_1 _5230_ (.A1(_1785_),
    .A2(_1786_),
    .B1(_1766_),
    .B2(_2090_),
    .X(_2092_));
 sky130_fd_sc_hd__inv_2 _5231_ (.A(_2090_),
    .Y(_2093_));
 sky130_fd_sc_hd__clkinv_2 _5232_ (.A(_1788_),
    .Y(_2094_));
 sky130_fd_sc_hd__clkinv_2 _5233_ (.A(\core_1.decode.oc_alu_mode[9] ),
    .Y(_2095_));
 sky130_fd_sc_hd__nor2_1 _5234_ (.A(_2095_),
    .B(_1777_),
    .Y(_2096_));
 sky130_fd_sc_hd__a221o_1 _5235_ (.A1(\core_1.decode.oc_alu_mode[7] ),
    .A2(_1693_),
    .B1(_1741_),
    .B2(_2094_),
    .C1(_2096_),
    .X(_2097_));
 sky130_fd_sc_hd__a221o_1 _5236_ (.A1(\core_1.decode.oc_alu_mode[2] ),
    .A2(_1778_),
    .B1(_2093_),
    .B2(\core_1.decode.oc_alu_mode[6] ),
    .C1(_2097_),
    .X(_2098_));
 sky130_fd_sc_hd__o21ba_1 _5237_ (.A1(_2091_),
    .A2(_2092_),
    .B1_N(_2098_),
    .X(_2099_));
 sky130_fd_sc_hd__o2bb2a_1 _5238_ (.A1_N(_1665_),
    .A2_N(_1712_),
    .B1(_1709_),
    .B2(_1650_),
    .X(_2100_));
 sky130_fd_sc_hd__o2bb2a_1 _5239_ (.A1_N(_1557_),
    .A2_N(_1712_),
    .B1(_1709_),
    .B2(_1885_),
    .X(_2101_));
 sky130_fd_sc_hd__mux2_1 _5240_ (.A0(_2100_),
    .A1(_2101_),
    .S(_1705_),
    .X(_2102_));
 sky130_fd_sc_hd__o2bb2a_1 _5241_ (.A1_N(_1723_),
    .A2_N(_1712_),
    .B1(_1709_),
    .B2(_1727_),
    .X(_2103_));
 sky130_fd_sc_hd__a2111o_1 _5242_ (.A1(_1693_),
    .A2(_1731_),
    .B1(_1703_),
    .C1(_1777_),
    .D1(_1705_),
    .X(_2104_));
 sky130_fd_sc_hd__o211a_1 _5243_ (.A1(_1691_),
    .A2(_2103_),
    .B1(_2104_),
    .C1(_1384_),
    .X(_2105_));
 sky130_fd_sc_hd__nor2_2 _5244_ (.A(_1361_),
    .B(_1735_),
    .Y(_2106_));
 sky130_fd_sc_hd__nand2_2 _5245_ (.A(_1369_),
    .B(_2106_),
    .Y(_2107_));
 sky130_fd_sc_hd__a211o_1 _5246_ (.A1(_1372_),
    .A2(_2102_),
    .B1(_2105_),
    .C1(_2107_),
    .X(_2108_));
 sky130_fd_sc_hd__o311a_1 _5247_ (.A1(_1758_),
    .A2(_1749_),
    .A3(_2089_),
    .B1(_2099_),
    .C1(_2108_),
    .X(_2109_));
 sky130_fd_sc_hd__o31a_2 _5248_ (.A1(_1369_),
    .A2(_1736_),
    .A3(_2088_),
    .B1(_2109_),
    .X(_2110_));
 sky130_fd_sc_hd__inv_2 _5249_ (.A(\core_1.execute.alu_mul_div.mul_res[0] ),
    .Y(_2111_));
 sky130_fd_sc_hd__a21o_1 _5250_ (.A1(_1688_),
    .A2(_2111_),
    .B1(\core_1.execute.alu_mul_div.i_div ),
    .X(_2112_));
 sky130_fd_sc_hd__a21oi_2 _5251_ (.A1(_2081_),
    .A2(_2110_),
    .B1(_2112_),
    .Y(_2113_));
 sky130_fd_sc_hd__o22a_2 _5252_ (.A1(_1686_),
    .A2(\core_1.execute.alu_mul_div.div_cur[0] ),
    .B1(_2080_),
    .B2(_2113_),
    .X(_2114_));
 sky130_fd_sc_hd__nor2_2 _5253_ (.A(\core_1.dec_sreg_jal_over ),
    .B(\core_1.dec_sreg_load ),
    .Y(_2115_));
 sky130_fd_sc_hd__buf_4 _5254_ (.A(_2115_),
    .X(_2116_));
 sky130_fd_sc_hd__buf_4 _5255_ (.A(_2116_),
    .X(_2117_));
 sky130_fd_sc_hd__mux2_1 _5256_ (.A0(_2079_),
    .A1(_2114_),
    .S(_2117_),
    .X(_2118_));
 sky130_fd_sc_hd__mux2_1 _5257_ (.A0(_2118_),
    .A1(net194),
    .S(_1147_),
    .X(_2119_));
 sky130_fd_sc_hd__buf_4 _5258_ (.A(_2008_),
    .X(_2120_));
 sky130_fd_sc_hd__mux2_1 _5259_ (.A0(\core_1.ew_data[0] ),
    .A1(_2119_),
    .S(_2120_),
    .X(_2121_));
 sky130_fd_sc_hd__clkbuf_1 _5260_ (.A(_2121_),
    .X(_0229_));
 sky130_fd_sc_hd__a21o_2 _5261_ (.A1(_1052_),
    .A2(_1056_),
    .B1(\core_1.dec_sreg_jal_over ),
    .X(_2122_));
 sky130_fd_sc_hd__and2_1 _5262_ (.A(net79),
    .B(_2122_),
    .X(_2123_));
 sky130_fd_sc_hd__and3_1 _5263_ (.A(\core_1.execute.alu_flag_reg.o_d[1] ),
    .B(_1056_),
    .C(_2066_),
    .X(_2124_));
 sky130_fd_sc_hd__and3_1 _5264_ (.A(\core_1.execute.sreg_irq_flags.o_d[1] ),
    .B(_1160_),
    .C(_2059_),
    .X(_2125_));
 sky130_fd_sc_hd__a221o_1 _5265_ (.A1(\core_1.execute.pc_high_buff_out[1] ),
    .A2(_2065_),
    .B1(_2071_),
    .B2(net8),
    .C1(_2125_),
    .X(_2126_));
 sky130_fd_sc_hd__and2_1 _5266_ (.A(_1052_),
    .B(_2060_),
    .X(_2127_));
 sky130_fd_sc_hd__a22o_1 _5267_ (.A1(\core_1.execute.sreg_irq_pc.o_d[1] ),
    .A2(_2057_),
    .B1(_2127_),
    .B2(\core_1.execute.trap_flag ),
    .X(_2128_));
 sky130_fd_sc_hd__and2_4 _5268_ (.A(_1056_),
    .B(_2064_),
    .X(_2129_));
 sky130_fd_sc_hd__and3_1 _5269_ (.A(\core_1.execute.sreg_scratch.o_d[1] ),
    .B(_2059_),
    .C(_2060_),
    .X(_2130_));
 sky130_fd_sc_hd__a221o_1 _5270_ (.A1(\core_1.execute.sreg_data_page ),
    .A2(_1161_),
    .B1(_2129_),
    .B2(\core_1.execute.pc_high_out[1] ),
    .C1(_2130_),
    .X(_2131_));
 sky130_fd_sc_hd__o41a_1 _5271_ (.A1(_2124_),
    .A2(_2126_),
    .A3(_2128_),
    .A4(_2131_),
    .B1(_2054_),
    .X(_2132_));
 sky130_fd_sc_hd__o21a_1 _5272_ (.A1(_2123_),
    .A2(_2132_),
    .B1(_1798_),
    .X(_2133_));
 sky130_fd_sc_hd__o2111ai_4 _5273_ (.A1(_1802_),
    .A2(_2133_),
    .B1(_2053_),
    .C1(\core_1.dec_sreg_jal_over ),
    .D1(_2077_),
    .Y(_2134_));
 sky130_fd_sc_hd__buf_4 _5274_ (.A(_2054_),
    .X(_2135_));
 sky130_fd_sc_hd__o21bai_1 _5275_ (.A1(_1802_),
    .A2(_2133_),
    .B1_N(_2116_),
    .Y(_2136_));
 sky130_fd_sc_hd__o21ai_1 _5276_ (.A1(_2135_),
    .A2(_2078_),
    .B1(_2136_),
    .Y(_2137_));
 sky130_fd_sc_hd__a22o_1 _5277_ (.A1(_1797_),
    .A2(_2117_),
    .B1(_2134_),
    .B2(_2137_),
    .X(_2138_));
 sky130_fd_sc_hd__mux2_1 _5278_ (.A0(_2138_),
    .A1(net201),
    .S(_1147_),
    .X(_2139_));
 sky130_fd_sc_hd__mux2_1 _5279_ (.A0(\core_1.ew_data[1] ),
    .A1(_2139_),
    .S(_2120_),
    .X(_2140_));
 sky130_fd_sc_hd__clkbuf_1 _5280_ (.A(_2140_),
    .X(_0230_));
 sky130_fd_sc_hd__a21o_1 _5281_ (.A1(net80),
    .A2(_2122_),
    .B1(\core_1.dec_sreg_irt ),
    .X(_2141_));
 sky130_fd_sc_hd__and3_1 _5282_ (.A(\core_1.execute.pc_high_buff_out[2] ),
    .B(_1160_),
    .C(_2064_),
    .X(_2142_));
 sky130_fd_sc_hd__a221o_1 _5283_ (.A1(\core_1.execute.sreg_irq_pc.o_d[2] ),
    .A2(_2057_),
    .B1(_2127_),
    .B2(_0671_),
    .C1(_2142_),
    .X(_2143_));
 sky130_fd_sc_hd__a22o_1 _5284_ (.A1(\core_1.execute.pc_high_out[2] ),
    .A2(_2129_),
    .B1(_2071_),
    .B2(net9),
    .X(_2144_));
 sky130_fd_sc_hd__and2_1 _5285_ (.A(_1056_),
    .B(_2066_),
    .X(_2145_));
 sky130_fd_sc_hd__and2_2 _5286_ (.A(_2066_),
    .B(_2060_),
    .X(_2146_));
 sky130_fd_sc_hd__a32o_1 _5287_ (.A1(\core_1.execute.sreg_irq_flags.o_d[2] ),
    .A2(_1160_),
    .A3(_2066_),
    .B1(_1161_),
    .B2(\core_1.execute.irq_en ),
    .X(_2147_));
 sky130_fd_sc_hd__a221o_1 _5288_ (.A1(\core_1.execute.alu_flag_reg.o_d[2] ),
    .A2(_2145_),
    .B1(_2146_),
    .B2(\core_1.execute.sreg_scratch.o_d[2] ),
    .C1(_2147_),
    .X(_2148_));
 sky130_fd_sc_hd__o31a_1 _5289_ (.A1(_2143_),
    .A2(_2144_),
    .A3(_2148_),
    .B1(_2054_),
    .X(_2149_));
 sky130_fd_sc_hd__o22a_1 _5290_ (.A1(\core_1.execute.sreg_irq_pc.o_d[2] ),
    .A2(_1798_),
    .B1(_2141_),
    .B2(_2149_),
    .X(_2150_));
 sky130_fd_sc_hd__xnor2_1 _5291_ (.A(_2134_),
    .B(_2150_),
    .Y(_2151_));
 sky130_fd_sc_hd__a21bo_1 _5292_ (.A1(\core_1.execute.alu_mul_div.div_res[2] ),
    .A2(_1685_),
    .B1_N(_0732_),
    .X(_2152_));
 sky130_fd_sc_hd__mux2_1 _5293_ (.A0(_2082_),
    .A1(_2101_),
    .S(_1691_),
    .X(_2153_));
 sky130_fd_sc_hd__mux2_1 _5294_ (.A0(_2100_),
    .A1(_2103_),
    .S(_1691_),
    .X(_2154_));
 sky130_fd_sc_hd__mux2_1 _5295_ (.A0(_2153_),
    .A1(_2154_),
    .S(_1384_),
    .X(_2155_));
 sky130_fd_sc_hd__nand2_1 _5296_ (.A(_1369_),
    .B(_2155_),
    .Y(_2156_));
 sky130_fd_sc_hd__mux2_1 _5297_ (.A0(_2084_),
    .A1(_2085_),
    .S(_1706_),
    .X(_2157_));
 sky130_fd_sc_hd__or2_1 _5298_ (.A(_1706_),
    .B(_2086_),
    .X(_2158_));
 sky130_fd_sc_hd__mux2_1 _5299_ (.A0(_2157_),
    .A1(_2158_),
    .S(_2087_),
    .X(_2159_));
 sky130_fd_sc_hd__a21oi_1 _5300_ (.A1(_1689_),
    .A2(_2159_),
    .B1(_1736_),
    .Y(_2160_));
 sky130_fd_sc_hd__o21a_1 _5301_ (.A1(_0988_),
    .A2(_1741_),
    .B1(_1748_),
    .X(_2161_));
 sky130_fd_sc_hd__o21a_1 _5302_ (.A1(_0988_),
    .A2(_1751_),
    .B1(_1748_),
    .X(_2162_));
 sky130_fd_sc_hd__o21a_1 _5303_ (.A1(_0988_),
    .A2(_1974_),
    .B1(_1748_),
    .X(_2163_));
 sky130_fd_sc_hd__mux2_1 _5304_ (.A0(_2162_),
    .A1(_2163_),
    .S(_1419_),
    .X(_2164_));
 sky130_fd_sc_hd__clkbuf_4 _5305_ (.A(_1982_),
    .X(_2165_));
 sky130_fd_sc_hd__a22o_1 _5306_ (.A1(_1694_),
    .A2(_2161_),
    .B1(_2164_),
    .B2(_2165_),
    .X(_2166_));
 sky130_fd_sc_hd__a21o_1 _5307_ (.A1(_1782_),
    .A2(_1779_),
    .B1(_1775_),
    .X(_2167_));
 sky130_fd_sc_hd__a2bb2o_1 _5308_ (.A1_N(_1785_),
    .A2_N(_2167_),
    .B1(_1899_),
    .B2(\core_1.decode.oc_alu_mode[11] ),
    .X(_2168_));
 sky130_fd_sc_hd__inv_2 _5309_ (.A(_1945_),
    .Y(_2169_));
 sky130_fd_sc_hd__nor2_1 _5310_ (.A(_2169_),
    .B(_1946_),
    .Y(_2170_));
 sky130_fd_sc_hd__o21a_1 _5311_ (.A1(_0931_),
    .A2(_2168_),
    .B1(_2170_),
    .X(_2171_));
 sky130_fd_sc_hd__buf_4 _5312_ (.A(_1786_),
    .X(_2172_));
 sky130_fd_sc_hd__o2bb2a_1 _5313_ (.A1_N(_0966_),
    .A2_N(_2167_),
    .B1(_1899_),
    .B2(_2172_),
    .X(_2173_));
 sky130_fd_sc_hd__nor2_1 _5314_ (.A(_2170_),
    .B(_2173_),
    .Y(_2174_));
 sky130_fd_sc_hd__nor2_1 _5315_ (.A(_1727_),
    .B(_1788_),
    .Y(_2175_));
 sky130_fd_sc_hd__a221o_1 _5316_ (.A1(_0937_),
    .A2(_2087_),
    .B1(_1945_),
    .B2(_0960_),
    .C1(_2175_),
    .X(_2176_));
 sky130_fd_sc_hd__a2111o_1 _5317_ (.A1(_1000_),
    .A2(_1946_),
    .B1(_2171_),
    .C1(_2174_),
    .D1(_2176_),
    .X(_2177_));
 sky130_fd_sc_hd__a31o_1 _5318_ (.A1(_1762_),
    .A2(_1765_),
    .A3(_2166_),
    .B1(_2177_),
    .X(_2178_));
 sky130_fd_sc_hd__a21oi_1 _5319_ (.A1(_2156_),
    .A2(_2160_),
    .B1(_2178_),
    .Y(_2179_));
 sky130_fd_sc_hd__nor2_1 _5320_ (.A(_1688_),
    .B(_2179_),
    .Y(_2180_));
 sky130_fd_sc_hd__a211o_1 _5321_ (.A1(_1688_),
    .A2(\core_1.execute.alu_mul_div.mul_res[2] ),
    .B1(_2180_),
    .C1(_0992_),
    .X(_2181_));
 sky130_fd_sc_hd__a22o_2 _5322_ (.A1(\core_1.execute.alu_mul_div.div_cur[2] ),
    .A2(\core_1.execute.alu_mul_div.i_mod ),
    .B1(_2152_),
    .B2(_2181_),
    .X(_2182_));
 sky130_fd_sc_hd__mux2_1 _5323_ (.A0(_2151_),
    .A1(_2182_),
    .S(_2117_),
    .X(_2183_));
 sky130_fd_sc_hd__mux2_1 _5324_ (.A0(_2183_),
    .A1(net202),
    .S(_1147_),
    .X(_2184_));
 sky130_fd_sc_hd__mux2_1 _5325_ (.A0(\core_1.ew_data[2] ),
    .A1(_2184_),
    .S(_2120_),
    .X(_2185_));
 sky130_fd_sc_hd__clkbuf_1 _5326_ (.A(_2185_),
    .X(_0231_));
 sky130_fd_sc_hd__or2b_1 _5327_ (.A(_2134_),
    .B_N(_2150_),
    .X(_2186_));
 sky130_fd_sc_hd__a22o_1 _5328_ (.A1(\core_1.execute.sreg_long_ptr_en ),
    .A2(_1161_),
    .B1(_2071_),
    .B2(net10),
    .X(_2187_));
 sky130_fd_sc_hd__a22o_1 _5329_ (.A1(\core_1.execute.sreg_scratch.o_d[3] ),
    .A2(_2146_),
    .B1(_2065_),
    .B2(\core_1.execute.pc_high_buff_out[3] ),
    .X(_2188_));
 sky130_fd_sc_hd__a32o_1 _5330_ (.A1(\core_1.execute.sreg_irq_flags.o_d[3] ),
    .A2(_1160_),
    .A3(_2066_),
    .B1(_2057_),
    .B2(\core_1.execute.sreg_irq_pc.o_d[3] ),
    .X(_2189_));
 sky130_fd_sc_hd__a22o_1 _5331_ (.A1(\core_1.execute.alu_flag_reg.o_d[3] ),
    .A2(_2145_),
    .B1(_2129_),
    .B2(\core_1.execute.pc_high_out[3] ),
    .X(_2190_));
 sky130_fd_sc_hd__or4_1 _5332_ (.A(_2187_),
    .B(_2188_),
    .C(_2189_),
    .D(_2190_),
    .X(_2191_));
 sky130_fd_sc_hd__a22o_1 _5333_ (.A1(net81),
    .A2(_2122_),
    .B1(_2191_),
    .B2(_2054_),
    .X(_2192_));
 sky130_fd_sc_hd__mux2_1 _5334_ (.A0(\core_1.execute.sreg_irq_pc.o_d[3] ),
    .A1(_2192_),
    .S(_1798_),
    .X(_2193_));
 sky130_fd_sc_hd__xnor2_1 _5335_ (.A(_2186_),
    .B(_2193_),
    .Y(_2194_));
 sky130_fd_sc_hd__a21bo_1 _5336_ (.A1(\core_1.execute.alu_mul_div.div_res[3] ),
    .A2(_1686_),
    .B1_N(_0732_),
    .X(_2195_));
 sky130_fd_sc_hd__nand2_1 _5337_ (.A(_1945_),
    .B(_1947_),
    .Y(_2196_));
 sky130_fd_sc_hd__or3_1 _5338_ (.A(_1785_),
    .B(_1903_),
    .C(_2196_),
    .X(_2197_));
 sky130_fd_sc_hd__a221o_1 _5339_ (.A1(_0937_),
    .A2(_1689_),
    .B1(_1901_),
    .B2(_1000_),
    .C1(_0960_),
    .X(_2198_));
 sky130_fd_sc_hd__nand2_1 _5340_ (.A(_1902_),
    .B(_2198_),
    .Y(_2199_));
 sky130_fd_sc_hd__a21o_1 _5341_ (.A1(_1898_),
    .A2(_1899_),
    .B1(_1900_),
    .X(_2200_));
 sky130_fd_sc_hd__a221o_1 _5342_ (.A1(_0981_),
    .A2(_2200_),
    .B1(_2196_),
    .B2(_0966_),
    .C1(\core_1.decode.oc_alu_mode[6] ),
    .X(_2201_));
 sky130_fd_sc_hd__nand2_1 _5343_ (.A(_1903_),
    .B(_2201_),
    .Y(_2202_));
 sky130_fd_sc_hd__o221a_1 _5344_ (.A1(_1643_),
    .A2(_1788_),
    .B1(_1904_),
    .B2(_2172_),
    .C1(_2202_),
    .X(_2203_));
 sky130_fd_sc_hd__mux2_1 _5345_ (.A0(_1715_),
    .A1(_1720_),
    .S(_1691_),
    .X(_2204_));
 sky130_fd_sc_hd__a31o_1 _5346_ (.A1(_1691_),
    .A2(_1708_),
    .A3(_1725_),
    .B1(_2087_),
    .X(_2205_));
 sky130_fd_sc_hd__a21oi_1 _5347_ (.A1(_1706_),
    .A2(_1718_),
    .B1(_2205_),
    .Y(_2206_));
 sky130_fd_sc_hd__a211o_1 _5348_ (.A1(_2087_),
    .A2(_2204_),
    .B1(_2206_),
    .C1(_2107_),
    .X(_2207_));
 sky130_fd_sc_hd__and4_1 _5349_ (.A(_2197_),
    .B(_2199_),
    .C(_2203_),
    .D(_2207_),
    .X(_2208_));
 sky130_fd_sc_hd__mux2_1 _5350_ (.A0(_1975_),
    .A1(_1978_),
    .S(_1419_),
    .X(_2209_));
 sky130_fd_sc_hd__mux2_1 _5351_ (.A0(_1753_),
    .A1(_2209_),
    .S(_2165_),
    .X(_2210_));
 sky130_fd_sc_hd__or3_1 _5352_ (.A(_2089_),
    .B(_1983_),
    .C(_2210_),
    .X(_2211_));
 sky130_fd_sc_hd__mux2_1 _5353_ (.A0(_1710_),
    .A1(_1714_),
    .S(_1691_),
    .X(_2212_));
 sky130_fd_sc_hd__nor2_1 _5354_ (.A(_1372_),
    .B(_2212_),
    .Y(_2213_));
 sky130_fd_sc_hd__a31o_1 _5355_ (.A1(_1372_),
    .A2(_1704_),
    .A3(_1730_),
    .B1(_2213_),
    .X(_2214_));
 sky130_fd_sc_hd__or3b_1 _5356_ (.A(_1369_),
    .B(_1736_),
    .C_N(_2214_),
    .X(_2215_));
 sky130_fd_sc_hd__and3_2 _5357_ (.A(_2208_),
    .B(_2211_),
    .C(_2215_),
    .X(_2216_));
 sky130_fd_sc_hd__nor2_1 _5358_ (.A(_1688_),
    .B(_2216_),
    .Y(_2217_));
 sky130_fd_sc_hd__a211o_1 _5359_ (.A1(_0959_),
    .A2(\core_1.execute.alu_mul_div.mul_res[3] ),
    .B1(_2217_),
    .C1(_0992_),
    .X(_2218_));
 sky130_fd_sc_hd__a22o_2 _5360_ (.A1(\core_1.execute.alu_mul_div.div_cur[3] ),
    .A2(_0964_),
    .B1(_2195_),
    .B2(_2218_),
    .X(_2219_));
 sky130_fd_sc_hd__mux2_1 _5361_ (.A0(_2194_),
    .A1(_2219_),
    .S(_2117_),
    .X(_2220_));
 sky130_fd_sc_hd__mux2_1 _5362_ (.A0(_2220_),
    .A1(net203),
    .S(_1147_),
    .X(_2221_));
 sky130_fd_sc_hd__mux2_1 _5363_ (.A0(\core_1.ew_data[3] ),
    .A1(_2221_),
    .S(_2120_),
    .X(_2222_));
 sky130_fd_sc_hd__clkbuf_1 _5364_ (.A(_2222_),
    .X(_0232_));
 sky130_fd_sc_hd__a21boi_1 _5365_ (.A1(\core_1.execute.alu_mul_div.div_res[4] ),
    .A2(_1685_),
    .B1_N(_0732_),
    .Y(_2223_));
 sky130_fd_sc_hd__and2_1 _5366_ (.A(_1748_),
    .B(_1977_),
    .X(_2224_));
 sky130_fd_sc_hd__mux2_1 _5367_ (.A0(_1979_),
    .A1(_2224_),
    .S(_1693_),
    .X(_2225_));
 sky130_fd_sc_hd__mux2_1 _5368_ (.A0(_2225_),
    .A1(_2164_),
    .S(_1740_),
    .X(_2226_));
 sky130_fd_sc_hd__a32o_1 _5369_ (.A1(_2087_),
    .A2(_1730_),
    .A3(_2161_),
    .B1(_1764_),
    .B2(_2226_),
    .X(_2227_));
 sky130_fd_sc_hd__mux2_1 _5370_ (.A0(_2086_),
    .A1(_2085_),
    .S(_1691_),
    .X(_2228_));
 sky130_fd_sc_hd__nor2_2 _5371_ (.A(_2087_),
    .B(_2228_),
    .Y(_2229_));
 sky130_fd_sc_hd__mux2_1 _5372_ (.A0(_2082_),
    .A1(_2084_),
    .S(_1706_),
    .X(_2230_));
 sky130_fd_sc_hd__a22oi_1 _5373_ (.A1(_1722_),
    .A2(_2230_),
    .B1(_2102_),
    .B2(_1734_),
    .Y(_2231_));
 sky130_fd_sc_hd__o211a_1 _5374_ (.A1(_1369_),
    .A2(_2229_),
    .B1(_2231_),
    .C1(_2106_),
    .X(_2232_));
 sky130_fd_sc_hd__and2_1 _5375_ (.A(_1905_),
    .B(_1948_),
    .X(_2233_));
 sky130_fd_sc_hd__nor2_1 _5376_ (.A(_1785_),
    .B(_2233_),
    .Y(_2234_));
 sky130_fd_sc_hd__o21a_1 _5377_ (.A1(_1905_),
    .A2(_1948_),
    .B1(_2234_),
    .X(_2235_));
 sky130_fd_sc_hd__mux2_1 _5378_ (.A0(_1905_),
    .A1(_1909_),
    .S(_1904_),
    .X(_2236_));
 sky130_fd_sc_hd__nor2_1 _5379_ (.A(_2172_),
    .B(_2236_),
    .Y(_2237_));
 sky130_fd_sc_hd__a21oi_1 _5380_ (.A1(_1364_),
    .A2(_1650_),
    .B1(_2095_),
    .Y(_2238_));
 sky130_fd_sc_hd__a221o_1 _5381_ (.A1(\core_1.decode.oc_alu_mode[7] ),
    .A2(_1361_),
    .B1(_1724_),
    .B2(_2094_),
    .C1(_2238_),
    .X(_2239_));
 sky130_fd_sc_hd__a221o_1 _5382_ (.A1(_1000_),
    .A2(_1953_),
    .B1(_1905_),
    .B2(_0931_),
    .C1(_2239_),
    .X(_2240_));
 sky130_fd_sc_hd__or3_1 _5383_ (.A(_2235_),
    .B(_2237_),
    .C(_2240_),
    .X(_2241_));
 sky130_fd_sc_hd__a211o_2 _5384_ (.A1(_1762_),
    .A2(_2227_),
    .B1(_2232_),
    .C1(_2241_),
    .X(_2242_));
 sky130_fd_sc_hd__a21o_1 _5385_ (.A1(_0958_),
    .A2(\core_1.execute.alu_mul_div.mul_res[4] ),
    .B1(\core_1.execute.alu_mul_div.i_div ),
    .X(_2243_));
 sky130_fd_sc_hd__a21oi_2 _5386_ (.A1(_2081_),
    .A2(_2242_),
    .B1(_2243_),
    .Y(_2244_));
 sky130_fd_sc_hd__o22a_2 _5387_ (.A1(_1359_),
    .A2(_1685_),
    .B1(_2223_),
    .B2(_2244_),
    .X(_2245_));
 sky130_fd_sc_hd__inv_2 _5388_ (.A(_2245_),
    .Y(_2246_));
 sky130_fd_sc_hd__and2_4 _5389_ (.A(_2066_),
    .B(_2056_),
    .X(_2247_));
 sky130_fd_sc_hd__a221o_1 _5390_ (.A1(\core_1.execute.sreg_irq_pc.o_d[4] ),
    .A2(_2057_),
    .B1(_2065_),
    .B2(\core_1.execute.pc_high_buff_out[4] ),
    .C1(_2247_),
    .X(_2248_));
 sky130_fd_sc_hd__a22o_1 _5391_ (.A1(\core_1.execute.sreg_scratch.o_d[4] ),
    .A2(_2146_),
    .B1(_2071_),
    .B2(net11),
    .X(_2249_));
 sky130_fd_sc_hd__and3_1 _5392_ (.A(\core_1.execute.sreg_irq_flags.o_d[4] ),
    .B(_1160_),
    .C(_2066_),
    .X(_2250_));
 sky130_fd_sc_hd__a221o_1 _5393_ (.A1(\core_1.execute.sreg_priv_control.o_d[4] ),
    .A2(_1161_),
    .B1(_2129_),
    .B2(\core_1.execute.pc_high_out[4] ),
    .C1(_2250_),
    .X(_2251_));
 sky130_fd_sc_hd__a2111o_1 _5394_ (.A1(\core_1.execute.alu_flag_reg.o_d[4] ),
    .A2(_2145_),
    .B1(_2248_),
    .C1(_2249_),
    .D1(_2251_),
    .X(_2252_));
 sky130_fd_sc_hd__a22o_1 _5395_ (.A1(net82),
    .A2(_2122_),
    .B1(_2252_),
    .B2(_2054_),
    .X(_2253_));
 sky130_fd_sc_hd__mux2_1 _5396_ (.A0(\core_1.execute.sreg_irq_pc.o_d[4] ),
    .A1(_2253_),
    .S(_1798_),
    .X(_2254_));
 sky130_fd_sc_hd__nand3b_1 _5397_ (.A_N(_2186_),
    .B(_2193_),
    .C(_2254_),
    .Y(_2255_));
 sky130_fd_sc_hd__and2b_1 _5398_ (.A_N(_2186_),
    .B(_2193_),
    .X(_2256_));
 sky130_fd_sc_hd__o21ba_1 _5399_ (.A1(_2256_),
    .A2(_2254_),
    .B1_N(_2115_),
    .X(_2257_));
 sky130_fd_sc_hd__a22oi_1 _5400_ (.A1(_2116_),
    .A2(_2246_),
    .B1(_2255_),
    .B2(_2257_),
    .Y(_2258_));
 sky130_fd_sc_hd__mux2_1 _5401_ (.A0(_2258_),
    .A1(_0633_),
    .S(\core_1.dec_mem_access ),
    .X(_2259_));
 sky130_fd_sc_hd__inv_2 _5402_ (.A(_2259_),
    .Y(_2260_));
 sky130_fd_sc_hd__mux2_1 _5403_ (.A0(\core_1.ew_data[4] ),
    .A1(_2260_),
    .S(_2120_),
    .X(_2261_));
 sky130_fd_sc_hd__clkbuf_1 _5404_ (.A(_2261_),
    .X(_0233_));
 sky130_fd_sc_hd__a22o_1 _5405_ (.A1(\core_1.execute.pc_high_out[5] ),
    .A2(_2129_),
    .B1(_2071_),
    .B2(net12),
    .X(_2262_));
 sky130_fd_sc_hd__a221o_1 _5406_ (.A1(\core_1.execute.sreg_irq_pc.o_d[5] ),
    .A2(_2057_),
    .B1(_2146_),
    .B2(\core_1.execute.sreg_scratch.o_d[5] ),
    .C1(_2262_),
    .X(_2263_));
 sky130_fd_sc_hd__a221o_1 _5407_ (.A1(\core_1.execute.sreg_priv_control.o_d[5] ),
    .A2(_1161_),
    .B1(_2065_),
    .B2(\core_1.execute.pc_high_buff_out[5] ),
    .C1(_2263_),
    .X(_2264_));
 sky130_fd_sc_hd__a22o_1 _5408_ (.A1(net83),
    .A2(_2122_),
    .B1(_2264_),
    .B2(_2054_),
    .X(_2265_));
 sky130_fd_sc_hd__and2_1 _5409_ (.A(\core_1.execute.sreg_irq_pc.o_d[5] ),
    .B(\core_1.dec_sreg_irt ),
    .X(_2266_));
 sky130_fd_sc_hd__a21oi_1 _5410_ (.A1(_1798_),
    .A2(_2265_),
    .B1(_2266_),
    .Y(_2267_));
 sky130_fd_sc_hd__nand2_1 _5411_ (.A(_2255_),
    .B(_2267_),
    .Y(_2268_));
 sky130_fd_sc_hd__or2_1 _5412_ (.A(_2255_),
    .B(_2267_),
    .X(_2269_));
 sky130_fd_sc_hd__and2_1 _5413_ (.A(_2268_),
    .B(_2269_),
    .X(_2270_));
 sky130_fd_sc_hd__a21bo_1 _5414_ (.A1(\core_1.execute.alu_mul_div.div_res[5] ),
    .A2(_1686_),
    .B1_N(_1407_),
    .X(_2271_));
 sky130_fd_sc_hd__mux2_1 _5415_ (.A0(_2163_),
    .A1(_2224_),
    .S(_1418_),
    .X(_2272_));
 sky130_fd_sc_hd__mux2_1 _5416_ (.A0(_1967_),
    .A1(_1979_),
    .S(_1692_),
    .X(_2273_));
 sky130_fd_sc_hd__mux2_1 _5417_ (.A0(_2272_),
    .A1(_2273_),
    .S(_1982_),
    .X(_2274_));
 sky130_fd_sc_hd__mux2_2 _5418_ (.A0(_1754_),
    .A1(_2274_),
    .S(_1764_),
    .X(_2275_));
 sky130_fd_sc_hd__or2_1 _5419_ (.A(_1953_),
    .B(_2233_),
    .X(_2276_));
 sky130_fd_sc_hd__o21ai_1 _5420_ (.A1(_1894_),
    .A2(_2276_),
    .B1(_0966_),
    .Y(_2277_));
 sky130_fd_sc_hd__a21oi_1 _5421_ (.A1(_1894_),
    .A2(_2276_),
    .B1(_2277_),
    .Y(_2278_));
 sky130_fd_sc_hd__a21o_1 _5422_ (.A1(_1904_),
    .A2(_1906_),
    .B1(_1905_),
    .X(_2279_));
 sky130_fd_sc_hd__a21oi_1 _5423_ (.A1(_1897_),
    .A2(_2279_),
    .B1(_2172_),
    .Y(_2280_));
 sky130_fd_sc_hd__o21a_1 _5424_ (.A1(_1897_),
    .A2(_2279_),
    .B1(_2280_),
    .X(_2281_));
 sky130_fd_sc_hd__a21oi_1 _5425_ (.A1(_2087_),
    .A2(_1716_),
    .B1(_1689_),
    .Y(_2282_));
 sky130_fd_sc_hd__nor2_1 _5426_ (.A(_1372_),
    .B(_1711_),
    .Y(_2283_));
 sky130_fd_sc_hd__nand2_1 _5427_ (.A(_1721_),
    .B(_1734_),
    .Y(_2284_));
 sky130_fd_sc_hd__o211a_1 _5428_ (.A1(_2282_),
    .A2(_2283_),
    .B1(_2284_),
    .C1(_2106_),
    .X(_2285_));
 sky130_fd_sc_hd__a22o_1 _5429_ (.A1(_0937_),
    .A2(_1696_),
    .B1(_1665_),
    .B2(_2094_),
    .X(_2286_));
 sky130_fd_sc_hd__a221o_1 _5430_ (.A1(_0960_),
    .A2(_1954_),
    .B1(_1894_),
    .B2(_0931_),
    .C1(_2286_),
    .X(_2287_));
 sky130_fd_sc_hd__a2111o_1 _5431_ (.A1(_1000_),
    .A2(_1952_),
    .B1(_2281_),
    .C1(_2285_),
    .D1(_2287_),
    .X(_2288_));
 sky130_fd_sc_hd__a211o_1 _5432_ (.A1(_1762_),
    .A2(_2275_),
    .B1(_2278_),
    .C1(_2288_),
    .X(_2289_));
 sky130_fd_sc_hd__a21o_1 _5433_ (.A1(_0958_),
    .A2(\core_1.execute.alu_mul_div.mul_res[5] ),
    .B1(\core_1.execute.alu_mul_div.i_div ),
    .X(_2290_));
 sky130_fd_sc_hd__a21o_2 _5434_ (.A1(_2081_),
    .A2(_2289_),
    .B1(_2290_),
    .X(_2291_));
 sky130_fd_sc_hd__a22o_2 _5435_ (.A1(\core_1.execute.alu_mul_div.div_cur[5] ),
    .A2(_0964_),
    .B1(_2271_),
    .B2(_2291_),
    .X(_2292_));
 sky130_fd_sc_hd__mux2_1 _5436_ (.A0(_2270_),
    .A1(_2292_),
    .S(_2117_),
    .X(_2293_));
 sky130_fd_sc_hd__mux2_1 _5437_ (.A0(_2293_),
    .A1(net205),
    .S(_1146_),
    .X(_2294_));
 sky130_fd_sc_hd__mux2_1 _5438_ (.A0(\core_1.ew_data[5] ),
    .A1(_2294_),
    .S(_2120_),
    .X(_2295_));
 sky130_fd_sc_hd__clkbuf_1 _5439_ (.A(_2295_),
    .X(_0234_));
 sky130_fd_sc_hd__clkbuf_4 _5440_ (.A(_2122_),
    .X(_2296_));
 sky130_fd_sc_hd__buf_4 _5441_ (.A(_2071_),
    .X(_2297_));
 sky130_fd_sc_hd__a22o_1 _5442_ (.A1(\core_1.execute.sreg_irq_pc.o_d[6] ),
    .A2(_2057_),
    .B1(_2065_),
    .B2(\core_1.execute.pc_high_buff_out[6] ),
    .X(_2298_));
 sky130_fd_sc_hd__a221o_1 _5443_ (.A1(\core_1.execute.sreg_scratch.o_d[6] ),
    .A2(_2146_),
    .B1(_2297_),
    .B2(net13),
    .C1(_2298_),
    .X(_2299_));
 sky130_fd_sc_hd__a221o_1 _5444_ (.A1(\core_1.execute.sreg_priv_control.o_d[6] ),
    .A2(_1161_),
    .B1(_2129_),
    .B2(\core_1.execute.pc_high_out[6] ),
    .C1(_2299_),
    .X(_2300_));
 sky130_fd_sc_hd__a22o_1 _5445_ (.A1(net84),
    .A2(_2296_),
    .B1(_2300_),
    .B2(_2054_),
    .X(_2301_));
 sky130_fd_sc_hd__mux2_1 _5446_ (.A0(\core_1.execute.sreg_irq_pc.o_d[6] ),
    .A1(_2301_),
    .S(_1798_),
    .X(_2302_));
 sky130_fd_sc_hd__xnor2_1 _5447_ (.A(_2269_),
    .B(_2302_),
    .Y(_2303_));
 sky130_fd_sc_hd__a21bo_1 _5448_ (.A1(\core_1.execute.alu_mul_div.div_res[6] ),
    .A2(_1686_),
    .B1_N(_1407_),
    .X(_2304_));
 sky130_fd_sc_hd__nor2_1 _5449_ (.A(_1893_),
    .B(_1911_),
    .Y(_2305_));
 sky130_fd_sc_hd__nand2_1 _5450_ (.A(_1893_),
    .B(_1911_),
    .Y(_2306_));
 sky130_fd_sc_hd__or3b_1 _5451_ (.A(_2305_),
    .B(_2172_),
    .C_N(_2306_),
    .X(_2307_));
 sky130_fd_sc_hd__and3_1 _5452_ (.A(_1419_),
    .B(_1748_),
    .C(_1965_),
    .X(_2308_));
 sky130_fd_sc_hd__a21o_1 _5453_ (.A1(_1693_),
    .A2(_1967_),
    .B1(_2308_),
    .X(_2309_));
 sky130_fd_sc_hd__mux2_1 _5454_ (.A0(_2225_),
    .A1(_2309_),
    .S(_2165_),
    .X(_2310_));
 sky130_fd_sc_hd__mux2_2 _5455_ (.A0(_2166_),
    .A1(_2310_),
    .S(_1764_),
    .X(_2311_));
 sky130_fd_sc_hd__and2_1 _5456_ (.A(_1948_),
    .B(_1949_),
    .X(_2312_));
 sky130_fd_sc_hd__o21ai_1 _5457_ (.A1(_2312_),
    .A2(_1955_),
    .B1(_1890_),
    .Y(_2313_));
 sky130_fd_sc_hd__o31a_1 _5458_ (.A1(_1890_),
    .A2(_2312_),
    .A3(_1955_),
    .B1(_0966_),
    .X(_2314_));
 sky130_fd_sc_hd__nor2_1 _5459_ (.A(_2087_),
    .B(_2158_),
    .Y(_2315_));
 sky130_fd_sc_hd__or2_1 _5460_ (.A(_1369_),
    .B(_2315_),
    .X(_2316_));
 sky130_fd_sc_hd__a22oi_1 _5461_ (.A1(_1722_),
    .A2(_2157_),
    .B1(_2153_),
    .B2(_1734_),
    .Y(_2317_));
 sky130_fd_sc_hd__a22o_1 _5462_ (.A1(_0937_),
    .A2(_1351_),
    .B1(_1658_),
    .B2(_2094_),
    .X(_2318_));
 sky130_fd_sc_hd__a221o_1 _5463_ (.A1(_0960_),
    .A2(_1889_),
    .B1(_1890_),
    .B2(_0931_),
    .C1(_2318_),
    .X(_2319_));
 sky130_fd_sc_hd__a31o_1 _5464_ (.A1(_2106_),
    .A2(_2316_),
    .A3(_2317_),
    .B1(_2319_),
    .X(_2320_));
 sky130_fd_sc_hd__a221o_1 _5465_ (.A1(_1000_),
    .A2(_1951_),
    .B1(_2313_),
    .B2(_2314_),
    .C1(_2320_),
    .X(_2321_));
 sky130_fd_sc_hd__a21oi_1 _5466_ (.A1(_1762_),
    .A2(_2311_),
    .B1(_2321_),
    .Y(_2322_));
 sky130_fd_sc_hd__nand2_1 _5467_ (.A(_2307_),
    .B(_2322_),
    .Y(_2323_));
 sky130_fd_sc_hd__a21o_1 _5468_ (.A1(_0958_),
    .A2(\core_1.execute.alu_mul_div.mul_res[6] ),
    .B1(\core_1.execute.alu_mul_div.i_div ),
    .X(_2324_));
 sky130_fd_sc_hd__a21o_1 _5469_ (.A1(_2081_),
    .A2(_2323_),
    .B1(_2324_),
    .X(_2325_));
 sky130_fd_sc_hd__a22o_2 _5470_ (.A1(\core_1.execute.alu_mul_div.div_cur[6] ),
    .A2(_0964_),
    .B1(_2304_),
    .B2(_2325_),
    .X(_2326_));
 sky130_fd_sc_hd__mux2_1 _5471_ (.A0(_2303_),
    .A1(_2326_),
    .S(_2117_),
    .X(_2327_));
 sky130_fd_sc_hd__mux2_1 _5472_ (.A0(_2327_),
    .A1(net206),
    .S(_1146_),
    .X(_2328_));
 sky130_fd_sc_hd__mux2_1 _5473_ (.A0(\core_1.ew_data[6] ),
    .A1(_2328_),
    .S(_2120_),
    .X(_2329_));
 sky130_fd_sc_hd__clkbuf_1 _5474_ (.A(_2329_),
    .X(_0235_));
 sky130_fd_sc_hd__and2b_1 _5475_ (.A_N(_2269_),
    .B(_2302_),
    .X(_2330_));
 sky130_fd_sc_hd__buf_4 _5476_ (.A(_2146_),
    .X(_2331_));
 sky130_fd_sc_hd__buf_4 _5477_ (.A(_2057_),
    .X(_2332_));
 sky130_fd_sc_hd__a22o_1 _5478_ (.A1(\core_1.execute.pc_high_out[7] ),
    .A2(_2129_),
    .B1(_2332_),
    .B2(\core_1.execute.sreg_irq_pc.o_d[7] ),
    .X(_2333_));
 sky130_fd_sc_hd__a221o_1 _5479_ (.A1(\core_1.execute.sreg_scratch.o_d[7] ),
    .A2(_2331_),
    .B1(_2297_),
    .B2(net14),
    .C1(_2333_),
    .X(_2334_));
 sky130_fd_sc_hd__a221o_1 _5480_ (.A1(\core_1.execute.sreg_priv_control.o_d[7] ),
    .A2(_1162_),
    .B1(_2065_),
    .B2(\core_1.execute.pc_high_buff_out[7] ),
    .C1(_2334_),
    .X(_2335_));
 sky130_fd_sc_hd__a22o_1 _5481_ (.A1(net85),
    .A2(_2296_),
    .B1(_2335_),
    .B2(_2135_),
    .X(_2336_));
 sky130_fd_sc_hd__and2_1 _5482_ (.A(\core_1.execute.sreg_irq_pc.o_d[7] ),
    .B(\core_1.dec_sreg_irt ),
    .X(_2337_));
 sky130_fd_sc_hd__a21oi_1 _5483_ (.A1(_1798_),
    .A2(_2336_),
    .B1(_2337_),
    .Y(_2338_));
 sky130_fd_sc_hd__xnor2_1 _5484_ (.A(_2330_),
    .B(_2338_),
    .Y(_2339_));
 sky130_fd_sc_hd__a21bo_1 _5485_ (.A1(\core_1.execute.alu_mul_div.div_res[7] ),
    .A2(_1686_),
    .B1_N(_1407_),
    .X(_2340_));
 sky130_fd_sc_hd__nand2_1 _5486_ (.A(_1888_),
    .B(_2313_),
    .Y(_2341_));
 sky130_fd_sc_hd__a21oi_1 _5487_ (.A1(_1883_),
    .A2(_2341_),
    .B1(_1785_),
    .Y(_2342_));
 sky130_fd_sc_hd__o21a_1 _5488_ (.A1(_1883_),
    .A2(_2341_),
    .B1(_2342_),
    .X(_2343_));
 sky130_fd_sc_hd__a21o_1 _5489_ (.A1(_1893_),
    .A2(_1911_),
    .B1(_1892_),
    .X(_2344_));
 sky130_fd_sc_hd__xnor2_1 _5490_ (.A(_1887_),
    .B(_2344_),
    .Y(_2345_));
 sky130_fd_sc_hd__nor2_1 _5491_ (.A(_2172_),
    .B(_2345_),
    .Y(_2346_));
 sky130_fd_sc_hd__or4_1 _5492_ (.A(_1692_),
    .B(_1745_),
    .C(_1746_),
    .D(_1971_),
    .X(_2347_));
 sky130_fd_sc_hd__o21ai_1 _5493_ (.A1(_1419_),
    .A2(_1966_),
    .B1(_2347_),
    .Y(_2348_));
 sky130_fd_sc_hd__mux2_1 _5494_ (.A0(_2273_),
    .A1(_2348_),
    .S(_1982_),
    .X(_2349_));
 sky130_fd_sc_hd__inv_2 _5495_ (.A(_2349_),
    .Y(_2350_));
 sky130_fd_sc_hd__mux2_1 _5496_ (.A0(_2210_),
    .A1(_2350_),
    .S(_1765_),
    .X(_2351_));
 sky130_fd_sc_hd__nor2_1 _5497_ (.A(_2089_),
    .B(_2351_),
    .Y(_2352_));
 sky130_fd_sc_hd__and3_1 _5498_ (.A(_1529_),
    .B(_1708_),
    .C(_1730_),
    .X(_2353_));
 sky130_fd_sc_hd__nand2_1 _5499_ (.A(_1384_),
    .B(_2353_),
    .Y(_2354_));
 sky130_fd_sc_hd__a221o_1 _5500_ (.A1(_1734_),
    .A2(_2204_),
    .B1(_2354_),
    .B2(_1689_),
    .C1(_1736_),
    .X(_2355_));
 sky130_fd_sc_hd__a21oi_1 _5501_ (.A1(_1722_),
    .A2(_2212_),
    .B1(_2355_),
    .Y(_2356_));
 sky130_fd_sc_hd__a221o_1 _5502_ (.A1(_0937_),
    .A2(_1697_),
    .B1(_1557_),
    .B2(_2094_),
    .C1(_0960_),
    .X(_2357_));
 sky130_fd_sc_hd__a22o_1 _5503_ (.A1(_0931_),
    .A2(_1883_),
    .B1(_2357_),
    .B2(_1956_),
    .X(_2358_));
 sky130_fd_sc_hd__a211o_1 _5504_ (.A1(_1000_),
    .A2(_1881_),
    .B1(_2356_),
    .C1(_2358_),
    .X(_2359_));
 sky130_fd_sc_hd__or4_2 _5505_ (.A(_2343_),
    .B(_2346_),
    .C(_2352_),
    .D(_2359_),
    .X(_2360_));
 sky130_fd_sc_hd__a21o_1 _5506_ (.A1(_0958_),
    .A2(\core_1.execute.alu_mul_div.mul_res[7] ),
    .B1(\core_1.execute.alu_mul_div.i_div ),
    .X(_2361_));
 sky130_fd_sc_hd__a21o_1 _5507_ (.A1(_2081_),
    .A2(_2360_),
    .B1(_2361_),
    .X(_2362_));
 sky130_fd_sc_hd__a22o_2 _5508_ (.A1(\core_1.execute.alu_mul_div.div_cur[7] ),
    .A2(_0964_),
    .B1(_2340_),
    .B2(_2362_),
    .X(_2363_));
 sky130_fd_sc_hd__mux2_1 _5509_ (.A0(_2339_),
    .A1(_2363_),
    .S(_2116_),
    .X(_2364_));
 sky130_fd_sc_hd__mux2_1 _5510_ (.A0(_2364_),
    .A1(net207),
    .S(_1146_),
    .X(_2365_));
 sky130_fd_sc_hd__mux2_1 _5511_ (.A0(\core_1.ew_data[7] ),
    .A1(_2365_),
    .S(_2120_),
    .X(_2366_));
 sky130_fd_sc_hd__clkbuf_1 _5512_ (.A(_2366_),
    .X(_0236_));
 sky130_fd_sc_hd__a21bo_1 _5513_ (.A1(\core_1.execute.alu_mul_div.div_res[8] ),
    .A2(_1686_),
    .B1_N(_1407_),
    .X(_2367_));
 sky130_fd_sc_hd__or4_1 _5514_ (.A(_1881_),
    .B(_1916_),
    .C(_1950_),
    .D(_1957_),
    .X(_2368_));
 sky130_fd_sc_hd__nand2_1 _5515_ (.A(_1958_),
    .B(_2368_),
    .Y(_2369_));
 sky130_fd_sc_hd__nor2_2 _5516_ (.A(_1757_),
    .B(_1999_),
    .Y(_2370_));
 sky130_fd_sc_hd__and3_1 _5517_ (.A(_1000_),
    .B(_1347_),
    .C(_1564_),
    .X(_2371_));
 sky130_fd_sc_hd__and2_2 _5518_ (.A(\core_1.decode.oc_alu_mode[3] ),
    .B(_1557_),
    .X(_2372_));
 sky130_fd_sc_hd__a221o_1 _5519_ (.A1(_0937_),
    .A2(_1347_),
    .B1(_1564_),
    .B2(_1787_),
    .C1(_2372_),
    .X(_2373_));
 sky130_fd_sc_hd__a211o_1 _5520_ (.A1(_0960_),
    .A2(_1915_),
    .B1(_2371_),
    .C1(_2373_),
    .X(_2374_));
 sky130_fd_sc_hd__a221oi_1 _5521_ (.A1(_0931_),
    .A2(_1916_),
    .B1(_2001_),
    .B2(_2370_),
    .C1(_2374_),
    .Y(_2375_));
 sky130_fd_sc_hd__o221a_1 _5522_ (.A1(_2089_),
    .A2(_1984_),
    .B1(_2088_),
    .B2(_2107_),
    .C1(_2375_),
    .X(_2376_));
 sky130_fd_sc_hd__or2_1 _5523_ (.A(_1913_),
    .B(_1919_),
    .X(_2377_));
 sky130_fd_sc_hd__a21oi_1 _5524_ (.A1(_1913_),
    .A2(_1919_),
    .B1(_2172_),
    .Y(_2378_));
 sky130_fd_sc_hd__nand2_1 _5525_ (.A(_2377_),
    .B(_2378_),
    .Y(_2379_));
 sky130_fd_sc_hd__o211a_1 _5526_ (.A1(_1785_),
    .A2(_2369_),
    .B1(_2376_),
    .C1(_2379_),
    .X(_2380_));
 sky130_fd_sc_hd__nor2_1 _5527_ (.A(_1688_),
    .B(_2380_),
    .Y(_2381_));
 sky130_fd_sc_hd__a211o_2 _5528_ (.A1(_0959_),
    .A2(\core_1.execute.alu_mul_div.mul_res[8] ),
    .B1(_2381_),
    .C1(_0992_),
    .X(_2382_));
 sky130_fd_sc_hd__a22o_2 _5529_ (.A1(\core_1.execute.alu_mul_div.div_cur[8] ),
    .A2(_0964_),
    .B1(_2367_),
    .B2(_2382_),
    .X(_2383_));
 sky130_fd_sc_hd__and2b_1 _5530_ (.A_N(_2338_),
    .B(_2330_),
    .X(_2384_));
 sky130_fd_sc_hd__a22o_1 _5531_ (.A1(\core_1.execute.sreg_scratch.o_d[8] ),
    .A2(_2331_),
    .B1(_2297_),
    .B2(net15),
    .X(_2385_));
 sky130_fd_sc_hd__a221o_1 _5532_ (.A1(\core_1.execute.sreg_priv_control.o_d[8] ),
    .A2(_1162_),
    .B1(_2332_),
    .B2(\core_1.execute.sreg_irq_pc.o_d[8] ),
    .C1(_2385_),
    .X(_2386_));
 sky130_fd_sc_hd__a22o_1 _5533_ (.A1(net86),
    .A2(_2296_),
    .B1(_2386_),
    .B2(_2135_),
    .X(_2387_));
 sky130_fd_sc_hd__mux2_1 _5534_ (.A0(\core_1.execute.sreg_irq_pc.o_d[8] ),
    .A1(_2387_),
    .S(_1799_),
    .X(_2388_));
 sky130_fd_sc_hd__or2_1 _5535_ (.A(_2384_),
    .B(_2388_),
    .X(_2389_));
 sky130_fd_sc_hd__a21oi_1 _5536_ (.A1(_2384_),
    .A2(_2388_),
    .B1(_2116_),
    .Y(_2390_));
 sky130_fd_sc_hd__a22o_1 _5537_ (.A1(_2117_),
    .A2(_2383_),
    .B1(_2389_),
    .B2(_2390_),
    .X(_2391_));
 sky130_fd_sc_hd__mux2_1 _5538_ (.A0(_2391_),
    .A1(net208),
    .S(_1146_),
    .X(_2392_));
 sky130_fd_sc_hd__mux2_1 _5539_ (.A0(\core_1.ew_data[8] ),
    .A1(_2392_),
    .S(_2120_),
    .X(_2393_));
 sky130_fd_sc_hd__clkbuf_1 _5540_ (.A(_2393_),
    .X(_0237_));
 sky130_fd_sc_hd__nand2_1 _5541_ (.A(_2384_),
    .B(_2388_),
    .Y(_2394_));
 sky130_fd_sc_hd__a22o_1 _5542_ (.A1(\core_1.execute.sreg_scratch.o_d[9] ),
    .A2(_2331_),
    .B1(_2297_),
    .B2(net16),
    .X(_2395_));
 sky130_fd_sc_hd__a221o_1 _5543_ (.A1(\core_1.execute.sreg_priv_control.o_d[9] ),
    .A2(_1162_),
    .B1(_2332_),
    .B2(\core_1.execute.sreg_irq_pc.o_d[9] ),
    .C1(_2395_),
    .X(_2396_));
 sky130_fd_sc_hd__a22o_1 _5544_ (.A1(net87),
    .A2(_2296_),
    .B1(_2396_),
    .B2(_2135_),
    .X(_2397_));
 sky130_fd_sc_hd__nand2_1 _5545_ (.A(\core_1.execute.sreg_irq_pc.o_d[9] ),
    .B(\core_1.dec_sreg_irt ),
    .Y(_2398_));
 sky130_fd_sc_hd__a21bo_1 _5546_ (.A1(_1799_),
    .A2(_2397_),
    .B1_N(_2398_),
    .X(_2399_));
 sky130_fd_sc_hd__xnor2_1 _5547_ (.A(_2394_),
    .B(_2399_),
    .Y(_2400_));
 sky130_fd_sc_hd__a21bo_1 _5548_ (.A1(\core_1.execute.alu_mul_div.div_res[9] ),
    .A2(_1685_),
    .B1_N(_0732_),
    .X(_2401_));
 sky130_fd_sc_hd__a21oi_1 _5549_ (.A1(_1914_),
    .A2(_1958_),
    .B1(_1877_),
    .Y(_2402_));
 sky130_fd_sc_hd__a31o_1 _5550_ (.A1(_1877_),
    .A2(_1914_),
    .A3(_1958_),
    .B1(_1785_),
    .X(_2403_));
 sky130_fd_sc_hd__nand3_1 _5551_ (.A(_1880_),
    .B(_1917_),
    .C(_2377_),
    .Y(_2404_));
 sky130_fd_sc_hd__a21o_1 _5552_ (.A1(_1917_),
    .A2(_2377_),
    .B1(_1880_),
    .X(_2405_));
 sky130_fd_sc_hd__inv_2 _5553_ (.A(_1875_),
    .Y(_2406_));
 sky130_fd_sc_hd__a221o_1 _5554_ (.A1(_0937_),
    .A2(_1343_),
    .B1(_1535_),
    .B2(_1787_),
    .C1(_0960_),
    .X(_2407_));
 sky130_fd_sc_hd__inv_2 _5555_ (.A(_1877_),
    .Y(_2408_));
 sky130_fd_sc_hd__a221o_1 _5556_ (.A1(_1000_),
    .A2(_1876_),
    .B1(_2408_),
    .B2(_0931_),
    .C1(_2372_),
    .X(_2409_));
 sky130_fd_sc_hd__nor2_1 _5557_ (.A(_1717_),
    .B(_2107_),
    .Y(_2410_));
 sky130_fd_sc_hd__a211o_1 _5558_ (.A1(_2406_),
    .A2(_2407_),
    .B1(_2409_),
    .C1(_2410_),
    .X(_2411_));
 sky130_fd_sc_hd__and3_1 _5559_ (.A(_1754_),
    .B(_1761_),
    .C(_1765_),
    .X(_2412_));
 sky130_fd_sc_hd__mux2_1 _5560_ (.A0(_1970_),
    .A1(_1986_),
    .S(_1419_),
    .X(_2413_));
 sky130_fd_sc_hd__nor2_1 _5561_ (.A(_2165_),
    .B(_2348_),
    .Y(_2414_));
 sky130_fd_sc_hd__a21oi_1 _5562_ (.A1(_2165_),
    .A2(_2413_),
    .B1(_2414_),
    .Y(_2415_));
 sky130_fd_sc_hd__or2_1 _5563_ (.A(_1764_),
    .B(_2274_),
    .X(_2416_));
 sky130_fd_sc_hd__o211a_1 _5564_ (.A1(_1983_),
    .A2(_2415_),
    .B1(_2416_),
    .C1(_1999_),
    .X(_2417_));
 sky130_fd_sc_hd__o21ba_1 _5565_ (.A1(_2412_),
    .A2(_2417_),
    .B1_N(_1757_),
    .X(_2418_));
 sky130_fd_sc_hd__a311o_1 _5566_ (.A1(_0981_),
    .A2(_2404_),
    .A3(_2405_),
    .B1(_2411_),
    .C1(_2418_),
    .X(_2419_));
 sky130_fd_sc_hd__o21ba_1 _5567_ (.A1(_2402_),
    .A2(_2403_),
    .B1_N(_2419_),
    .X(_2420_));
 sky130_fd_sc_hd__nor2_1 _5568_ (.A(_1688_),
    .B(_2420_),
    .Y(_2421_));
 sky130_fd_sc_hd__a211o_2 _5569_ (.A1(_1688_),
    .A2(\core_1.execute.alu_mul_div.mul_res[9] ),
    .B1(_2421_),
    .C1(_0992_),
    .X(_2422_));
 sky130_fd_sc_hd__a22o_2 _5570_ (.A1(\core_1.execute.alu_mul_div.div_cur[9] ),
    .A2(\core_1.execute.alu_mul_div.i_mod ),
    .B1(_2401_),
    .B2(_2422_),
    .X(_2423_));
 sky130_fd_sc_hd__mux2_1 _5571_ (.A0(_2400_),
    .A1(_2423_),
    .S(_2116_),
    .X(_2424_));
 sky130_fd_sc_hd__mux2_1 _5572_ (.A0(_2424_),
    .A1(net209),
    .S(_1146_),
    .X(_2425_));
 sky130_fd_sc_hd__mux2_1 _5573_ (.A0(\core_1.ew_data[9] ),
    .A1(_2425_),
    .S(_2120_),
    .X(_2426_));
 sky130_fd_sc_hd__clkbuf_1 _5574_ (.A(_2426_),
    .X(_0238_));
 sky130_fd_sc_hd__and3_1 _5575_ (.A(_2384_),
    .B(_2388_),
    .C(_2399_),
    .X(_2427_));
 sky130_fd_sc_hd__a22o_1 _5576_ (.A1(\core_1.execute.sreg_scratch.o_d[10] ),
    .A2(_2331_),
    .B1(_2297_),
    .B2(net2),
    .X(_2428_));
 sky130_fd_sc_hd__a221o_1 _5577_ (.A1(\core_1.execute.sreg_priv_control.o_d[10] ),
    .A2(_1162_),
    .B1(_2332_),
    .B2(\core_1.execute.sreg_irq_pc.o_d[10] ),
    .C1(_2428_),
    .X(_2429_));
 sky130_fd_sc_hd__a22o_1 _5578_ (.A1(net73),
    .A2(_2296_),
    .B1(_2429_),
    .B2(_2135_),
    .X(_2430_));
 sky130_fd_sc_hd__and2_1 _5579_ (.A(\core_1.execute.sreg_irq_pc.o_d[10] ),
    .B(_1057_),
    .X(_2431_));
 sky130_fd_sc_hd__a21oi_1 _5580_ (.A1(_1799_),
    .A2(_2430_),
    .B1(_2431_),
    .Y(_2432_));
 sky130_fd_sc_hd__xnor2_1 _5581_ (.A(_2427_),
    .B(_2432_),
    .Y(_2433_));
 sky130_fd_sc_hd__a21bo_1 _5582_ (.A1(\core_1.execute.alu_mul_div.div_res[10] ),
    .A2(_1685_),
    .B1_N(_0732_),
    .X(_2434_));
 sky130_fd_sc_hd__xor2_1 _5583_ (.A(_1921_),
    .B(_1927_),
    .X(_2435_));
 sky130_fd_sc_hd__o2bb2a_1 _5584_ (.A1_N(_1694_),
    .A2_N(_2161_),
    .B1(_1976_),
    .B2(_1740_),
    .X(_2436_));
 sky130_fd_sc_hd__nor2_1 _5585_ (.A(_1765_),
    .B(_2310_),
    .Y(_2437_));
 sky130_fd_sc_hd__o211a_1 _5586_ (.A1(_1693_),
    .A2(_1970_),
    .B1(_1972_),
    .C1(_1740_),
    .X(_2438_));
 sky130_fd_sc_hd__a21oi_1 _5587_ (.A1(_2165_),
    .A2(_1988_),
    .B1(_2438_),
    .Y(_2439_));
 sky130_fd_sc_hd__o21ai_1 _5588_ (.A1(_1983_),
    .A2(_2439_),
    .B1(_1999_),
    .Y(_2440_));
 sky130_fd_sc_hd__o32a_1 _5589_ (.A1(_1999_),
    .A2(_1983_),
    .A3(_2436_),
    .B1(_2437_),
    .B2(_2440_),
    .X(_2441_));
 sky130_fd_sc_hd__inv_2 _5590_ (.A(\core_1.decode.oc_alu_mode[6] ),
    .Y(_2442_));
 sky130_fd_sc_hd__a221o_1 _5591_ (.A1(\core_1.decode.oc_alu_mode[7] ),
    .A2(_1340_),
    .B1(_1543_),
    .B2(_1787_),
    .C1(_2372_),
    .X(_2443_));
 sky130_fd_sc_hd__a21oi_1 _5592_ (.A1(\core_1.decode.oc_alu_mode[2] ),
    .A2(_1922_),
    .B1(_2443_),
    .Y(_2444_));
 sky130_fd_sc_hd__o221a_1 _5593_ (.A1(_2095_),
    .A2(_1923_),
    .B1(_1924_),
    .B2(_2442_),
    .C1(_2444_),
    .X(_2445_));
 sky130_fd_sc_hd__o21a_1 _5594_ (.A1(_2107_),
    .A2(_2159_),
    .B1(_2445_),
    .X(_2446_));
 sky130_fd_sc_hd__o21ai_1 _5595_ (.A1(_1757_),
    .A2(_2441_),
    .B1(_2446_),
    .Y(_2447_));
 sky130_fd_sc_hd__a31o_1 _5596_ (.A1(_1944_),
    .A2(_1914_),
    .A3(_1958_),
    .B1(_1875_),
    .X(_2448_));
 sky130_fd_sc_hd__nand2_1 _5597_ (.A(_1924_),
    .B(_2448_),
    .Y(_2449_));
 sky130_fd_sc_hd__and3b_1 _5598_ (.A_N(_1959_),
    .B(_2449_),
    .C(_0966_),
    .X(_2450_));
 sky130_fd_sc_hd__a211o_1 _5599_ (.A1(_0981_),
    .A2(_2435_),
    .B1(_2447_),
    .C1(_2450_),
    .X(_2451_));
 sky130_fd_sc_hd__a21o_1 _5600_ (.A1(_0958_),
    .A2(\core_1.execute.alu_mul_div.mul_res[10] ),
    .B1(\core_1.execute.alu_mul_div.i_div ),
    .X(_2452_));
 sky130_fd_sc_hd__a21o_1 _5601_ (.A1(_2081_),
    .A2(_2451_),
    .B1(_2452_),
    .X(_2453_));
 sky130_fd_sc_hd__a22o_2 _5602_ (.A1(\core_1.execute.alu_mul_div.div_cur[10] ),
    .A2(\core_1.execute.alu_mul_div.i_mod ),
    .B1(_2434_),
    .B2(_2453_),
    .X(_2454_));
 sky130_fd_sc_hd__mux2_1 _5603_ (.A0(_2433_),
    .A1(_2454_),
    .S(_2116_),
    .X(_2455_));
 sky130_fd_sc_hd__mux2_1 _5604_ (.A0(_2455_),
    .A1(net195),
    .S(_1146_),
    .X(_2456_));
 sky130_fd_sc_hd__buf_6 _5605_ (.A(_2008_),
    .X(_2457_));
 sky130_fd_sc_hd__mux2_1 _5606_ (.A0(\core_1.ew_data[10] ),
    .A1(_2456_),
    .S(_2457_),
    .X(_2458_));
 sky130_fd_sc_hd__clkbuf_1 _5607_ (.A(_2458_),
    .X(_0239_));
 sky130_fd_sc_hd__inv_2 _5608_ (.A(\core_1.ew_data[11] ),
    .Y(_2459_));
 sky130_fd_sc_hd__a21bo_1 _5609_ (.A1(\core_1.execute.alu_mul_div.div_res[11] ),
    .A2(_1686_),
    .B1_N(_1407_),
    .X(_2460_));
 sky130_fd_sc_hd__o21a_1 _5610_ (.A1(_1922_),
    .A2(_1959_),
    .B1(_1870_),
    .X(_2461_));
 sky130_fd_sc_hd__o31ai_1 _5611_ (.A1(_1870_),
    .A2(_1922_),
    .A3(_1959_),
    .B1(_0966_),
    .Y(_2462_));
 sky130_fd_sc_hd__nor2_1 _5612_ (.A(_1765_),
    .B(_2349_),
    .Y(_2463_));
 sky130_fd_sc_hd__mux2_1 _5613_ (.A0(_1987_),
    .A1(_1989_),
    .S(_1419_),
    .X(_2464_));
 sky130_fd_sc_hd__mux2_1 _5614_ (.A0(_2413_),
    .A1(_2464_),
    .S(_2165_),
    .X(_2465_));
 sky130_fd_sc_hd__a21o_1 _5615_ (.A1(_1764_),
    .A2(_2465_),
    .B1(_1761_),
    .X(_2466_));
 sky130_fd_sc_hd__o32a_1 _5616_ (.A1(_1999_),
    .A2(_1983_),
    .A3(_2210_),
    .B1(_2463_),
    .B2(_2466_),
    .X(_2467_));
 sky130_fd_sc_hd__nor2_2 _5617_ (.A(_1689_),
    .B(_1736_),
    .Y(_2468_));
 sky130_fd_sc_hd__a221o_1 _5618_ (.A1(\core_1.decode.oc_alu_mode[7] ),
    .A2(_1866_),
    .B1(_1586_),
    .B2(_1787_),
    .C1(\core_1.decode.oc_alu_mode[9] ),
    .X(_2469_));
 sky130_fd_sc_hd__a221o_1 _5619_ (.A1(\core_1.decode.oc_alu_mode[2] ),
    .A2(_1869_),
    .B1(_1870_),
    .B2(\core_1.decode.oc_alu_mode[6] ),
    .C1(_2372_),
    .X(_2470_));
 sky130_fd_sc_hd__a221o_1 _5620_ (.A1(_2468_),
    .A2(_2214_),
    .B1(_2469_),
    .B2(_1867_),
    .C1(_2470_),
    .X(_2471_));
 sky130_fd_sc_hd__o21ba_1 _5621_ (.A1(_1757_),
    .A2(_2467_),
    .B1_N(_2471_),
    .X(_2472_));
 sky130_fd_sc_hd__a21oi_1 _5622_ (.A1(_1921_),
    .A2(_1927_),
    .B1(_1925_),
    .Y(_2473_));
 sky130_fd_sc_hd__xnor2_1 _5623_ (.A(_1873_),
    .B(_2473_),
    .Y(_2474_));
 sky130_fd_sc_hd__nand2_1 _5624_ (.A(_0981_),
    .B(_2474_),
    .Y(_2475_));
 sky130_fd_sc_hd__o211a_1 _5625_ (.A1(_2461_),
    .A2(_2462_),
    .B1(_2472_),
    .C1(_2475_),
    .X(_2476_));
 sky130_fd_sc_hd__nor2_1 _5626_ (.A(_0959_),
    .B(_2476_),
    .Y(_2477_));
 sky130_fd_sc_hd__a211o_1 _5627_ (.A1(_0959_),
    .A2(\core_1.execute.alu_mul_div.mul_res[11] ),
    .B1(_2477_),
    .C1(_0992_),
    .X(_2478_));
 sky130_fd_sc_hd__a22o_2 _5628_ (.A1(\core_1.execute.alu_mul_div.div_cur[11] ),
    .A2(_0964_),
    .B1(_2460_),
    .B2(_2478_),
    .X(_2479_));
 sky130_fd_sc_hd__and2b_1 _5629_ (.A_N(_2432_),
    .B(_2427_),
    .X(_2480_));
 sky130_fd_sc_hd__a22o_1 _5630_ (.A1(\core_1.execute.sreg_scratch.o_d[11] ),
    .A2(_2331_),
    .B1(_2297_),
    .B2(net3),
    .X(_2481_));
 sky130_fd_sc_hd__a221o_1 _5631_ (.A1(\core_1.execute.sreg_priv_control.o_d[11] ),
    .A2(_1162_),
    .B1(_2332_),
    .B2(\core_1.execute.sreg_irq_pc.o_d[11] ),
    .C1(_2481_),
    .X(_2482_));
 sky130_fd_sc_hd__a22o_1 _5632_ (.A1(net74),
    .A2(_2296_),
    .B1(_2482_),
    .B2(_2135_),
    .X(_2483_));
 sky130_fd_sc_hd__mux2_1 _5633_ (.A0(\core_1.execute.sreg_irq_pc.o_d[11] ),
    .A1(_2483_),
    .S(_1799_),
    .X(_2484_));
 sky130_fd_sc_hd__nand2_1 _5634_ (.A(_2480_),
    .B(_2484_),
    .Y(_2485_));
 sky130_fd_sc_hd__o21ba_1 _5635_ (.A1(_2480_),
    .A2(_2484_),
    .B1_N(_2117_),
    .X(_2486_));
 sky130_fd_sc_hd__a221oi_1 _5636_ (.A1(_2117_),
    .A2(_2479_),
    .B1(_2485_),
    .B2(_2486_),
    .C1(_1147_),
    .Y(_2487_));
 sky130_fd_sc_hd__a211o_1 _5637_ (.A1(_1147_),
    .A2(_0585_),
    .B1(_1846_),
    .C1(_2487_),
    .X(_2488_));
 sky130_fd_sc_hd__o21ai_1 _5638_ (.A1(_2459_),
    .A2(_2009_),
    .B1(_2488_),
    .Y(_0240_));
 sky130_fd_sc_hd__a22o_1 _5639_ (.A1(\core_1.execute.sreg_scratch.o_d[12] ),
    .A2(_2331_),
    .B1(_2297_),
    .B2(net4),
    .X(_2489_));
 sky130_fd_sc_hd__a221o_1 _5640_ (.A1(\core_1.execute.sreg_priv_control.o_d[12] ),
    .A2(_1162_),
    .B1(_2332_),
    .B2(\core_1.execute.sreg_irq_pc.o_d[12] ),
    .C1(_2489_),
    .X(_2490_));
 sky130_fd_sc_hd__a22o_1 _5641_ (.A1(net75),
    .A2(_2296_),
    .B1(_2490_),
    .B2(_2135_),
    .X(_2491_));
 sky130_fd_sc_hd__nand2_1 _5642_ (.A(\core_1.execute.sreg_irq_pc.o_d[12] ),
    .B(_1057_),
    .Y(_2492_));
 sky130_fd_sc_hd__a21bo_1 _5643_ (.A1(_1799_),
    .A2(_2491_),
    .B1_N(_2492_),
    .X(_2493_));
 sky130_fd_sc_hd__xnor2_1 _5644_ (.A(_2485_),
    .B(_2493_),
    .Y(_2494_));
 sky130_fd_sc_hd__a21bo_1 _5645_ (.A1(\core_1.execute.alu_mul_div.div_res[12] ),
    .A2(_1686_),
    .B1_N(_1407_),
    .X(_2495_));
 sky130_fd_sc_hd__a21oi_1 _5646_ (.A1(_1929_),
    .A2(_1935_),
    .B1(_2172_),
    .Y(_2496_));
 sky130_fd_sc_hd__o21a_1 _5647_ (.A1(_1929_),
    .A2(_1935_),
    .B1(_2496_),
    .X(_2497_));
 sky130_fd_sc_hd__o21a_1 _5648_ (.A1(_1943_),
    .A2(_1959_),
    .B1(_1867_),
    .X(_2498_));
 sky130_fd_sc_hd__nor2_1 _5649_ (.A(_1932_),
    .B(_2498_),
    .Y(_2499_));
 sky130_fd_sc_hd__or3_1 _5650_ (.A(_1785_),
    .B(_1960_),
    .C(_2499_),
    .X(_2500_));
 sky130_fd_sc_hd__inv_2 _5651_ (.A(_1931_),
    .Y(_2501_));
 sky130_fd_sc_hd__a221o_1 _5652_ (.A1(_0937_),
    .A2(_1329_),
    .B1(_2501_),
    .B2(_0960_),
    .C1(_2372_),
    .X(_2502_));
 sky130_fd_sc_hd__a22o_1 _5653_ (.A1(_1580_),
    .A2(_1787_),
    .B1(_1930_),
    .B2(_1000_),
    .X(_2503_));
 sky130_fd_sc_hd__a221o_1 _5654_ (.A1(_0931_),
    .A2(_1932_),
    .B1(_2468_),
    .B2(_2229_),
    .C1(_2503_),
    .X(_2504_));
 sky130_fd_sc_hd__nor2_1 _5655_ (.A(_2502_),
    .B(_2504_),
    .Y(_2505_));
 sky130_fd_sc_hd__mux4_1 _5656_ (.A0(_1969_),
    .A1(_1973_),
    .A2(_1988_),
    .A3(_1991_),
    .S0(_2165_),
    .S1(_1765_),
    .X(_2506_));
 sky130_fd_sc_hd__nor2_1 _5657_ (.A(_1999_),
    .B(_2227_),
    .Y(_2507_));
 sky130_fd_sc_hd__a211o_1 _5658_ (.A1(_1999_),
    .A2(_2506_),
    .B1(_2507_),
    .C1(_1757_),
    .X(_2508_));
 sky130_fd_sc_hd__and4b_1 _5659_ (.A_N(_2497_),
    .B(_2500_),
    .C(_2505_),
    .D(_2508_),
    .X(_2509_));
 sky130_fd_sc_hd__nor2_1 _5660_ (.A(_1688_),
    .B(_2509_),
    .Y(_2510_));
 sky130_fd_sc_hd__a211o_2 _5661_ (.A1(_0959_),
    .A2(\core_1.execute.alu_mul_div.mul_res[12] ),
    .B1(_2510_),
    .C1(_0992_),
    .X(_2511_));
 sky130_fd_sc_hd__a22oi_4 _5662_ (.A1(\core_1.execute.alu_mul_div.div_cur[12] ),
    .A2(_0964_),
    .B1(_2495_),
    .B2(_2511_),
    .Y(_2512_));
 sky130_fd_sc_hd__inv_2 _5663_ (.A(_2512_),
    .Y(_2513_));
 sky130_fd_sc_hd__mux2_1 _5664_ (.A0(_2494_),
    .A1(_2513_),
    .S(_2117_),
    .X(_2514_));
 sky130_fd_sc_hd__nand2_1 _5665_ (.A(_1147_),
    .B(_0577_),
    .Y(_2515_));
 sky130_fd_sc_hd__o211a_1 _5666_ (.A1(_1147_),
    .A2(_2514_),
    .B1(_2515_),
    .C1(_0228_),
    .X(_2516_));
 sky130_fd_sc_hd__a21o_1 _5667_ (.A1(\core_1.ew_data[12] ),
    .A2(_1846_),
    .B1(_2516_),
    .X(_0241_));
 sky130_fd_sc_hd__and3_1 _5668_ (.A(_2480_),
    .B(_2484_),
    .C(_2493_),
    .X(_2517_));
 sky130_fd_sc_hd__a221o_1 _5669_ (.A1(\core_1.execute.sreg_scratch.o_d[13] ),
    .A2(_2331_),
    .B1(_2297_),
    .B2(net5),
    .C1(_2247_),
    .X(_2518_));
 sky130_fd_sc_hd__a221o_1 _5670_ (.A1(\core_1.execute.sreg_priv_control.o_d[13] ),
    .A2(_1162_),
    .B1(_2332_),
    .B2(\core_1.execute.sreg_irq_pc.o_d[13] ),
    .C1(_2518_),
    .X(_2519_));
 sky130_fd_sc_hd__a22o_1 _5671_ (.A1(net76),
    .A2(_2296_),
    .B1(_2519_),
    .B2(_2135_),
    .X(_2520_));
 sky130_fd_sc_hd__and2_1 _5672_ (.A(\core_1.execute.sreg_irq_pc.o_d[13] ),
    .B(_1057_),
    .X(_2521_));
 sky130_fd_sc_hd__a21o_1 _5673_ (.A1(_1799_),
    .A2(_2520_),
    .B1(_2521_),
    .X(_2522_));
 sky130_fd_sc_hd__xor2_1 _5674_ (.A(_2517_),
    .B(_2522_),
    .X(_2523_));
 sky130_fd_sc_hd__a21bo_1 _5675_ (.A1(\core_1.execute.alu_mul_div.div_res[13] ),
    .A2(_1686_),
    .B1_N(_1407_),
    .X(_2524_));
 sky130_fd_sc_hd__a21oi_1 _5676_ (.A1(_1929_),
    .A2(_1935_),
    .B1(_1934_),
    .Y(_2525_));
 sky130_fd_sc_hd__xnor2_1 _5677_ (.A(_1865_),
    .B(_2525_),
    .Y(_2526_));
 sky130_fd_sc_hd__or3_1 _5678_ (.A(_1862_),
    .B(_1930_),
    .C(_1960_),
    .X(_2527_));
 sky130_fd_sc_hd__o21ai_1 _5679_ (.A1(_1930_),
    .A2(_1960_),
    .B1(_1862_),
    .Y(_2528_));
 sky130_fd_sc_hd__a221o_1 _5680_ (.A1(\core_1.decode.oc_alu_mode[7] ),
    .A2(_1699_),
    .B1(_1854_),
    .B2(_1787_),
    .C1(_2372_),
    .X(_2529_));
 sky130_fd_sc_hd__a221o_1 _5681_ (.A1(\core_1.decode.oc_alu_mode[9] ),
    .A2(_1859_),
    .B1(_1861_),
    .B2(\core_1.decode.oc_alu_mode[2] ),
    .C1(_2529_),
    .X(_2530_));
 sky130_fd_sc_hd__a21o_1 _5682_ (.A1(\core_1.decode.oc_alu_mode[6] ),
    .A2(_1862_),
    .B1(_2530_),
    .X(_2531_));
 sky130_fd_sc_hd__a21o_1 _5683_ (.A1(_2468_),
    .A2(_2283_),
    .B1(_2531_),
    .X(_2532_));
 sky130_fd_sc_hd__a21o_1 _5684_ (.A1(_2275_),
    .A2(_2370_),
    .B1(_2532_),
    .X(_2533_));
 sky130_fd_sc_hd__mux2_1 _5685_ (.A0(_1990_),
    .A1(_1993_),
    .S(_1419_),
    .X(_2534_));
 sky130_fd_sc_hd__mux2_1 _5686_ (.A0(_2464_),
    .A1(_2534_),
    .S(_2165_),
    .X(_2535_));
 sky130_fd_sc_hd__nand2_1 _5687_ (.A(_1765_),
    .B(_2535_),
    .Y(_2536_));
 sky130_fd_sc_hd__o211a_1 _5688_ (.A1(_1765_),
    .A2(_2415_),
    .B1(_2536_),
    .C1(_1762_),
    .X(_2537_));
 sky130_fd_sc_hd__a311o_1 _5689_ (.A1(_0966_),
    .A2(_2527_),
    .A3(_2528_),
    .B1(_2533_),
    .C1(_2537_),
    .X(_2538_));
 sky130_fd_sc_hd__a21oi_2 _5690_ (.A1(_0981_),
    .A2(_2526_),
    .B1(_2538_),
    .Y(_2539_));
 sky130_fd_sc_hd__nor2_1 _5691_ (.A(_1688_),
    .B(_2539_),
    .Y(_2540_));
 sky130_fd_sc_hd__a211o_1 _5692_ (.A1(_0959_),
    .A2(\core_1.execute.alu_mul_div.mul_res[13] ),
    .B1(_2540_),
    .C1(_0992_),
    .X(_2541_));
 sky130_fd_sc_hd__a22o_4 _5693_ (.A1(\core_1.execute.alu_mul_div.div_cur[13] ),
    .A2(_0964_),
    .B1(_2524_),
    .B2(_2541_),
    .X(_2542_));
 sky130_fd_sc_hd__mux2_1 _5694_ (.A0(_2523_),
    .A1(_2542_),
    .S(_2116_),
    .X(_2543_));
 sky130_fd_sc_hd__mux2_1 _5695_ (.A0(_2543_),
    .A1(net198),
    .S(_1146_),
    .X(_2544_));
 sky130_fd_sc_hd__mux2_1 _5696_ (.A0(\core_1.ew_data[13] ),
    .A1(_2544_),
    .S(_2457_),
    .X(_2545_));
 sky130_fd_sc_hd__clkbuf_1 _5697_ (.A(_2545_),
    .X(_0242_));
 sky130_fd_sc_hd__nand2_1 _5698_ (.A(_2517_),
    .B(_2522_),
    .Y(_2546_));
 sky130_fd_sc_hd__a221o_1 _5699_ (.A1(\core_1.execute.sreg_scratch.o_d[14] ),
    .A2(_2331_),
    .B1(_2297_),
    .B2(net6),
    .C1(_2247_),
    .X(_2547_));
 sky130_fd_sc_hd__a221o_1 _5700_ (.A1(\core_1.execute.sreg_priv_control.o_d[14] ),
    .A2(_1162_),
    .B1(_2332_),
    .B2(\core_1.execute.sreg_irq_pc.o_d[14] ),
    .C1(_2547_),
    .X(_2548_));
 sky130_fd_sc_hd__a22o_1 _5701_ (.A1(net77),
    .A2(_2296_),
    .B1(_2548_),
    .B2(_2135_),
    .X(_2549_));
 sky130_fd_sc_hd__nand2_1 _5702_ (.A(\core_1.execute.sreg_irq_pc.o_d[14] ),
    .B(_1057_),
    .Y(_2550_));
 sky130_fd_sc_hd__a21bo_1 _5703_ (.A1(_1799_),
    .A2(_2549_),
    .B1_N(_2550_),
    .X(_2551_));
 sky130_fd_sc_hd__xnor2_1 _5704_ (.A(_2546_),
    .B(_2551_),
    .Y(_2552_));
 sky130_fd_sc_hd__o31a_1 _5705_ (.A1(_1861_),
    .A2(_1930_),
    .A3(_1960_),
    .B1(_1859_),
    .X(_2553_));
 sky130_fd_sc_hd__nor2_1 _5706_ (.A(_1857_),
    .B(_2553_),
    .Y(_2554_));
 sky130_fd_sc_hd__a21oi_1 _5707_ (.A1(_1938_),
    .A2(_1858_),
    .B1(_1937_),
    .Y(_2555_));
 sky130_fd_sc_hd__a31o_1 _5708_ (.A1(_1938_),
    .A2(_1858_),
    .A3(_1937_),
    .B1(_2172_),
    .X(_2556_));
 sky130_fd_sc_hd__mux2_1 _5709_ (.A0(_1991_),
    .A1(_1995_),
    .S(_1982_),
    .X(_2557_));
 sky130_fd_sc_hd__inv_2 _5710_ (.A(_2557_),
    .Y(_2558_));
 sky130_fd_sc_hd__mux2_1 _5711_ (.A0(_2439_),
    .A1(_2558_),
    .S(_1764_),
    .X(_2559_));
 sky130_fd_sc_hd__inv_2 _5712_ (.A(_1856_),
    .Y(_2560_));
 sky130_fd_sc_hd__a221o_1 _5713_ (.A1(\core_1.decode.oc_alu_mode[7] ),
    .A2(_1323_),
    .B1(_2560_),
    .B2(\core_1.decode.oc_alu_mode[9] ),
    .C1(_2372_),
    .X(_2561_));
 sky130_fd_sc_hd__a221o_1 _5714_ (.A1(\core_1.decode.oc_alu_mode[2] ),
    .A2(_1855_),
    .B1(_1857_),
    .B2(\core_1.decode.oc_alu_mode[6] ),
    .C1(_2561_),
    .X(_2562_));
 sky130_fd_sc_hd__a221o_1 _5715_ (.A1(_1594_),
    .A2(_1787_),
    .B1(_2468_),
    .B2(_2315_),
    .C1(_2562_),
    .X(_2563_));
 sky130_fd_sc_hd__a221o_1 _5716_ (.A1(_2311_),
    .A2(_2370_),
    .B1(_2559_),
    .B2(_1762_),
    .C1(_2563_),
    .X(_2564_));
 sky130_fd_sc_hd__o21ba_1 _5717_ (.A1(_2555_),
    .A2(_2556_),
    .B1_N(_2564_),
    .X(_2565_));
 sky130_fd_sc_hd__o31ai_4 _5718_ (.A1(_1785_),
    .A2(_1961_),
    .A3(_2554_),
    .B1(_2565_),
    .Y(_2566_));
 sky130_fd_sc_hd__a21o_1 _5719_ (.A1(_0958_),
    .A2(\core_1.execute.alu_mul_div.mul_res[14] ),
    .B1(\core_1.execute.alu_mul_div.i_div ),
    .X(_2567_));
 sky130_fd_sc_hd__a21oi_1 _5720_ (.A1(_2081_),
    .A2(_2566_),
    .B1(_2567_),
    .Y(_2568_));
 sky130_fd_sc_hd__a21boi_1 _5721_ (.A1(\core_1.execute.alu_mul_div.div_res[14] ),
    .A2(_1685_),
    .B1_N(_0732_),
    .Y(_2569_));
 sky130_fd_sc_hd__o2bb2a_2 _5722_ (.A1_N(\core_1.execute.alu_mul_div.div_cur[14] ),
    .A2_N(\core_1.execute.alu_mul_div.i_mod ),
    .B1(_2568_),
    .B2(_2569_),
    .X(_2570_));
 sky130_fd_sc_hd__clkinv_2 _5723_ (.A(_2570_),
    .Y(_2571_));
 sky130_fd_sc_hd__mux2_1 _5724_ (.A0(_2552_),
    .A1(_2571_),
    .S(_2116_),
    .X(_2572_));
 sky130_fd_sc_hd__mux2_1 _5725_ (.A0(_2572_),
    .A1(net199),
    .S(_1146_),
    .X(_2573_));
 sky130_fd_sc_hd__mux2_1 _5726_ (.A0(\core_1.ew_data[14] ),
    .A1(_2573_),
    .S(_2457_),
    .X(_2574_));
 sky130_fd_sc_hd__clkbuf_1 _5727_ (.A(_2574_),
    .X(_0243_));
 sky130_fd_sc_hd__or2b_1 _5728_ (.A(_2546_),
    .B_N(_2551_),
    .X(_2575_));
 sky130_fd_sc_hd__a221o_1 _5729_ (.A1(\core_1.execute.sreg_scratch.o_d[15] ),
    .A2(_2331_),
    .B1(_2297_),
    .B2(net7),
    .C1(_2247_),
    .X(_2576_));
 sky130_fd_sc_hd__a221o_1 _5730_ (.A1(\core_1.execute.sreg_priv_control.o_d[15] ),
    .A2(_1162_),
    .B1(_2332_),
    .B2(\core_1.execute.sreg_irq_pc.o_d[15] ),
    .C1(_2576_),
    .X(_2577_));
 sky130_fd_sc_hd__a22o_1 _5731_ (.A1(net78),
    .A2(_2296_),
    .B1(_2577_),
    .B2(_2135_),
    .X(_2578_));
 sky130_fd_sc_hd__mux2_1 _5732_ (.A0(\core_1.execute.sreg_irq_pc.o_d[15] ),
    .A1(_2578_),
    .S(_1799_),
    .X(_2579_));
 sky130_fd_sc_hd__xnor2_1 _5733_ (.A(_2575_),
    .B(_2579_),
    .Y(_2580_));
 sky130_fd_sc_hd__nor2_1 _5734_ (.A(_1853_),
    .B(_1940_),
    .Y(_2581_));
 sky130_fd_sc_hd__xnor2_1 _5735_ (.A(_1939_),
    .B(_2581_),
    .Y(_2582_));
 sky130_fd_sc_hd__a21o_1 _5736_ (.A1(\core_1.decode.oc_alu_mode[2] ),
    .A2(_1529_),
    .B1(_0937_),
    .X(_2583_));
 sky130_fd_sc_hd__a221o_1 _5737_ (.A1(_0960_),
    .A2(_1962_),
    .B1(_2583_),
    .B2(_1849_),
    .C1(_2372_),
    .X(_2584_));
 sky130_fd_sc_hd__a32o_1 _5738_ (.A1(_1384_),
    .A2(_2468_),
    .A3(_2353_),
    .B1(_1852_),
    .B2(_0931_),
    .X(_2585_));
 sky130_fd_sc_hd__nor2_1 _5739_ (.A(_2584_),
    .B(_2585_),
    .Y(_2586_));
 sky130_fd_sc_hd__nor2_1 _5740_ (.A(_1693_),
    .B(_1996_),
    .Y(_2587_));
 sky130_fd_sc_hd__a211o_1 _5741_ (.A1(_1693_),
    .A2(_1994_),
    .B1(_2587_),
    .C1(_1740_),
    .X(_2588_));
 sky130_fd_sc_hd__o211a_1 _5742_ (.A1(_2165_),
    .A2(_2534_),
    .B1(_2588_),
    .C1(_1765_),
    .X(_2589_));
 sky130_fd_sc_hd__a211o_1 _5743_ (.A1(_1983_),
    .A2(_2465_),
    .B1(_2589_),
    .C1(_2089_),
    .X(_2590_));
 sky130_fd_sc_hd__o311a_2 _5744_ (.A1(_1757_),
    .A2(_1999_),
    .A3(_2351_),
    .B1(_2586_),
    .C1(_2590_),
    .X(_2591_));
 sky130_fd_sc_hd__o21ai_1 _5745_ (.A1(_1855_),
    .A2(_1961_),
    .B1(_1852_),
    .Y(_2592_));
 sky130_fd_sc_hd__o31a_1 _5746_ (.A1(_1852_),
    .A2(_1855_),
    .A3(_1961_),
    .B1(_0966_),
    .X(_2593_));
 sky130_fd_sc_hd__nand2_1 _5747_ (.A(_2592_),
    .B(_2593_),
    .Y(_2594_));
 sky130_fd_sc_hd__o211a_1 _5748_ (.A1(_2172_),
    .A2(_2582_),
    .B1(_2591_),
    .C1(_2594_),
    .X(_2595_));
 sky130_fd_sc_hd__a21bo_2 _5749_ (.A1(_1529_),
    .A2(_1787_),
    .B1_N(_2595_),
    .X(_2596_));
 sky130_fd_sc_hd__a21o_1 _5750_ (.A1(_0958_),
    .A2(\core_1.execute.alu_mul_div.mul_res[15] ),
    .B1(\core_1.execute.alu_mul_div.i_div ),
    .X(_2597_));
 sky130_fd_sc_hd__a21o_1 _5751_ (.A1(_2081_),
    .A2(_2596_),
    .B1(_2597_),
    .X(_2598_));
 sky130_fd_sc_hd__a21bo_1 _5752_ (.A1(\core_1.execute.alu_mul_div.div_res[15] ),
    .A2(_1685_),
    .B1_N(_0732_),
    .X(_2599_));
 sky130_fd_sc_hd__a22o_4 _5753_ (.A1(\core_1.execute.alu_mul_div.div_cur[15] ),
    .A2(\core_1.execute.alu_mul_div.i_mod ),
    .B1(_2598_),
    .B2(_2599_),
    .X(_2600_));
 sky130_fd_sc_hd__mux2_1 _5754_ (.A0(_2580_),
    .A1(_2600_),
    .S(_2116_),
    .X(_2601_));
 sky130_fd_sc_hd__mux2_1 _5755_ (.A0(_2601_),
    .A1(net200),
    .S(_1146_),
    .X(_2602_));
 sky130_fd_sc_hd__mux2_1 _5756_ (.A0(\core_1.ew_data[15] ),
    .A1(_2602_),
    .S(_2457_),
    .X(_2603_));
 sky130_fd_sc_hd__clkbuf_1 _5757_ (.A(_2603_),
    .X(_0244_));
 sky130_fd_sc_hd__mux2_1 _5758_ (.A0(\core_1.ew_addr[0] ),
    .A1(_2114_),
    .S(_2457_),
    .X(_2604_));
 sky130_fd_sc_hd__clkbuf_1 _5759_ (.A(_2604_),
    .X(_0245_));
 sky130_fd_sc_hd__mux2_1 _5760_ (.A0(net116),
    .A1(_1797_),
    .S(_2457_),
    .X(_2605_));
 sky130_fd_sc_hd__clkbuf_1 _5761_ (.A(_2605_),
    .X(_0246_));
 sky130_fd_sc_hd__mux2_1 _5762_ (.A0(net123),
    .A1(_2182_),
    .S(_2457_),
    .X(_2606_));
 sky130_fd_sc_hd__clkbuf_1 _5763_ (.A(_2606_),
    .X(_0247_));
 sky130_fd_sc_hd__mux2_1 _5764_ (.A0(net124),
    .A1(_2219_),
    .S(_2457_),
    .X(_2607_));
 sky130_fd_sc_hd__clkbuf_1 _5765_ (.A(_2607_),
    .X(_0248_));
 sky130_fd_sc_hd__mux2_1 _5766_ (.A0(net125),
    .A1(_2246_),
    .S(_2457_),
    .X(_2608_));
 sky130_fd_sc_hd__clkbuf_1 _5767_ (.A(_2608_),
    .X(_0249_));
 sky130_fd_sc_hd__mux2_1 _5768_ (.A0(net126),
    .A1(_2292_),
    .S(_2457_),
    .X(_2609_));
 sky130_fd_sc_hd__clkbuf_1 _5769_ (.A(_2609_),
    .X(_0250_));
 sky130_fd_sc_hd__buf_4 _5770_ (.A(_2008_),
    .X(_2610_));
 sky130_fd_sc_hd__mux2_1 _5771_ (.A0(net127),
    .A1(_2326_),
    .S(_2610_),
    .X(_2611_));
 sky130_fd_sc_hd__clkbuf_1 _5772_ (.A(_2611_),
    .X(_0251_));
 sky130_fd_sc_hd__mux2_1 _5773_ (.A0(net128),
    .A1(_2363_),
    .S(_2610_),
    .X(_2612_));
 sky130_fd_sc_hd__clkbuf_1 _5774_ (.A(_2612_),
    .X(_0252_));
 sky130_fd_sc_hd__mux2_1 _5775_ (.A0(net129),
    .A1(_2383_),
    .S(_2610_),
    .X(_2613_));
 sky130_fd_sc_hd__clkbuf_1 _5776_ (.A(_2613_),
    .X(_0253_));
 sky130_fd_sc_hd__mux2_1 _5777_ (.A0(net130),
    .A1(_2423_),
    .S(_2610_),
    .X(_2614_));
 sky130_fd_sc_hd__clkbuf_1 _5778_ (.A(_2614_),
    .X(_0254_));
 sky130_fd_sc_hd__mux2_1 _5779_ (.A0(net131),
    .A1(_2454_),
    .S(_2610_),
    .X(_2615_));
 sky130_fd_sc_hd__clkbuf_1 _5780_ (.A(_2615_),
    .X(_0255_));
 sky130_fd_sc_hd__mux2_1 _5781_ (.A0(net117),
    .A1(_2479_),
    .S(_2610_),
    .X(_2616_));
 sky130_fd_sc_hd__clkbuf_1 _5782_ (.A(_2616_),
    .X(_0256_));
 sky130_fd_sc_hd__mux2_1 _5783_ (.A0(net118),
    .A1(_2513_),
    .S(_2610_),
    .X(_2617_));
 sky130_fd_sc_hd__clkbuf_1 _5784_ (.A(_2617_),
    .X(_0257_));
 sky130_fd_sc_hd__mux2_1 _5785_ (.A0(net119),
    .A1(_2542_),
    .S(_2610_),
    .X(_2618_));
 sky130_fd_sc_hd__clkbuf_1 _5786_ (.A(_2618_),
    .X(_0258_));
 sky130_fd_sc_hd__mux2_1 _5787_ (.A0(net120),
    .A1(_2571_),
    .S(_2610_),
    .X(_2619_));
 sky130_fd_sc_hd__clkbuf_1 _5788_ (.A(_2619_),
    .X(_0259_));
 sky130_fd_sc_hd__mux2_1 _5789_ (.A0(net121),
    .A1(_2600_),
    .S(_2610_),
    .X(_2620_));
 sky130_fd_sc_hd__clkbuf_1 _5790_ (.A(_2620_),
    .X(_0260_));
 sky130_fd_sc_hd__mux2_1 _5791_ (.A0(\core_1.dec_rf_ie[0] ),
    .A1(\core_1.ew_reg_ie[0] ),
    .S(_1846_),
    .X(_2621_));
 sky130_fd_sc_hd__clkbuf_1 _5792_ (.A(_2621_),
    .X(_0261_));
 sky130_fd_sc_hd__mux2_1 _5793_ (.A0(\core_1.dec_rf_ie[1] ),
    .A1(\core_1.ew_reg_ie[1] ),
    .S(_1846_),
    .X(_2622_));
 sky130_fd_sc_hd__clkbuf_1 _5794_ (.A(_2622_),
    .X(_0262_));
 sky130_fd_sc_hd__mux2_1 _5795_ (.A0(\core_1.dec_rf_ie[2] ),
    .A1(\core_1.ew_reg_ie[2] ),
    .S(_1846_),
    .X(_2623_));
 sky130_fd_sc_hd__clkbuf_1 _5796_ (.A(_2623_),
    .X(_0263_));
 sky130_fd_sc_hd__mux2_1 _5797_ (.A0(\core_1.dec_rf_ie[3] ),
    .A1(\core_1.ew_reg_ie[3] ),
    .S(_1846_),
    .X(_2624_));
 sky130_fd_sc_hd__clkbuf_1 _5798_ (.A(_2624_),
    .X(_0264_));
 sky130_fd_sc_hd__mux2_1 _5799_ (.A0(\core_1.dec_rf_ie[4] ),
    .A1(\core_1.ew_reg_ie[4] ),
    .S(_1846_),
    .X(_2625_));
 sky130_fd_sc_hd__clkbuf_1 _5800_ (.A(_2625_),
    .X(_0265_));
 sky130_fd_sc_hd__mux2_1 _5801_ (.A0(\core_1.dec_rf_ie[5] ),
    .A1(\core_1.ew_reg_ie[5] ),
    .S(_1845_),
    .X(_2626_));
 sky130_fd_sc_hd__clkbuf_1 _5802_ (.A(_2626_),
    .X(_0266_));
 sky130_fd_sc_hd__mux2_1 _5803_ (.A0(\core_1.dec_rf_ie[6] ),
    .A1(\core_1.ew_reg_ie[6] ),
    .S(_1845_),
    .X(_2627_));
 sky130_fd_sc_hd__clkbuf_1 _5804_ (.A(_2627_),
    .X(_0267_));
 sky130_fd_sc_hd__mux2_1 _5805_ (.A0(\core_1.dec_rf_ie[7] ),
    .A1(\core_1.ew_reg_ie[7] ),
    .S(_1845_),
    .X(_2628_));
 sky130_fd_sc_hd__clkbuf_1 _5806_ (.A(_2628_),
    .X(_0268_));
 sky130_fd_sc_hd__mux2_1 _5807_ (.A0(_1147_),
    .A1(_1310_),
    .S(_1845_),
    .X(_2629_));
 sky130_fd_sc_hd__clkbuf_1 _5808_ (.A(_2629_),
    .X(_0269_));
 sky130_fd_sc_hd__mux2_1 _5809_ (.A0(\core_1.dec_mem_width ),
    .A1(\core_1.ew_mem_width ),
    .S(_1845_),
    .X(_2630_));
 sky130_fd_sc_hd__clkbuf_1 _5810_ (.A(_2630_),
    .X(_0270_));
 sky130_fd_sc_hd__and3_1 _5811_ (.A(\core_1.execute.sreg_long_ptr_en ),
    .B(\core_1.dec_mem_long ),
    .C(_2009_),
    .X(_2631_));
 sky130_fd_sc_hd__a21o_1 _5812_ (.A1(net155),
    .A2(_1846_),
    .B1(_2631_),
    .X(_0271_));
 sky130_fd_sc_hd__nor2_1 _5813_ (.A(_1128_),
    .B(_1158_),
    .Y(_0272_));
 sky130_fd_sc_hd__mux2_2 _5814_ (.A0(\core_1.ew_submit ),
    .A1(net20),
    .S(\core_1.ew_mem_access ),
    .X(_2632_));
 sky130_fd_sc_hd__buf_6 _5815_ (.A(_2632_),
    .X(_2633_));
 sky130_fd_sc_hd__nand2_4 _5816_ (.A(\core_1.ew_reg_ie[7] ),
    .B(_2633_),
    .Y(_2634_));
 sky130_fd_sc_hd__mux2_1 _5817_ (.A0(net35),
    .A1(net21),
    .S(_1008_),
    .X(_2635_));
 sky130_fd_sc_hd__mux2_1 _5818_ (.A0(\core_1.ew_data[0] ),
    .A1(_2635_),
    .S(_1309_),
    .X(_2636_));
 sky130_fd_sc_hd__buf_4 _5819_ (.A(_2636_),
    .X(_2637_));
 sky130_fd_sc_hd__and2_2 _5820_ (.A(\core_1.ew_reg_ie[7] ),
    .B(_2632_),
    .X(_2638_));
 sky130_fd_sc_hd__buf_4 _5821_ (.A(_2638_),
    .X(_2639_));
 sky130_fd_sc_hd__or2_1 _5822_ (.A(\core_1.execute.rf.reg_outputs[7][0] ),
    .B(_2639_),
    .X(_2640_));
 sky130_fd_sc_hd__o211a_1 _5823_ (.A1(_2634_),
    .A2(_2637_),
    .B1(_2640_),
    .C1(_1834_),
    .X(_0273_));
 sky130_fd_sc_hd__mux2_1 _5824_ (.A0(net36),
    .A1(net28),
    .S(_1008_),
    .X(_2641_));
 sky130_fd_sc_hd__mux2_1 _5825_ (.A0(\core_1.ew_data[1] ),
    .A1(_2641_),
    .S(_1309_),
    .X(_2642_));
 sky130_fd_sc_hd__clkbuf_4 _5826_ (.A(_2642_),
    .X(_2643_));
 sky130_fd_sc_hd__or2_1 _5827_ (.A(\core_1.execute.rf.reg_outputs[7][1] ),
    .B(_2639_),
    .X(_2644_));
 sky130_fd_sc_hd__buf_4 _5828_ (.A(_1307_),
    .X(_2645_));
 sky130_fd_sc_hd__o211a_1 _5829_ (.A1(_2634_),
    .A2(_2643_),
    .B1(_2644_),
    .C1(_2645_),
    .X(_0274_));
 sky130_fd_sc_hd__mux2_1 _5830_ (.A0(net22),
    .A1(net29),
    .S(_1007_),
    .X(_2646_));
 sky130_fd_sc_hd__mux2_1 _5831_ (.A0(\core_1.ew_data[2] ),
    .A1(_2646_),
    .S(_1309_),
    .X(_2647_));
 sky130_fd_sc_hd__clkbuf_4 _5832_ (.A(_2647_),
    .X(_2648_));
 sky130_fd_sc_hd__or2_1 _5833_ (.A(\core_1.execute.rf.reg_outputs[7][2] ),
    .B(_2639_),
    .X(_2649_));
 sky130_fd_sc_hd__o211a_1 _5834_ (.A1(_2634_),
    .A2(_2648_),
    .B1(_2649_),
    .C1(_2645_),
    .X(_0275_));
 sky130_fd_sc_hd__mux2_1 _5835_ (.A0(net23),
    .A1(net30),
    .S(_1007_),
    .X(_2650_));
 sky130_fd_sc_hd__mux2_1 _5836_ (.A0(\core_1.ew_data[3] ),
    .A1(_2650_),
    .S(_1309_),
    .X(_2651_));
 sky130_fd_sc_hd__buf_4 _5837_ (.A(_2651_),
    .X(_2652_));
 sky130_fd_sc_hd__or2_1 _5838_ (.A(\core_1.execute.rf.reg_outputs[7][3] ),
    .B(_2639_),
    .X(_2653_));
 sky130_fd_sc_hd__o211a_1 _5839_ (.A1(_2634_),
    .A2(_2652_),
    .B1(_2653_),
    .C1(_2645_),
    .X(_0276_));
 sky130_fd_sc_hd__mux2_1 _5840_ (.A0(net24),
    .A1(net31),
    .S(_1007_),
    .X(_2654_));
 sky130_fd_sc_hd__mux2_1 _5841_ (.A0(\core_1.ew_data[4] ),
    .A1(_2654_),
    .S(_1309_),
    .X(_2655_));
 sky130_fd_sc_hd__buf_2 _5842_ (.A(_2655_),
    .X(_2656_));
 sky130_fd_sc_hd__or2_1 _5843_ (.A(\core_1.execute.rf.reg_outputs[7][4] ),
    .B(_2638_),
    .X(_2657_));
 sky130_fd_sc_hd__o211a_1 _5844_ (.A1(_2634_),
    .A2(_2656_),
    .B1(_2657_),
    .C1(_2645_),
    .X(_0277_));
 sky130_fd_sc_hd__mux2_1 _5845_ (.A0(net25),
    .A1(net32),
    .S(_1007_),
    .X(_2658_));
 sky130_fd_sc_hd__mux2_1 _5846_ (.A0(\core_1.ew_data[5] ),
    .A1(_2658_),
    .S(_1309_),
    .X(_2659_));
 sky130_fd_sc_hd__buf_2 _5847_ (.A(_2659_),
    .X(_2660_));
 sky130_fd_sc_hd__or2_1 _5848_ (.A(\core_1.execute.rf.reg_outputs[7][5] ),
    .B(_2638_),
    .X(_2661_));
 sky130_fd_sc_hd__o211a_1 _5849_ (.A1(_2634_),
    .A2(_2660_),
    .B1(_2661_),
    .C1(_2645_),
    .X(_0278_));
 sky130_fd_sc_hd__mux2_1 _5850_ (.A0(net26),
    .A1(net33),
    .S(_1007_),
    .X(_2662_));
 sky130_fd_sc_hd__mux2_1 _5851_ (.A0(\core_1.ew_data[6] ),
    .A1(_2662_),
    .S(_1309_),
    .X(_2663_));
 sky130_fd_sc_hd__clkbuf_4 _5852_ (.A(_2663_),
    .X(_2664_));
 sky130_fd_sc_hd__or2_1 _5853_ (.A(\core_1.execute.rf.reg_outputs[7][6] ),
    .B(_2638_),
    .X(_2665_));
 sky130_fd_sc_hd__o211a_1 _5854_ (.A1(_2634_),
    .A2(_2664_),
    .B1(_2665_),
    .C1(_2645_),
    .X(_0279_));
 sky130_fd_sc_hd__mux2_1 _5855_ (.A0(net27),
    .A1(net34),
    .S(_1007_),
    .X(_2666_));
 sky130_fd_sc_hd__mux2_1 _5856_ (.A0(\core_1.ew_data[7] ),
    .A1(_2666_),
    .S(_1309_),
    .X(_2667_));
 sky130_fd_sc_hd__clkbuf_4 _5857_ (.A(_2667_),
    .X(_2668_));
 sky130_fd_sc_hd__or2_1 _5858_ (.A(\core_1.execute.rf.reg_outputs[7][7] ),
    .B(_2638_),
    .X(_2669_));
 sky130_fd_sc_hd__o211a_1 _5859_ (.A1(_2634_),
    .A2(_2668_),
    .B1(_2669_),
    .C1(_2645_),
    .X(_0280_));
 sky130_fd_sc_hd__buf_4 _5860_ (.A(_2638_),
    .X(_2670_));
 sky130_fd_sc_hd__and2b_1 _5861_ (.A_N(\core_1.ew_mem_width ),
    .B(_1309_),
    .X(_2671_));
 sky130_fd_sc_hd__buf_4 _5862_ (.A(_2671_),
    .X(_2672_));
 sky130_fd_sc_hd__inv_2 _5863_ (.A(\core_1.ew_data[8] ),
    .Y(_2673_));
 sky130_fd_sc_hd__o2bb2a_4 _5864_ (.A1_N(net35),
    .A2_N(_2672_),
    .B1(_2673_),
    .B2(_1310_),
    .X(_2674_));
 sky130_fd_sc_hd__nand2_1 _5865_ (.A(_2670_),
    .B(_2674_),
    .Y(_2675_));
 sky130_fd_sc_hd__o211a_1 _5866_ (.A1(\core_1.execute.rf.reg_outputs[7][8] ),
    .A2(_2670_),
    .B1(_2675_),
    .C1(_2645_),
    .X(_0281_));
 sky130_fd_sc_hd__inv_2 _5867_ (.A(\core_1.ew_data[9] ),
    .Y(_2676_));
 sky130_fd_sc_hd__o2bb2a_4 _5868_ (.A1_N(net36),
    .A2_N(_2672_),
    .B1(_2676_),
    .B2(_1310_),
    .X(_2677_));
 sky130_fd_sc_hd__nand2_1 _5869_ (.A(_2670_),
    .B(_2677_),
    .Y(_2678_));
 sky130_fd_sc_hd__o211a_1 _5870_ (.A1(\core_1.execute.rf.reg_outputs[7][9] ),
    .A2(_2670_),
    .B1(_2678_),
    .C1(_2645_),
    .X(_0282_));
 sky130_fd_sc_hd__inv_2 _5871_ (.A(\core_1.ew_data[10] ),
    .Y(_2679_));
 sky130_fd_sc_hd__o2bb2a_4 _5872_ (.A1_N(net22),
    .A2_N(_2672_),
    .B1(_2679_),
    .B2(_1310_),
    .X(_2680_));
 sky130_fd_sc_hd__nand2_1 _5873_ (.A(_2639_),
    .B(_2680_),
    .Y(_2681_));
 sky130_fd_sc_hd__o211a_1 _5874_ (.A1(\core_1.execute.rf.reg_outputs[7][10] ),
    .A2(_2670_),
    .B1(_2681_),
    .C1(_2645_),
    .X(_0283_));
 sky130_fd_sc_hd__o2bb2a_4 _5875_ (.A1_N(net23),
    .A2_N(_2672_),
    .B1(_2459_),
    .B2(_1310_),
    .X(_2682_));
 sky130_fd_sc_hd__nand2_1 _5876_ (.A(_2639_),
    .B(_2682_),
    .Y(_2683_));
 sky130_fd_sc_hd__buf_4 _5877_ (.A(_1307_),
    .X(_2684_));
 sky130_fd_sc_hd__o211a_1 _5878_ (.A1(\core_1.execute.rf.reg_outputs[7][11] ),
    .A2(_2670_),
    .B1(_2683_),
    .C1(_2684_),
    .X(_0284_));
 sky130_fd_sc_hd__inv_2 _5879_ (.A(\core_1.ew_data[12] ),
    .Y(_2685_));
 sky130_fd_sc_hd__o2bb2a_4 _5880_ (.A1_N(net24),
    .A2_N(_2672_),
    .B1(_2685_),
    .B2(_1310_),
    .X(_2686_));
 sky130_fd_sc_hd__nand2_1 _5881_ (.A(_2639_),
    .B(_2686_),
    .Y(_2687_));
 sky130_fd_sc_hd__o211a_1 _5882_ (.A1(\core_1.execute.rf.reg_outputs[7][12] ),
    .A2(_2670_),
    .B1(_2687_),
    .C1(_2684_),
    .X(_0285_));
 sky130_fd_sc_hd__inv_2 _5883_ (.A(\core_1.ew_data[13] ),
    .Y(_2688_));
 sky130_fd_sc_hd__o2bb2a_4 _5884_ (.A1_N(net25),
    .A2_N(_2672_),
    .B1(_2688_),
    .B2(_1310_),
    .X(_2689_));
 sky130_fd_sc_hd__nand2_1 _5885_ (.A(_2639_),
    .B(_2689_),
    .Y(_2690_));
 sky130_fd_sc_hd__o211a_1 _5886_ (.A1(\core_1.execute.rf.reg_outputs[7][13] ),
    .A2(_2670_),
    .B1(_2690_),
    .C1(_2684_),
    .X(_0286_));
 sky130_fd_sc_hd__inv_2 _5887_ (.A(\core_1.ew_data[14] ),
    .Y(_2691_));
 sky130_fd_sc_hd__o2bb2a_4 _5888_ (.A1_N(net26),
    .A2_N(_2672_),
    .B1(_2691_),
    .B2(_1310_),
    .X(_2692_));
 sky130_fd_sc_hd__nand2_1 _5889_ (.A(_2639_),
    .B(_2692_),
    .Y(_2693_));
 sky130_fd_sc_hd__o211a_1 _5890_ (.A1(\core_1.execute.rf.reg_outputs[7][14] ),
    .A2(_2670_),
    .B1(_2693_),
    .C1(_2684_),
    .X(_0287_));
 sky130_fd_sc_hd__inv_2 _5891_ (.A(\core_1.ew_data[15] ),
    .Y(_2694_));
 sky130_fd_sc_hd__o2bb2a_4 _5892_ (.A1_N(net27),
    .A2_N(_2672_),
    .B1(_2694_),
    .B2(_1310_),
    .X(_2695_));
 sky130_fd_sc_hd__nand2_1 _5893_ (.A(_2639_),
    .B(_2695_),
    .Y(_2696_));
 sky130_fd_sc_hd__o211a_1 _5894_ (.A1(\core_1.execute.rf.reg_outputs[7][15] ),
    .A2(_2670_),
    .B1(_2696_),
    .C1(_2684_),
    .X(_0288_));
 sky130_fd_sc_hd__nand2_4 _5895_ (.A(\core_1.ew_reg_ie[6] ),
    .B(_2633_),
    .Y(_2697_));
 sky130_fd_sc_hd__and2_2 _5896_ (.A(\core_1.ew_reg_ie[6] ),
    .B(_2633_),
    .X(_2698_));
 sky130_fd_sc_hd__buf_4 _5897_ (.A(_2698_),
    .X(_2699_));
 sky130_fd_sc_hd__or2_1 _5898_ (.A(\core_1.execute.rf.reg_outputs[6][0] ),
    .B(_2699_),
    .X(_2700_));
 sky130_fd_sc_hd__o211a_1 _5899_ (.A1(_2637_),
    .A2(_2697_),
    .B1(_2700_),
    .C1(_2684_),
    .X(_0289_));
 sky130_fd_sc_hd__or2_1 _5900_ (.A(\core_1.execute.rf.reg_outputs[6][1] ),
    .B(_2699_),
    .X(_2701_));
 sky130_fd_sc_hd__o211a_1 _5901_ (.A1(_2643_),
    .A2(_2697_),
    .B1(_2701_),
    .C1(_2684_),
    .X(_0290_));
 sky130_fd_sc_hd__or2_1 _5902_ (.A(\core_1.execute.rf.reg_outputs[6][2] ),
    .B(_2699_),
    .X(_2702_));
 sky130_fd_sc_hd__o211a_1 _5903_ (.A1(_2648_),
    .A2(_2697_),
    .B1(_2702_),
    .C1(_2684_),
    .X(_0291_));
 sky130_fd_sc_hd__or2_1 _5904_ (.A(\core_1.execute.rf.reg_outputs[6][3] ),
    .B(_2699_),
    .X(_2703_));
 sky130_fd_sc_hd__o211a_1 _5905_ (.A1(_2652_),
    .A2(_2697_),
    .B1(_2703_),
    .C1(_2684_),
    .X(_0292_));
 sky130_fd_sc_hd__or2_1 _5906_ (.A(\core_1.execute.rf.reg_outputs[6][4] ),
    .B(_2698_),
    .X(_2704_));
 sky130_fd_sc_hd__o211a_1 _5907_ (.A1(_2656_),
    .A2(_2697_),
    .B1(_2704_),
    .C1(_2684_),
    .X(_0293_));
 sky130_fd_sc_hd__or2_1 _5908_ (.A(\core_1.execute.rf.reg_outputs[6][5] ),
    .B(_2698_),
    .X(_2705_));
 sky130_fd_sc_hd__buf_4 _5909_ (.A(_1307_),
    .X(_2706_));
 sky130_fd_sc_hd__o211a_1 _5910_ (.A1(_2660_),
    .A2(_2697_),
    .B1(_2705_),
    .C1(_2706_),
    .X(_0294_));
 sky130_fd_sc_hd__or2_1 _5911_ (.A(\core_1.execute.rf.reg_outputs[6][6] ),
    .B(_2698_),
    .X(_2707_));
 sky130_fd_sc_hd__o211a_1 _5912_ (.A1(_2664_),
    .A2(_2697_),
    .B1(_2707_),
    .C1(_2706_),
    .X(_0295_));
 sky130_fd_sc_hd__or2_1 _5913_ (.A(\core_1.execute.rf.reg_outputs[6][7] ),
    .B(_2698_),
    .X(_2708_));
 sky130_fd_sc_hd__o211a_1 _5914_ (.A1(_2668_),
    .A2(_2697_),
    .B1(_2708_),
    .C1(_2706_),
    .X(_0296_));
 sky130_fd_sc_hd__buf_4 _5915_ (.A(_2698_),
    .X(_2709_));
 sky130_fd_sc_hd__nand2_1 _5916_ (.A(_2674_),
    .B(_2709_),
    .Y(_2710_));
 sky130_fd_sc_hd__o211a_1 _5917_ (.A1(\core_1.execute.rf.reg_outputs[6][8] ),
    .A2(_2709_),
    .B1(_2710_),
    .C1(_2706_),
    .X(_0297_));
 sky130_fd_sc_hd__nand2_1 _5918_ (.A(_2677_),
    .B(_2709_),
    .Y(_2711_));
 sky130_fd_sc_hd__o211a_1 _5919_ (.A1(\core_1.execute.rf.reg_outputs[6][9] ),
    .A2(_2709_),
    .B1(_2711_),
    .C1(_2706_),
    .X(_0298_));
 sky130_fd_sc_hd__nand2_1 _5920_ (.A(_2680_),
    .B(_2699_),
    .Y(_2712_));
 sky130_fd_sc_hd__o211a_1 _5921_ (.A1(\core_1.execute.rf.reg_outputs[6][10] ),
    .A2(_2709_),
    .B1(_2712_),
    .C1(_2706_),
    .X(_0299_));
 sky130_fd_sc_hd__nand2_1 _5922_ (.A(_2682_),
    .B(_2699_),
    .Y(_2713_));
 sky130_fd_sc_hd__o211a_1 _5923_ (.A1(\core_1.execute.rf.reg_outputs[6][11] ),
    .A2(_2709_),
    .B1(_2713_),
    .C1(_2706_),
    .X(_0300_));
 sky130_fd_sc_hd__nand2_1 _5924_ (.A(_2686_),
    .B(_2699_),
    .Y(_2714_));
 sky130_fd_sc_hd__o211a_1 _5925_ (.A1(\core_1.execute.rf.reg_outputs[6][12] ),
    .A2(_2709_),
    .B1(_2714_),
    .C1(_2706_),
    .X(_0301_));
 sky130_fd_sc_hd__nand2_1 _5926_ (.A(_2689_),
    .B(_2699_),
    .Y(_2715_));
 sky130_fd_sc_hd__o211a_1 _5927_ (.A1(\core_1.execute.rf.reg_outputs[6][13] ),
    .A2(_2709_),
    .B1(_2715_),
    .C1(_2706_),
    .X(_0302_));
 sky130_fd_sc_hd__nand2_1 _5928_ (.A(_2692_),
    .B(_2699_),
    .Y(_2716_));
 sky130_fd_sc_hd__o211a_1 _5929_ (.A1(\core_1.execute.rf.reg_outputs[6][14] ),
    .A2(_2709_),
    .B1(_2716_),
    .C1(_2706_),
    .X(_0303_));
 sky130_fd_sc_hd__nand2_1 _5930_ (.A(_2695_),
    .B(_2699_),
    .Y(_2717_));
 sky130_fd_sc_hd__clkbuf_4 _5931_ (.A(_0662_),
    .X(_2718_));
 sky130_fd_sc_hd__buf_4 _5932_ (.A(_2718_),
    .X(_2719_));
 sky130_fd_sc_hd__o211a_1 _5933_ (.A1(\core_1.execute.rf.reg_outputs[6][15] ),
    .A2(_2709_),
    .B1(_2717_),
    .C1(_2719_),
    .X(_0304_));
 sky130_fd_sc_hd__nand2_4 _5934_ (.A(\core_1.ew_reg_ie[5] ),
    .B(_2633_),
    .Y(_2720_));
 sky130_fd_sc_hd__and2_2 _5935_ (.A(\core_1.ew_reg_ie[5] ),
    .B(_2633_),
    .X(_2721_));
 sky130_fd_sc_hd__buf_4 _5936_ (.A(_2721_),
    .X(_2722_));
 sky130_fd_sc_hd__or2_1 _5937_ (.A(\core_1.execute.rf.reg_outputs[5][0] ),
    .B(_2722_),
    .X(_2723_));
 sky130_fd_sc_hd__o211a_1 _5938_ (.A1(_2637_),
    .A2(_2720_),
    .B1(_2723_),
    .C1(_2719_),
    .X(_0305_));
 sky130_fd_sc_hd__or2_1 _5939_ (.A(\core_1.execute.rf.reg_outputs[5][1] ),
    .B(_2722_),
    .X(_2724_));
 sky130_fd_sc_hd__o211a_1 _5940_ (.A1(_2643_),
    .A2(_2720_),
    .B1(_2724_),
    .C1(_2719_),
    .X(_0306_));
 sky130_fd_sc_hd__or2_1 _5941_ (.A(\core_1.execute.rf.reg_outputs[5][2] ),
    .B(_2722_),
    .X(_2725_));
 sky130_fd_sc_hd__o211a_1 _5942_ (.A1(_2648_),
    .A2(_2720_),
    .B1(_2725_),
    .C1(_2719_),
    .X(_0307_));
 sky130_fd_sc_hd__or2_1 _5943_ (.A(\core_1.execute.rf.reg_outputs[5][3] ),
    .B(_2722_),
    .X(_2726_));
 sky130_fd_sc_hd__o211a_1 _5944_ (.A1(_2652_),
    .A2(_2720_),
    .B1(_2726_),
    .C1(_2719_),
    .X(_0308_));
 sky130_fd_sc_hd__or2_1 _5945_ (.A(\core_1.execute.rf.reg_outputs[5][4] ),
    .B(_2721_),
    .X(_2727_));
 sky130_fd_sc_hd__o211a_1 _5946_ (.A1(_2656_),
    .A2(_2720_),
    .B1(_2727_),
    .C1(_2719_),
    .X(_0309_));
 sky130_fd_sc_hd__or2_1 _5947_ (.A(\core_1.execute.rf.reg_outputs[5][5] ),
    .B(_2721_),
    .X(_2728_));
 sky130_fd_sc_hd__o211a_1 _5948_ (.A1(_2660_),
    .A2(_2720_),
    .B1(_2728_),
    .C1(_2719_),
    .X(_0310_));
 sky130_fd_sc_hd__or2_1 _5949_ (.A(\core_1.execute.rf.reg_outputs[5][6] ),
    .B(_2721_),
    .X(_2729_));
 sky130_fd_sc_hd__o211a_1 _5950_ (.A1(_2664_),
    .A2(_2720_),
    .B1(_2729_),
    .C1(_2719_),
    .X(_0311_));
 sky130_fd_sc_hd__or2_1 _5951_ (.A(\core_1.execute.rf.reg_outputs[5][7] ),
    .B(_2721_),
    .X(_2730_));
 sky130_fd_sc_hd__o211a_1 _5952_ (.A1(_2668_),
    .A2(_2720_),
    .B1(_2730_),
    .C1(_2719_),
    .X(_0312_));
 sky130_fd_sc_hd__buf_4 _5953_ (.A(_2721_),
    .X(_2731_));
 sky130_fd_sc_hd__nand2_1 _5954_ (.A(_2674_),
    .B(_2731_),
    .Y(_2732_));
 sky130_fd_sc_hd__o211a_1 _5955_ (.A1(\core_1.execute.rf.reg_outputs[5][8] ),
    .A2(_2731_),
    .B1(_2732_),
    .C1(_2719_),
    .X(_0313_));
 sky130_fd_sc_hd__nand2_1 _5956_ (.A(_2677_),
    .B(_2731_),
    .Y(_2733_));
 sky130_fd_sc_hd__buf_4 _5957_ (.A(_2718_),
    .X(_2734_));
 sky130_fd_sc_hd__o211a_1 _5958_ (.A1(\core_1.execute.rf.reg_outputs[5][9] ),
    .A2(_2731_),
    .B1(_2733_),
    .C1(_2734_),
    .X(_0314_));
 sky130_fd_sc_hd__nand2_1 _5959_ (.A(_2680_),
    .B(_2722_),
    .Y(_2735_));
 sky130_fd_sc_hd__o211a_1 _5960_ (.A1(\core_1.execute.rf.reg_outputs[5][10] ),
    .A2(_2731_),
    .B1(_2735_),
    .C1(_2734_),
    .X(_0315_));
 sky130_fd_sc_hd__nand2_1 _5961_ (.A(_2682_),
    .B(_2722_),
    .Y(_2736_));
 sky130_fd_sc_hd__o211a_1 _5962_ (.A1(\core_1.execute.rf.reg_outputs[5][11] ),
    .A2(_2731_),
    .B1(_2736_),
    .C1(_2734_),
    .X(_0316_));
 sky130_fd_sc_hd__nand2_1 _5963_ (.A(_2686_),
    .B(_2722_),
    .Y(_2737_));
 sky130_fd_sc_hd__o211a_1 _5964_ (.A1(\core_1.execute.rf.reg_outputs[5][12] ),
    .A2(_2731_),
    .B1(_2737_),
    .C1(_2734_),
    .X(_0317_));
 sky130_fd_sc_hd__nand2_1 _5965_ (.A(_2689_),
    .B(_2722_),
    .Y(_2738_));
 sky130_fd_sc_hd__o211a_1 _5966_ (.A1(\core_1.execute.rf.reg_outputs[5][13] ),
    .A2(_2731_),
    .B1(_2738_),
    .C1(_2734_),
    .X(_0318_));
 sky130_fd_sc_hd__nand2_1 _5967_ (.A(_2692_),
    .B(_2722_),
    .Y(_2739_));
 sky130_fd_sc_hd__o211a_1 _5968_ (.A1(\core_1.execute.rf.reg_outputs[5][14] ),
    .A2(_2731_),
    .B1(_2739_),
    .C1(_2734_),
    .X(_0319_));
 sky130_fd_sc_hd__nand2_1 _5969_ (.A(_2695_),
    .B(_2722_),
    .Y(_2740_));
 sky130_fd_sc_hd__o211a_1 _5970_ (.A1(\core_1.execute.rf.reg_outputs[5][15] ),
    .A2(_2731_),
    .B1(_2740_),
    .C1(_2734_),
    .X(_0320_));
 sky130_fd_sc_hd__nand2_4 _5971_ (.A(\core_1.ew_reg_ie[4] ),
    .B(_2633_),
    .Y(_2741_));
 sky130_fd_sc_hd__and2_2 _5972_ (.A(\core_1.ew_reg_ie[4] ),
    .B(_2632_),
    .X(_2742_));
 sky130_fd_sc_hd__buf_4 _5973_ (.A(_2742_),
    .X(_2743_));
 sky130_fd_sc_hd__or2_1 _5974_ (.A(\core_1.execute.rf.reg_outputs[4][0] ),
    .B(_2743_),
    .X(_2744_));
 sky130_fd_sc_hd__o211a_1 _5975_ (.A1(_2637_),
    .A2(_2741_),
    .B1(_2744_),
    .C1(_2734_),
    .X(_0321_));
 sky130_fd_sc_hd__or2_1 _5976_ (.A(\core_1.execute.rf.reg_outputs[4][1] ),
    .B(_2743_),
    .X(_2745_));
 sky130_fd_sc_hd__o211a_1 _5977_ (.A1(_2643_),
    .A2(_2741_),
    .B1(_2745_),
    .C1(_2734_),
    .X(_0322_));
 sky130_fd_sc_hd__or2_1 _5978_ (.A(\core_1.execute.rf.reg_outputs[4][2] ),
    .B(_2743_),
    .X(_2746_));
 sky130_fd_sc_hd__o211a_1 _5979_ (.A1(_2648_),
    .A2(_2741_),
    .B1(_2746_),
    .C1(_2734_),
    .X(_0323_));
 sky130_fd_sc_hd__or2_1 _5980_ (.A(\core_1.execute.rf.reg_outputs[4][3] ),
    .B(_2743_),
    .X(_2747_));
 sky130_fd_sc_hd__buf_4 _5981_ (.A(_2718_),
    .X(_2748_));
 sky130_fd_sc_hd__o211a_1 _5982_ (.A1(_2652_),
    .A2(_2741_),
    .B1(_2747_),
    .C1(_2748_),
    .X(_0324_));
 sky130_fd_sc_hd__or2_1 _5983_ (.A(\core_1.execute.rf.reg_outputs[4][4] ),
    .B(_2742_),
    .X(_2749_));
 sky130_fd_sc_hd__o211a_1 _5984_ (.A1(_2656_),
    .A2(_2741_),
    .B1(_2749_),
    .C1(_2748_),
    .X(_0325_));
 sky130_fd_sc_hd__or2_1 _5985_ (.A(\core_1.execute.rf.reg_outputs[4][5] ),
    .B(_2742_),
    .X(_2750_));
 sky130_fd_sc_hd__o211a_1 _5986_ (.A1(_2660_),
    .A2(_2741_),
    .B1(_2750_),
    .C1(_2748_),
    .X(_0326_));
 sky130_fd_sc_hd__or2_1 _5987_ (.A(\core_1.execute.rf.reg_outputs[4][6] ),
    .B(_2742_),
    .X(_2751_));
 sky130_fd_sc_hd__o211a_1 _5988_ (.A1(_2664_),
    .A2(_2741_),
    .B1(_2751_),
    .C1(_2748_),
    .X(_0327_));
 sky130_fd_sc_hd__or2_1 _5989_ (.A(\core_1.execute.rf.reg_outputs[4][7] ),
    .B(_2742_),
    .X(_2752_));
 sky130_fd_sc_hd__o211a_1 _5990_ (.A1(_2668_),
    .A2(_2741_),
    .B1(_2752_),
    .C1(_2748_),
    .X(_0328_));
 sky130_fd_sc_hd__clkbuf_4 _5991_ (.A(_2742_),
    .X(_2753_));
 sky130_fd_sc_hd__nand2_1 _5992_ (.A(_2674_),
    .B(_2753_),
    .Y(_2754_));
 sky130_fd_sc_hd__o211a_1 _5993_ (.A1(\core_1.execute.rf.reg_outputs[4][8] ),
    .A2(_2753_),
    .B1(_2754_),
    .C1(_2748_),
    .X(_0329_));
 sky130_fd_sc_hd__nand2_1 _5994_ (.A(_2677_),
    .B(_2753_),
    .Y(_2755_));
 sky130_fd_sc_hd__o211a_1 _5995_ (.A1(\core_1.execute.rf.reg_outputs[4][9] ),
    .A2(_2753_),
    .B1(_2755_),
    .C1(_2748_),
    .X(_0330_));
 sky130_fd_sc_hd__nand2_1 _5996_ (.A(_2680_),
    .B(_2743_),
    .Y(_2756_));
 sky130_fd_sc_hd__o211a_1 _5997_ (.A1(\core_1.execute.rf.reg_outputs[4][10] ),
    .A2(_2753_),
    .B1(_2756_),
    .C1(_2748_),
    .X(_0331_));
 sky130_fd_sc_hd__nand2_1 _5998_ (.A(_2682_),
    .B(_2743_),
    .Y(_2757_));
 sky130_fd_sc_hd__o211a_1 _5999_ (.A1(\core_1.execute.rf.reg_outputs[4][11] ),
    .A2(_2753_),
    .B1(_2757_),
    .C1(_2748_),
    .X(_0332_));
 sky130_fd_sc_hd__nand2_1 _6000_ (.A(_2686_),
    .B(_2743_),
    .Y(_2758_));
 sky130_fd_sc_hd__o211a_1 _6001_ (.A1(\core_1.execute.rf.reg_outputs[4][12] ),
    .A2(_2753_),
    .B1(_2758_),
    .C1(_2748_),
    .X(_0333_));
 sky130_fd_sc_hd__nand2_1 _6002_ (.A(_2689_),
    .B(_2743_),
    .Y(_2759_));
 sky130_fd_sc_hd__buf_4 _6003_ (.A(_2718_),
    .X(_2760_));
 sky130_fd_sc_hd__o211a_1 _6004_ (.A1(\core_1.execute.rf.reg_outputs[4][13] ),
    .A2(_2753_),
    .B1(_2759_),
    .C1(_2760_),
    .X(_0334_));
 sky130_fd_sc_hd__nand2_1 _6005_ (.A(_2692_),
    .B(_2743_),
    .Y(_2761_));
 sky130_fd_sc_hd__o211a_1 _6006_ (.A1(\core_1.execute.rf.reg_outputs[4][14] ),
    .A2(_2753_),
    .B1(_2761_),
    .C1(_2760_),
    .X(_0335_));
 sky130_fd_sc_hd__nand2_1 _6007_ (.A(_2695_),
    .B(_2743_),
    .Y(_2762_));
 sky130_fd_sc_hd__o211a_1 _6008_ (.A1(\core_1.execute.rf.reg_outputs[4][15] ),
    .A2(_2753_),
    .B1(_2762_),
    .C1(_2760_),
    .X(_0336_));
 sky130_fd_sc_hd__nand2_4 _6009_ (.A(\core_1.ew_reg_ie[3] ),
    .B(_2633_),
    .Y(_2763_));
 sky130_fd_sc_hd__and2_2 _6010_ (.A(\core_1.ew_reg_ie[3] ),
    .B(_2632_),
    .X(_2764_));
 sky130_fd_sc_hd__buf_4 _6011_ (.A(_2764_),
    .X(_2765_));
 sky130_fd_sc_hd__or2_1 _6012_ (.A(\core_1.execute.rf.reg_outputs[3][0] ),
    .B(_2765_),
    .X(_2766_));
 sky130_fd_sc_hd__o211a_1 _6013_ (.A1(_2637_),
    .A2(_2763_),
    .B1(_2766_),
    .C1(_2760_),
    .X(_0337_));
 sky130_fd_sc_hd__or2_1 _6014_ (.A(\core_1.execute.rf.reg_outputs[3][1] ),
    .B(_2765_),
    .X(_2767_));
 sky130_fd_sc_hd__o211a_1 _6015_ (.A1(_2643_),
    .A2(_2763_),
    .B1(_2767_),
    .C1(_2760_),
    .X(_0338_));
 sky130_fd_sc_hd__or2_1 _6016_ (.A(\core_1.execute.rf.reg_outputs[3][2] ),
    .B(_2765_),
    .X(_2768_));
 sky130_fd_sc_hd__o211a_1 _6017_ (.A1(_2648_),
    .A2(_2763_),
    .B1(_2768_),
    .C1(_2760_),
    .X(_0339_));
 sky130_fd_sc_hd__or2_1 _6018_ (.A(\core_1.execute.rf.reg_outputs[3][3] ),
    .B(_2765_),
    .X(_2769_));
 sky130_fd_sc_hd__o211a_1 _6019_ (.A1(_2652_),
    .A2(_2763_),
    .B1(_2769_),
    .C1(_2760_),
    .X(_0340_));
 sky130_fd_sc_hd__or2_1 _6020_ (.A(\core_1.execute.rf.reg_outputs[3][4] ),
    .B(_2764_),
    .X(_2770_));
 sky130_fd_sc_hd__o211a_1 _6021_ (.A1(_2656_),
    .A2(_2763_),
    .B1(_2770_),
    .C1(_2760_),
    .X(_0341_));
 sky130_fd_sc_hd__or2_1 _6022_ (.A(\core_1.execute.rf.reg_outputs[3][5] ),
    .B(_2764_),
    .X(_2771_));
 sky130_fd_sc_hd__o211a_1 _6023_ (.A1(_2660_),
    .A2(_2763_),
    .B1(_2771_),
    .C1(_2760_),
    .X(_0342_));
 sky130_fd_sc_hd__or2_1 _6024_ (.A(\core_1.execute.rf.reg_outputs[3][6] ),
    .B(_2764_),
    .X(_2772_));
 sky130_fd_sc_hd__o211a_1 _6025_ (.A1(_2664_),
    .A2(_2763_),
    .B1(_2772_),
    .C1(_2760_),
    .X(_0343_));
 sky130_fd_sc_hd__or2_1 _6026_ (.A(\core_1.execute.rf.reg_outputs[3][7] ),
    .B(_2764_),
    .X(_2773_));
 sky130_fd_sc_hd__buf_4 _6027_ (.A(_2718_),
    .X(_2774_));
 sky130_fd_sc_hd__o211a_1 _6028_ (.A1(_2668_),
    .A2(_2763_),
    .B1(_2773_),
    .C1(_2774_),
    .X(_0344_));
 sky130_fd_sc_hd__clkbuf_4 _6029_ (.A(_2764_),
    .X(_2775_));
 sky130_fd_sc_hd__nand2_1 _6030_ (.A(_2674_),
    .B(_2775_),
    .Y(_2776_));
 sky130_fd_sc_hd__o211a_1 _6031_ (.A1(\core_1.execute.rf.reg_outputs[3][8] ),
    .A2(_2775_),
    .B1(_2776_),
    .C1(_2774_),
    .X(_0345_));
 sky130_fd_sc_hd__nand2_1 _6032_ (.A(_2677_),
    .B(_2775_),
    .Y(_2777_));
 sky130_fd_sc_hd__o211a_1 _6033_ (.A1(\core_1.execute.rf.reg_outputs[3][9] ),
    .A2(_2775_),
    .B1(_2777_),
    .C1(_2774_),
    .X(_0346_));
 sky130_fd_sc_hd__nand2_1 _6034_ (.A(_2680_),
    .B(_2765_),
    .Y(_2778_));
 sky130_fd_sc_hd__o211a_1 _6035_ (.A1(\core_1.execute.rf.reg_outputs[3][10] ),
    .A2(_2775_),
    .B1(_2778_),
    .C1(_2774_),
    .X(_0347_));
 sky130_fd_sc_hd__nand2_1 _6036_ (.A(_2682_),
    .B(_2765_),
    .Y(_2779_));
 sky130_fd_sc_hd__o211a_1 _6037_ (.A1(\core_1.execute.rf.reg_outputs[3][11] ),
    .A2(_2775_),
    .B1(_2779_),
    .C1(_2774_),
    .X(_0348_));
 sky130_fd_sc_hd__nand2_1 _6038_ (.A(_2686_),
    .B(_2765_),
    .Y(_2780_));
 sky130_fd_sc_hd__o211a_1 _6039_ (.A1(\core_1.execute.rf.reg_outputs[3][12] ),
    .A2(_2775_),
    .B1(_2780_),
    .C1(_2774_),
    .X(_0349_));
 sky130_fd_sc_hd__nand2_1 _6040_ (.A(_2689_),
    .B(_2765_),
    .Y(_2781_));
 sky130_fd_sc_hd__o211a_1 _6041_ (.A1(\core_1.execute.rf.reg_outputs[3][13] ),
    .A2(_2775_),
    .B1(_2781_),
    .C1(_2774_),
    .X(_0350_));
 sky130_fd_sc_hd__nand2_1 _6042_ (.A(_2692_),
    .B(_2765_),
    .Y(_2782_));
 sky130_fd_sc_hd__o211a_1 _6043_ (.A1(\core_1.execute.rf.reg_outputs[3][14] ),
    .A2(_2775_),
    .B1(_2782_),
    .C1(_2774_),
    .X(_0351_));
 sky130_fd_sc_hd__nand2_1 _6044_ (.A(_2695_),
    .B(_2765_),
    .Y(_2783_));
 sky130_fd_sc_hd__o211a_1 _6045_ (.A1(\core_1.execute.rf.reg_outputs[3][15] ),
    .A2(_2775_),
    .B1(_2783_),
    .C1(_2774_),
    .X(_0352_));
 sky130_fd_sc_hd__nand2_4 _6046_ (.A(\core_1.ew_reg_ie[2] ),
    .B(_2633_),
    .Y(_2784_));
 sky130_fd_sc_hd__and2_2 _6047_ (.A(\core_1.ew_reg_ie[2] ),
    .B(_2632_),
    .X(_2785_));
 sky130_fd_sc_hd__buf_4 _6048_ (.A(_2785_),
    .X(_2786_));
 sky130_fd_sc_hd__or2_1 _6049_ (.A(\core_1.execute.rf.reg_outputs[2][0] ),
    .B(_2786_),
    .X(_2787_));
 sky130_fd_sc_hd__o211a_1 _6050_ (.A1(_2637_),
    .A2(_2784_),
    .B1(_2787_),
    .C1(_2774_),
    .X(_0353_));
 sky130_fd_sc_hd__or2_1 _6051_ (.A(\core_1.execute.rf.reg_outputs[2][1] ),
    .B(_2786_),
    .X(_2788_));
 sky130_fd_sc_hd__buf_4 _6052_ (.A(_2718_),
    .X(_2789_));
 sky130_fd_sc_hd__o211a_1 _6053_ (.A1(_2643_),
    .A2(_2784_),
    .B1(_2788_),
    .C1(_2789_),
    .X(_0354_));
 sky130_fd_sc_hd__or2_1 _6054_ (.A(\core_1.execute.rf.reg_outputs[2][2] ),
    .B(_2786_),
    .X(_2790_));
 sky130_fd_sc_hd__o211a_1 _6055_ (.A1(_2648_),
    .A2(_2784_),
    .B1(_2790_),
    .C1(_2789_),
    .X(_0355_));
 sky130_fd_sc_hd__or2_1 _6056_ (.A(\core_1.execute.rf.reg_outputs[2][3] ),
    .B(_2786_),
    .X(_2791_));
 sky130_fd_sc_hd__o211a_1 _6057_ (.A1(_2652_),
    .A2(_2784_),
    .B1(_2791_),
    .C1(_2789_),
    .X(_0356_));
 sky130_fd_sc_hd__or2_1 _6058_ (.A(\core_1.execute.rf.reg_outputs[2][4] ),
    .B(_2785_),
    .X(_2792_));
 sky130_fd_sc_hd__o211a_1 _6059_ (.A1(_2656_),
    .A2(_2784_),
    .B1(_2792_),
    .C1(_2789_),
    .X(_0357_));
 sky130_fd_sc_hd__or2_1 _6060_ (.A(\core_1.execute.rf.reg_outputs[2][5] ),
    .B(_2785_),
    .X(_2793_));
 sky130_fd_sc_hd__o211a_1 _6061_ (.A1(_2660_),
    .A2(_2784_),
    .B1(_2793_),
    .C1(_2789_),
    .X(_0358_));
 sky130_fd_sc_hd__or2_1 _6062_ (.A(\core_1.execute.rf.reg_outputs[2][6] ),
    .B(_2785_),
    .X(_2794_));
 sky130_fd_sc_hd__o211a_1 _6063_ (.A1(_2664_),
    .A2(_2784_),
    .B1(_2794_),
    .C1(_2789_),
    .X(_0359_));
 sky130_fd_sc_hd__or2_1 _6064_ (.A(\core_1.execute.rf.reg_outputs[2][7] ),
    .B(_2785_),
    .X(_2795_));
 sky130_fd_sc_hd__o211a_1 _6065_ (.A1(_2668_),
    .A2(_2784_),
    .B1(_2795_),
    .C1(_2789_),
    .X(_0360_));
 sky130_fd_sc_hd__clkbuf_4 _6066_ (.A(_2785_),
    .X(_2796_));
 sky130_fd_sc_hd__nand2_1 _6067_ (.A(_2674_),
    .B(_2796_),
    .Y(_2797_));
 sky130_fd_sc_hd__o211a_1 _6068_ (.A1(\core_1.execute.rf.reg_outputs[2][8] ),
    .A2(_2796_),
    .B1(_2797_),
    .C1(_2789_),
    .X(_0361_));
 sky130_fd_sc_hd__nand2_1 _6069_ (.A(_2677_),
    .B(_2796_),
    .Y(_2798_));
 sky130_fd_sc_hd__o211a_1 _6070_ (.A1(\core_1.execute.rf.reg_outputs[2][9] ),
    .A2(_2796_),
    .B1(_2798_),
    .C1(_2789_),
    .X(_0362_));
 sky130_fd_sc_hd__nand2_1 _6071_ (.A(_2680_),
    .B(_2786_),
    .Y(_2799_));
 sky130_fd_sc_hd__o211a_1 _6072_ (.A1(\core_1.execute.rf.reg_outputs[2][10] ),
    .A2(_2796_),
    .B1(_2799_),
    .C1(_2789_),
    .X(_0363_));
 sky130_fd_sc_hd__nand2_1 _6073_ (.A(_2682_),
    .B(_2786_),
    .Y(_2800_));
 sky130_fd_sc_hd__buf_4 _6074_ (.A(_2718_),
    .X(_2801_));
 sky130_fd_sc_hd__o211a_1 _6075_ (.A1(\core_1.execute.rf.reg_outputs[2][11] ),
    .A2(_2796_),
    .B1(_2800_),
    .C1(_2801_),
    .X(_0364_));
 sky130_fd_sc_hd__nand2_1 _6076_ (.A(_2686_),
    .B(_2786_),
    .Y(_2802_));
 sky130_fd_sc_hd__o211a_1 _6077_ (.A1(\core_1.execute.rf.reg_outputs[2][12] ),
    .A2(_2796_),
    .B1(_2802_),
    .C1(_2801_),
    .X(_0365_));
 sky130_fd_sc_hd__nand2_1 _6078_ (.A(_2689_),
    .B(_2786_),
    .Y(_2803_));
 sky130_fd_sc_hd__o211a_1 _6079_ (.A1(\core_1.execute.rf.reg_outputs[2][13] ),
    .A2(_2796_),
    .B1(_2803_),
    .C1(_2801_),
    .X(_0366_));
 sky130_fd_sc_hd__nand2_1 _6080_ (.A(_2692_),
    .B(_2786_),
    .Y(_2804_));
 sky130_fd_sc_hd__o211a_1 _6081_ (.A1(\core_1.execute.rf.reg_outputs[2][14] ),
    .A2(_2796_),
    .B1(_2804_),
    .C1(_2801_),
    .X(_0367_));
 sky130_fd_sc_hd__nand2_1 _6082_ (.A(_2695_),
    .B(_2786_),
    .Y(_2805_));
 sky130_fd_sc_hd__o211a_1 _6083_ (.A1(\core_1.execute.rf.reg_outputs[2][15] ),
    .A2(_2796_),
    .B1(_2805_),
    .C1(_2801_),
    .X(_0368_));
 sky130_fd_sc_hd__nand2_4 _6084_ (.A(\core_1.ew_reg_ie[1] ),
    .B(_2633_),
    .Y(_2806_));
 sky130_fd_sc_hd__and2_2 _6085_ (.A(\core_1.ew_reg_ie[1] ),
    .B(_2632_),
    .X(_2807_));
 sky130_fd_sc_hd__buf_4 _6086_ (.A(_2807_),
    .X(_2808_));
 sky130_fd_sc_hd__or2_1 _6087_ (.A(\core_1.execute.rf.reg_outputs[1][0] ),
    .B(_2808_),
    .X(_2809_));
 sky130_fd_sc_hd__o211a_1 _6088_ (.A1(_2637_),
    .A2(_2806_),
    .B1(_2809_),
    .C1(_2801_),
    .X(_0369_));
 sky130_fd_sc_hd__or2_1 _6089_ (.A(\core_1.execute.rf.reg_outputs[1][1] ),
    .B(_2808_),
    .X(_2810_));
 sky130_fd_sc_hd__o211a_1 _6090_ (.A1(_2643_),
    .A2(_2806_),
    .B1(_2810_),
    .C1(_2801_),
    .X(_0370_));
 sky130_fd_sc_hd__or2_1 _6091_ (.A(\core_1.execute.rf.reg_outputs[1][2] ),
    .B(_2808_),
    .X(_2811_));
 sky130_fd_sc_hd__o211a_1 _6092_ (.A1(_2648_),
    .A2(_2806_),
    .B1(_2811_),
    .C1(_2801_),
    .X(_0371_));
 sky130_fd_sc_hd__or2_1 _6093_ (.A(\core_1.execute.rf.reg_outputs[1][3] ),
    .B(_2808_),
    .X(_2812_));
 sky130_fd_sc_hd__o211a_1 _6094_ (.A1(_2652_),
    .A2(_2806_),
    .B1(_2812_),
    .C1(_2801_),
    .X(_0372_));
 sky130_fd_sc_hd__or2_1 _6095_ (.A(\core_1.execute.rf.reg_outputs[1][4] ),
    .B(_2807_),
    .X(_2813_));
 sky130_fd_sc_hd__o211a_1 _6096_ (.A1(_2656_),
    .A2(_2806_),
    .B1(_2813_),
    .C1(_2801_),
    .X(_0373_));
 sky130_fd_sc_hd__or2_1 _6097_ (.A(\core_1.execute.rf.reg_outputs[1][5] ),
    .B(_2807_),
    .X(_2814_));
 sky130_fd_sc_hd__clkbuf_4 _6098_ (.A(_2718_),
    .X(_2815_));
 sky130_fd_sc_hd__o211a_1 _6099_ (.A1(_2660_),
    .A2(_2806_),
    .B1(_2814_),
    .C1(_2815_),
    .X(_0374_));
 sky130_fd_sc_hd__or2_1 _6100_ (.A(\core_1.execute.rf.reg_outputs[1][6] ),
    .B(_2807_),
    .X(_2816_));
 sky130_fd_sc_hd__o211a_1 _6101_ (.A1(_2664_),
    .A2(_2806_),
    .B1(_2816_),
    .C1(_2815_),
    .X(_0375_));
 sky130_fd_sc_hd__or2_1 _6102_ (.A(\core_1.execute.rf.reg_outputs[1][7] ),
    .B(_2807_),
    .X(_2817_));
 sky130_fd_sc_hd__o211a_1 _6103_ (.A1(_2668_),
    .A2(_2806_),
    .B1(_2817_),
    .C1(_2815_),
    .X(_0376_));
 sky130_fd_sc_hd__buf_2 _6104_ (.A(_2807_),
    .X(_2818_));
 sky130_fd_sc_hd__nand2_1 _6105_ (.A(_2674_),
    .B(_2818_),
    .Y(_2819_));
 sky130_fd_sc_hd__o211a_1 _6106_ (.A1(\core_1.execute.rf.reg_outputs[1][8] ),
    .A2(_2818_),
    .B1(_2819_),
    .C1(_2815_),
    .X(_0377_));
 sky130_fd_sc_hd__nand2_1 _6107_ (.A(_2677_),
    .B(_2818_),
    .Y(_2820_));
 sky130_fd_sc_hd__o211a_1 _6108_ (.A1(\core_1.execute.rf.reg_outputs[1][9] ),
    .A2(_2818_),
    .B1(_2820_),
    .C1(_2815_),
    .X(_0378_));
 sky130_fd_sc_hd__nand2_1 _6109_ (.A(_2680_),
    .B(_2808_),
    .Y(_2821_));
 sky130_fd_sc_hd__o211a_1 _6110_ (.A1(\core_1.execute.rf.reg_outputs[1][10] ),
    .A2(_2818_),
    .B1(_2821_),
    .C1(_2815_),
    .X(_0379_));
 sky130_fd_sc_hd__nand2_1 _6111_ (.A(_2682_),
    .B(_2808_),
    .Y(_2822_));
 sky130_fd_sc_hd__o211a_1 _6112_ (.A1(\core_1.execute.rf.reg_outputs[1][11] ),
    .A2(_2818_),
    .B1(_2822_),
    .C1(_2815_),
    .X(_0380_));
 sky130_fd_sc_hd__nand2_1 _6113_ (.A(_2686_),
    .B(_2808_),
    .Y(_2823_));
 sky130_fd_sc_hd__o211a_1 _6114_ (.A1(\core_1.execute.rf.reg_outputs[1][12] ),
    .A2(_2818_),
    .B1(_2823_),
    .C1(_2815_),
    .X(_0381_));
 sky130_fd_sc_hd__nand2_1 _6115_ (.A(_2689_),
    .B(_2808_),
    .Y(_2824_));
 sky130_fd_sc_hd__o211a_1 _6116_ (.A1(\core_1.execute.rf.reg_outputs[1][13] ),
    .A2(_2818_),
    .B1(_2824_),
    .C1(_2815_),
    .X(_0382_));
 sky130_fd_sc_hd__nand2_1 _6117_ (.A(_2692_),
    .B(_2808_),
    .Y(_2825_));
 sky130_fd_sc_hd__o211a_1 _6118_ (.A1(\core_1.execute.rf.reg_outputs[1][14] ),
    .A2(_2818_),
    .B1(_2825_),
    .C1(_2815_),
    .X(_0383_));
 sky130_fd_sc_hd__nand2_1 _6119_ (.A(_2695_),
    .B(_2808_),
    .Y(_2826_));
 sky130_fd_sc_hd__clkbuf_4 _6120_ (.A(_2718_),
    .X(_2827_));
 sky130_fd_sc_hd__o211a_1 _6121_ (.A1(\core_1.execute.rf.reg_outputs[1][15] ),
    .A2(_2818_),
    .B1(_2826_),
    .C1(_2827_),
    .X(_0384_));
 sky130_fd_sc_hd__nand2_2 _6122_ (.A(\core_1.ew_reg_ie[0] ),
    .B(_2633_),
    .Y(_2828_));
 sky130_fd_sc_hd__and2_2 _6123_ (.A(\core_1.ew_reg_ie[0] ),
    .B(_2632_),
    .X(_2829_));
 sky130_fd_sc_hd__clkbuf_4 _6124_ (.A(_2829_),
    .X(_2830_));
 sky130_fd_sc_hd__or2_1 _6125_ (.A(net88),
    .B(_2830_),
    .X(_2831_));
 sky130_fd_sc_hd__o211a_1 _6126_ (.A1(_2637_),
    .A2(_2828_),
    .B1(_2831_),
    .C1(_2827_),
    .X(_0385_));
 sky130_fd_sc_hd__or2_1 _6127_ (.A(net95),
    .B(_2830_),
    .X(_2832_));
 sky130_fd_sc_hd__o211a_1 _6128_ (.A1(_2643_),
    .A2(_2828_),
    .B1(_2832_),
    .C1(_2827_),
    .X(_0386_));
 sky130_fd_sc_hd__or2_1 _6129_ (.A(net96),
    .B(_2830_),
    .X(_2833_));
 sky130_fd_sc_hd__o211a_1 _6130_ (.A1(_2648_),
    .A2(_2828_),
    .B1(_2833_),
    .C1(_2827_),
    .X(_0387_));
 sky130_fd_sc_hd__or2_1 _6131_ (.A(net97),
    .B(_2830_),
    .X(_2834_));
 sky130_fd_sc_hd__o211a_1 _6132_ (.A1(_2652_),
    .A2(_2828_),
    .B1(_2834_),
    .C1(_2827_),
    .X(_0388_));
 sky130_fd_sc_hd__or2_1 _6133_ (.A(net98),
    .B(_2829_),
    .X(_2835_));
 sky130_fd_sc_hd__o211a_1 _6134_ (.A1(_2656_),
    .A2(_2828_),
    .B1(_2835_),
    .C1(_2827_),
    .X(_0389_));
 sky130_fd_sc_hd__or2_1 _6135_ (.A(net99),
    .B(_2829_),
    .X(_2836_));
 sky130_fd_sc_hd__o211a_1 _6136_ (.A1(_2660_),
    .A2(_2828_),
    .B1(_2836_),
    .C1(_2827_),
    .X(_0390_));
 sky130_fd_sc_hd__or2_1 _6137_ (.A(net100),
    .B(_2829_),
    .X(_2837_));
 sky130_fd_sc_hd__o211a_1 _6138_ (.A1(_2664_),
    .A2(_2828_),
    .B1(_2837_),
    .C1(_2827_),
    .X(_0391_));
 sky130_fd_sc_hd__or2_1 _6139_ (.A(net101),
    .B(_2829_),
    .X(_2838_));
 sky130_fd_sc_hd__o211a_1 _6140_ (.A1(_2668_),
    .A2(_2828_),
    .B1(_2838_),
    .C1(_2827_),
    .X(_0392_));
 sky130_fd_sc_hd__buf_2 _6141_ (.A(_2829_),
    .X(_2839_));
 sky130_fd_sc_hd__nand2_1 _6142_ (.A(_2674_),
    .B(_2839_),
    .Y(_2840_));
 sky130_fd_sc_hd__o211a_1 _6143_ (.A1(net102),
    .A2(_2839_),
    .B1(_2840_),
    .C1(_2827_),
    .X(_0393_));
 sky130_fd_sc_hd__nand2_1 _6144_ (.A(_2677_),
    .B(_2839_),
    .Y(_2841_));
 sky130_fd_sc_hd__buf_6 _6145_ (.A(_2718_),
    .X(_2842_));
 sky130_fd_sc_hd__o211a_1 _6146_ (.A1(net103),
    .A2(_2839_),
    .B1(_2841_),
    .C1(_2842_),
    .X(_0394_));
 sky130_fd_sc_hd__nand2_1 _6147_ (.A(_2680_),
    .B(_2830_),
    .Y(_2843_));
 sky130_fd_sc_hd__o211a_1 _6148_ (.A1(net89),
    .A2(_2839_),
    .B1(_2843_),
    .C1(_2842_),
    .X(_0395_));
 sky130_fd_sc_hd__nand2_1 _6149_ (.A(_2682_),
    .B(_2830_),
    .Y(_2844_));
 sky130_fd_sc_hd__o211a_1 _6150_ (.A1(net90),
    .A2(_2839_),
    .B1(_2844_),
    .C1(_2842_),
    .X(_0396_));
 sky130_fd_sc_hd__nand2_1 _6151_ (.A(_2686_),
    .B(_2830_),
    .Y(_2845_));
 sky130_fd_sc_hd__o211a_1 _6152_ (.A1(net91),
    .A2(_2839_),
    .B1(_2845_),
    .C1(_2842_),
    .X(_0397_));
 sky130_fd_sc_hd__nand2_1 _6153_ (.A(_2689_),
    .B(_2830_),
    .Y(_2846_));
 sky130_fd_sc_hd__o211a_1 _6154_ (.A1(net92),
    .A2(_2839_),
    .B1(_2846_),
    .C1(_2842_),
    .X(_0398_));
 sky130_fd_sc_hd__nand2_1 _6155_ (.A(_2692_),
    .B(_2830_),
    .Y(_2847_));
 sky130_fd_sc_hd__o211a_1 _6156_ (.A1(net93),
    .A2(_2839_),
    .B1(_2847_),
    .C1(_2842_),
    .X(_0399_));
 sky130_fd_sc_hd__nand2_1 _6157_ (.A(_2695_),
    .B(_2830_),
    .Y(_2848_));
 sky130_fd_sc_hd__o211a_1 _6158_ (.A1(net94),
    .A2(_2839_),
    .B1(_2848_),
    .C1(_2842_),
    .X(_0400_));
 sky130_fd_sc_hd__a21oi_1 _6159_ (.A1(_1155_),
    .A2(_1029_),
    .B1(\core_1.execute.irq_en ),
    .Y(_2849_));
 sky130_fd_sc_hd__a21oi_1 _6160_ (.A1(_1163_),
    .A2(_2849_),
    .B1(_1168_),
    .Y(_2850_));
 sky130_fd_sc_hd__o31a_1 _6161_ (.A1(_1155_),
    .A2(net202),
    .A3(_1163_),
    .B1(_2850_),
    .X(_0401_));
 sky130_fd_sc_hd__and2_2 _6162_ (.A(\core_1.decode.o_submit ),
    .B(_0959_),
    .X(_2851_));
 sky130_fd_sc_hd__a21o_1 _6163_ (.A1(_1566_),
    .A2(_1428_),
    .B1(_2851_),
    .X(_2852_));
 sky130_fd_sc_hd__mux2_1 _6164_ (.A0(_2852_),
    .A1(_1203_),
    .S(_1806_),
    .X(_2853_));
 sky130_fd_sc_hd__clkbuf_1 _6165_ (.A(_2853_),
    .X(_0402_));
 sky130_fd_sc_hd__nand2_1 _6166_ (.A(_1808_),
    .B(_1317_),
    .Y(_2854_));
 sky130_fd_sc_hd__or2_4 _6167_ (.A(\core_1.execute.alu_mul_div.cbit[0] ),
    .B(\core_1.execute.alu_mul_div.cbit[1] ),
    .X(_2855_));
 sky130_fd_sc_hd__or2_1 _6168_ (.A(_2855_),
    .B(_1329_),
    .X(_2856_));
 sky130_fd_sc_hd__o221a_1 _6169_ (.A1(_1323_),
    .A2(_1636_),
    .B1(_1604_),
    .B2(_1699_),
    .C1(_2856_),
    .X(_2857_));
 sky130_fd_sc_hd__o22a_1 _6170_ (.A1(_2855_),
    .A2(_1361_),
    .B1(_1604_),
    .B2(_1696_),
    .X(_2858_));
 sky130_fd_sc_hd__a21oi_1 _6171_ (.A1(_1808_),
    .A2(_1349_),
    .B1(_1200_),
    .Y(_2859_));
 sky130_fd_sc_hd__o211a_1 _6172_ (.A1(_1351_),
    .A2(_1636_),
    .B1(_2858_),
    .C1(_2859_),
    .X(_2860_));
 sky130_fd_sc_hd__a311o_1 _6173_ (.A1(_1200_),
    .A2(_2854_),
    .A3(_2857_),
    .B1(_2860_),
    .C1(_1202_),
    .X(_2861_));
 sky130_fd_sc_hd__o22a_1 _6174_ (.A1(_1205_),
    .A2(_1689_),
    .B1(_2087_),
    .B2(_1636_),
    .X(_2862_));
 sky130_fd_sc_hd__o22a_1 _6175_ (.A1(_2855_),
    .A2(_1693_),
    .B1(_1604_),
    .B2(_1706_),
    .X(_2863_));
 sky130_fd_sc_hd__o22a_1 _6176_ (.A1(_1205_),
    .A2(_1866_),
    .B1(_1340_),
    .B2(_1636_),
    .X(_2864_));
 sky130_fd_sc_hd__o22a_1 _6177_ (.A1(_2855_),
    .A2(_1347_),
    .B1(_1604_),
    .B2(_1343_),
    .X(_2865_));
 sky130_fd_sc_hd__a31o_1 _6178_ (.A1(_1200_),
    .A2(_2864_),
    .A3(_2865_),
    .B1(_1810_),
    .X(_2866_));
 sky130_fd_sc_hd__a31o_1 _6179_ (.A1(_1608_),
    .A2(_2862_),
    .A3(_2863_),
    .B1(_2866_),
    .X(_2867_));
 sky130_fd_sc_hd__nand4_2 _6180_ (.A(_0959_),
    .B(\core_1.execute.alu_mul_div.comp ),
    .C(_2861_),
    .D(_2867_),
    .Y(_2868_));
 sky130_fd_sc_hd__and2_1 _6181_ (.A(_0734_),
    .B(_2868_),
    .X(_2869_));
 sky130_fd_sc_hd__buf_4 _6182_ (.A(_2869_),
    .X(_2870_));
 sky130_fd_sc_hd__clkbuf_4 _6183_ (.A(_2870_),
    .X(_2871_));
 sky130_fd_sc_hd__nor2_4 _6184_ (.A(_0734_),
    .B(_1419_),
    .Y(_2872_));
 sky130_fd_sc_hd__clkbuf_4 _6185_ (.A(_2872_),
    .X(_2873_));
 sky130_fd_sc_hd__nor2_1 _6186_ (.A(\core_1.decode.o_submit ),
    .B(_2868_),
    .Y(_2874_));
 sky130_fd_sc_hd__or2_1 _6187_ (.A(\core_1.execute.alu_mul_div.cbit[3] ),
    .B(\core_1.execute.alu_mul_div.cbit[2] ),
    .X(_2875_));
 sky130_fd_sc_hd__or4_1 _6188_ (.A(_2111_),
    .B(_2855_),
    .C(_1635_),
    .D(_2875_),
    .X(_2876_));
 sky130_fd_sc_hd__nor2_2 _6189_ (.A(_1570_),
    .B(_2855_),
    .Y(_2877_));
 sky130_fd_sc_hd__a31o_1 _6190_ (.A1(_1608_),
    .A2(_2877_),
    .A3(_1741_),
    .B1(\core_1.execute.alu_mul_div.mul_res[0] ),
    .X(_2878_));
 sky130_fd_sc_hd__and3_1 _6191_ (.A(_2874_),
    .B(_2876_),
    .C(_2878_),
    .X(_2879_));
 sky130_fd_sc_hd__a221o_1 _6192_ (.A1(\core_1.execute.alu_mul_div.mul_res[0] ),
    .A2(_2871_),
    .B1(_2873_),
    .B2(_1741_),
    .C1(_2879_),
    .X(_0403_));
 sky130_fd_sc_hd__o311a_1 _6193_ (.A1(_1630_),
    .A2(_1632_),
    .A3(_1633_),
    .B1(_1634_),
    .C1(\core_1.execute.alu_mul_div.cbit[0] ),
    .X(_2880_));
 sky130_fd_sc_hd__a31o_1 _6194_ (.A1(_1565_),
    .A2(_1618_),
    .A3(_1625_),
    .B1(_2880_),
    .X(_2881_));
 sky130_fd_sc_hd__and4_1 _6195_ (.A(_1201_),
    .B(_1602_),
    .C(\core_1.execute.alu_mul_div.mul_res[1] ),
    .D(_2881_),
    .X(_2882_));
 sky130_fd_sc_hd__a41oi_2 _6196_ (.A1(_1569_),
    .A2(_1201_),
    .A3(_1603_),
    .A4(_2881_),
    .B1(\core_1.execute.alu_mul_div.mul_res[1] ),
    .Y(_2883_));
 sky130_fd_sc_hd__a21o_1 _6197_ (.A1(_1608_),
    .A2(_2882_),
    .B1(_2883_),
    .X(_2884_));
 sky130_fd_sc_hd__a21oi_1 _6198_ (.A1(_2876_),
    .A2(_2884_),
    .B1(_2868_),
    .Y(_2885_));
 sky130_fd_sc_hd__clkbuf_4 _6199_ (.A(_0734_),
    .X(_2886_));
 sky130_fd_sc_hd__o211a_1 _6200_ (.A1(_2876_),
    .A2(_2884_),
    .B1(_2885_),
    .C1(_2886_),
    .X(_2887_));
 sky130_fd_sc_hd__a221o_1 _6201_ (.A1(\core_1.execute.alu_mul_div.mul_res[1] ),
    .A2(_2871_),
    .B1(_2873_),
    .B2(_1751_),
    .C1(_2887_),
    .X(_0404_));
 sky130_fd_sc_hd__inv_2 _6202_ (.A(\core_1.execute.alu_mul_div.mul_res[2] ),
    .Y(_2888_));
 sky130_fd_sc_hd__and4bb_1 _6203_ (.A_N(_2888_),
    .B_N(_1637_),
    .C(_1569_),
    .D(_1201_),
    .X(_2889_));
 sky130_fd_sc_hd__o31a_1 _6204_ (.A1(\core_1.execute.alu_mul_div.cbit[3] ),
    .A2(_1570_),
    .A3(_1637_),
    .B1(_2888_),
    .X(_2890_));
 sky130_fd_sc_hd__o2bb2a_1 _6205_ (.A1_N(_1569_),
    .A2_N(_2882_),
    .B1(_2883_),
    .B2(_2876_),
    .X(_2891_));
 sky130_fd_sc_hd__o21a_1 _6206_ (.A1(_2889_),
    .A2(_2890_),
    .B1(_2891_),
    .X(_2892_));
 sky130_fd_sc_hd__nor3_1 _6207_ (.A(_2889_),
    .B(_2890_),
    .C(_2891_),
    .Y(_2893_));
 sky130_fd_sc_hd__a21oi_1 _6208_ (.A1(_1974_),
    .A2(_2873_),
    .B1(_2870_),
    .Y(_2894_));
 sky130_fd_sc_hd__o31a_1 _6209_ (.A1(_2851_),
    .A2(_2892_),
    .A3(_2893_),
    .B1(_2894_),
    .X(_2895_));
 sky130_fd_sc_hd__a21oi_1 _6210_ (.A1(_2888_),
    .A2(_2871_),
    .B1(_2895_),
    .Y(_0405_));
 sky130_fd_sc_hd__inv_2 _6211_ (.A(\core_1.execute.alu_mul_div.mul_res[3] ),
    .Y(_2896_));
 sky130_fd_sc_hd__mux4_2 _6212_ (.A0(_1731_),
    .A1(_1635_),
    .A2(_1643_),
    .A3(_1727_),
    .S0(\core_1.execute.alu_mul_div.cbit[0] ),
    .S1(_1602_),
    .X(_2897_));
 sky130_fd_sc_hd__or4_1 _6213_ (.A(\core_1.execute.alu_mul_div.cbit[3] ),
    .B(\core_1.execute.alu_mul_div.cbit[2] ),
    .C(_2896_),
    .D(_2897_),
    .X(_2898_));
 sky130_fd_sc_hd__o31ai_1 _6214_ (.A1(_1199_),
    .A2(_1570_),
    .A3(_2897_),
    .B1(_2896_),
    .Y(_2899_));
 sky130_fd_sc_hd__nand2_1 _6215_ (.A(_2898_),
    .B(_2899_),
    .Y(_2900_));
 sky130_fd_sc_hd__o21bai_1 _6216_ (.A1(_2889_),
    .A2(_2893_),
    .B1_N(_2900_),
    .Y(_2901_));
 sky130_fd_sc_hd__or3b_1 _6217_ (.A(_2889_),
    .B(_2893_),
    .C_N(_2900_),
    .X(_2902_));
 sky130_fd_sc_hd__a32o_1 _6218_ (.A1(_2886_),
    .A2(_2901_),
    .A3(_2902_),
    .B1(_1723_),
    .B2(_2873_),
    .X(_2903_));
 sky130_fd_sc_hd__mux2_1 _6219_ (.A0(_2903_),
    .A1(\core_1.execute.alu_mul_div.mul_res[3] ),
    .S(_2871_),
    .X(_2904_));
 sky130_fd_sc_hd__clkbuf_1 _6220_ (.A(_2904_),
    .X(_0406_));
 sky130_fd_sc_hd__mux4_1 _6221_ (.A0(_1731_),
    .A1(_1727_),
    .A2(_1643_),
    .A3(_1650_),
    .S0(_1565_),
    .S1(_1602_),
    .X(_2905_));
 sky130_fd_sc_hd__nor2_1 _6222_ (.A(_2855_),
    .B(_1635_),
    .Y(_2906_));
 sky130_fd_sc_hd__nand2_1 _6223_ (.A(\core_1.execute.alu_mul_div.cbit[2] ),
    .B(_2906_),
    .Y(_2907_));
 sky130_fd_sc_hd__o21ai_2 _6224_ (.A1(_1570_),
    .A2(_2905_),
    .B1(_2907_),
    .Y(_2908_));
 sky130_fd_sc_hd__and3_1 _6225_ (.A(_1569_),
    .B(\core_1.execute.alu_mul_div.mul_res[4] ),
    .C(_2908_),
    .X(_2909_));
 sky130_fd_sc_hd__a21oi_1 _6226_ (.A1(_1569_),
    .A2(_2908_),
    .B1(\core_1.execute.alu_mul_div.mul_res[4] ),
    .Y(_2910_));
 sky130_fd_sc_hd__or2_1 _6227_ (.A(_2909_),
    .B(_2910_),
    .X(_2911_));
 sky130_fd_sc_hd__and3_1 _6228_ (.A(_2898_),
    .B(_2901_),
    .C(_2911_),
    .X(_2912_));
 sky130_fd_sc_hd__a21oi_1 _6229_ (.A1(_2898_),
    .A2(_2901_),
    .B1(_2911_),
    .Y(_2913_));
 sky130_fd_sc_hd__or3_1 _6230_ (.A(_2851_),
    .B(_2912_),
    .C(_2913_),
    .X(_2914_));
 sky130_fd_sc_hd__a21bo_1 _6231_ (.A1(_1724_),
    .A2(_2873_),
    .B1_N(_2914_),
    .X(_2915_));
 sky130_fd_sc_hd__mux2_1 _6232_ (.A0(_2915_),
    .A1(\core_1.execute.alu_mul_div.mul_res[4] ),
    .S(_2871_),
    .X(_2916_));
 sky130_fd_sc_hd__clkbuf_1 _6233_ (.A(_2916_),
    .X(_0407_));
 sky130_fd_sc_hd__nand2_1 _6234_ (.A(_1603_),
    .B(_2881_),
    .Y(_2917_));
 sky130_fd_sc_hd__mux4_1 _6235_ (.A0(_1974_),
    .A1(_1723_),
    .A2(_1724_),
    .A3(_1665_),
    .S0(_1565_),
    .S1(_1602_),
    .X(_2918_));
 sky130_fd_sc_hd__clkinv_2 _6236_ (.A(_2918_),
    .Y(_2919_));
 sky130_fd_sc_hd__mux2_1 _6237_ (.A0(_2917_),
    .A1(_2919_),
    .S(_1201_),
    .X(_2920_));
 sky130_fd_sc_hd__or3b_1 _6238_ (.A(_2920_),
    .B(_1199_),
    .C_N(\core_1.execute.alu_mul_div.mul_res[5] ),
    .X(_2921_));
 sky130_fd_sc_hd__o21bai_1 _6239_ (.A1(_1199_),
    .A2(_2920_),
    .B1_N(\core_1.execute.alu_mul_div.mul_res[5] ),
    .Y(_2922_));
 sky130_fd_sc_hd__o211ai_1 _6240_ (.A1(_2909_),
    .A2(_2913_),
    .B1(_2921_),
    .C1(_2922_),
    .Y(_2923_));
 sky130_fd_sc_hd__a211o_1 _6241_ (.A1(_2921_),
    .A2(_2922_),
    .B1(_2909_),
    .C1(_2913_),
    .X(_2924_));
 sky130_fd_sc_hd__and3_1 _6242_ (.A(_2874_),
    .B(_2923_),
    .C(_2924_),
    .X(_2925_));
 sky130_fd_sc_hd__a221o_1 _6243_ (.A1(\core_1.execute.alu_mul_div.mul_res[5] ),
    .A2(_2871_),
    .B1(_2873_),
    .B2(_1665_),
    .C1(_2925_),
    .X(_0408_));
 sky130_fd_sc_hd__nor2_1 _6244_ (.A(_1199_),
    .B(_1669_),
    .Y(_2926_));
 sky130_fd_sc_hd__xnor2_1 _6245_ (.A(\core_1.execute.alu_mul_div.mul_res[6] ),
    .B(_2926_),
    .Y(_2927_));
 sky130_fd_sc_hd__and3_1 _6246_ (.A(_2921_),
    .B(_2923_),
    .C(_2927_),
    .X(_2928_));
 sky130_fd_sc_hd__a21oi_1 _6247_ (.A1(_2921_),
    .A2(_2923_),
    .B1(_2927_),
    .Y(_2929_));
 sky130_fd_sc_hd__nor2_1 _6248_ (.A(_2928_),
    .B(_2929_),
    .Y(_2930_));
 sky130_fd_sc_hd__a22o_1 _6249_ (.A1(_1658_),
    .A2(_2872_),
    .B1(_2930_),
    .B2(_2886_),
    .X(_2931_));
 sky130_fd_sc_hd__mux2_1 _6250_ (.A0(_2931_),
    .A1(\core_1.execute.alu_mul_div.mul_res[6] ),
    .S(_2871_),
    .X(_2932_));
 sky130_fd_sc_hd__clkbuf_1 _6251_ (.A(_2932_),
    .X(_0409_));
 sky130_fd_sc_hd__and2_1 _6252_ (.A(\core_1.execute.alu_mul_div.mul_res[6] ),
    .B(_2926_),
    .X(_2933_));
 sky130_fd_sc_hd__clkinv_2 _6253_ (.A(_2897_),
    .Y(_2934_));
 sky130_fd_sc_hd__mux4_1 _6254_ (.A0(_1658_),
    .A1(_1724_),
    .A2(_1557_),
    .A3(_1665_),
    .S0(\core_1.execute.alu_mul_div.cbit[1] ),
    .S1(_1566_),
    .X(_2935_));
 sky130_fd_sc_hd__mux2_1 _6255_ (.A0(_2934_),
    .A1(_2935_),
    .S(_1202_),
    .X(_2936_));
 sky130_fd_sc_hd__and3_1 _6256_ (.A(_1608_),
    .B(\core_1.execute.alu_mul_div.mul_res[7] ),
    .C(_2936_),
    .X(_2937_));
 sky130_fd_sc_hd__a21oi_1 _6257_ (.A1(_1608_),
    .A2(_2936_),
    .B1(\core_1.execute.alu_mul_div.mul_res[7] ),
    .Y(_2938_));
 sky130_fd_sc_hd__or2_1 _6258_ (.A(_2937_),
    .B(_2938_),
    .X(_2939_));
 sky130_fd_sc_hd__o21ba_1 _6259_ (.A1(_2933_),
    .A2(_2929_),
    .B1_N(_2939_),
    .X(_2940_));
 sky130_fd_sc_hd__or3b_1 _6260_ (.A(_2933_),
    .B(_2929_),
    .C_N(_2939_),
    .X(_2941_));
 sky130_fd_sc_hd__nand2_1 _6261_ (.A(_2886_),
    .B(_2941_),
    .Y(_2942_));
 sky130_fd_sc_hd__a2bb2o_1 _6262_ (.A1_N(_2940_),
    .A2_N(_2942_),
    .B1(_1557_),
    .B2(_2872_),
    .X(_2943_));
 sky130_fd_sc_hd__mux2_1 _6263_ (.A0(_2943_),
    .A1(\core_1.execute.alu_mul_div.mul_res[7] ),
    .S(_2870_),
    .X(_2944_));
 sky130_fd_sc_hd__clkbuf_1 _6264_ (.A(_2944_),
    .X(_0410_));
 sky130_fd_sc_hd__mux2_1 _6265_ (.A0(_1666_),
    .A1(_1567_),
    .S(_1603_),
    .X(_2945_));
 sky130_fd_sc_hd__nor2_1 _6266_ (.A(_1571_),
    .B(_2905_),
    .Y(_2946_));
 sky130_fd_sc_hd__a31o_1 _6267_ (.A1(_1199_),
    .A2(_1202_),
    .A3(_2906_),
    .B1(_2946_),
    .X(_2947_));
 sky130_fd_sc_hd__a21o_1 _6268_ (.A1(_1607_),
    .A2(_2945_),
    .B1(_2947_),
    .X(_2948_));
 sky130_fd_sc_hd__and2_1 _6269_ (.A(\core_1.execute.alu_mul_div.mul_res[8] ),
    .B(_2948_),
    .X(_2949_));
 sky130_fd_sc_hd__nor2_1 _6270_ (.A(\core_1.execute.alu_mul_div.mul_res[8] ),
    .B(_2948_),
    .Y(_2950_));
 sky130_fd_sc_hd__nor2_1 _6271_ (.A(_2949_),
    .B(_2950_),
    .Y(_2951_));
 sky130_fd_sc_hd__o21a_1 _6272_ (.A1(_2937_),
    .A2(_2940_),
    .B1(_2951_),
    .X(_2952_));
 sky130_fd_sc_hd__o31ai_1 _6273_ (.A1(_2937_),
    .A2(_2940_),
    .A3(_2951_),
    .B1(_0734_),
    .Y(_2953_));
 sky130_fd_sc_hd__a2bb2o_1 _6274_ (.A1_N(_2952_),
    .A2_N(_2953_),
    .B1(_1564_),
    .B2(_2872_),
    .X(_2954_));
 sky130_fd_sc_hd__mux2_1 _6275_ (.A0(_2954_),
    .A1(\core_1.execute.alu_mul_div.mul_res[8] ),
    .S(_2870_),
    .X(_2955_));
 sky130_fd_sc_hd__clkbuf_1 _6276_ (.A(_2955_),
    .X(_0411_));
 sky130_fd_sc_hd__mux4_1 _6277_ (.A0(_1658_),
    .A1(_1557_),
    .A2(_1564_),
    .A3(_1535_),
    .S0(_1566_),
    .S1(_1603_),
    .X(_2956_));
 sky130_fd_sc_hd__a31o_1 _6278_ (.A1(_1202_),
    .A2(_1603_),
    .A3(_2881_),
    .B1(_1608_),
    .X(_2957_));
 sky130_fd_sc_hd__o221a_1 _6279_ (.A1(_1571_),
    .A2(_2918_),
    .B1(_2956_),
    .B2(_2875_),
    .C1(_2957_),
    .X(_2958_));
 sky130_fd_sc_hd__nand2_1 _6280_ (.A(\core_1.execute.alu_mul_div.mul_res[9] ),
    .B(_2958_),
    .Y(_2959_));
 sky130_fd_sc_hd__or2_1 _6281_ (.A(\core_1.execute.alu_mul_div.mul_res[9] ),
    .B(_2958_),
    .X(_2960_));
 sky130_fd_sc_hd__nand2_1 _6282_ (.A(_2959_),
    .B(_2960_),
    .Y(_2961_));
 sky130_fd_sc_hd__o21bai_1 _6283_ (.A1(_2949_),
    .A2(_2952_),
    .B1_N(_2961_),
    .Y(_2962_));
 sky130_fd_sc_hd__or3b_1 _6284_ (.A(_2949_),
    .B(_2952_),
    .C_N(_2961_),
    .X(_2963_));
 sky130_fd_sc_hd__a32o_1 _6285_ (.A1(_2886_),
    .A2(_2962_),
    .A3(_2963_),
    .B1(_1535_),
    .B2(_2873_),
    .X(_2964_));
 sky130_fd_sc_hd__mux2_1 _6286_ (.A0(_2964_),
    .A1(\core_1.execute.alu_mul_div.mul_res[9] ),
    .S(_2870_),
    .X(_2965_));
 sky130_fd_sc_hd__clkbuf_1 _6287_ (.A(_2965_),
    .X(_0412_));
 sky130_fd_sc_hd__inv_2 _6288_ (.A(\core_1.execute.alu_mul_div.mul_res[10] ),
    .Y(_2966_));
 sky130_fd_sc_hd__or2_1 _6289_ (.A(_1570_),
    .B(_1637_),
    .X(_2967_));
 sky130_fd_sc_hd__a21o_1 _6290_ (.A1(_1570_),
    .A2(_1668_),
    .B1(_1199_),
    .X(_2968_));
 sky130_fd_sc_hd__a2bb2o_1 _6291_ (.A1_N(_1568_),
    .A2_N(_2875_),
    .B1(_2967_),
    .B2(_2968_),
    .X(_2969_));
 sky130_fd_sc_hd__nor2_1 _6292_ (.A(_2966_),
    .B(_2969_),
    .Y(_2970_));
 sky130_fd_sc_hd__and2_1 _6293_ (.A(_2966_),
    .B(_2969_),
    .X(_2971_));
 sky130_fd_sc_hd__or2_1 _6294_ (.A(_2970_),
    .B(_2971_),
    .X(_2972_));
 sky130_fd_sc_hd__and3_1 _6295_ (.A(_2959_),
    .B(_2962_),
    .C(_2972_),
    .X(_2973_));
 sky130_fd_sc_hd__a21oi_1 _6296_ (.A1(_2959_),
    .A2(_2962_),
    .B1(_2972_),
    .Y(_2974_));
 sky130_fd_sc_hd__or3_1 _6297_ (.A(_2851_),
    .B(_2973_),
    .C(_2974_),
    .X(_2975_));
 sky130_fd_sc_hd__a21oi_1 _6298_ (.A1(_1543_),
    .A2(_2873_),
    .B1(_2871_),
    .Y(_2976_));
 sky130_fd_sc_hd__a22oi_1 _6299_ (.A1(_2966_),
    .A2(_2871_),
    .B1(_2975_),
    .B2(_2976_),
    .Y(_0413_));
 sky130_fd_sc_hd__or2_1 _6300_ (.A(_2970_),
    .B(_2974_),
    .X(_2977_));
 sky130_fd_sc_hd__o21ai_1 _6301_ (.A1(_1570_),
    .A2(_2897_),
    .B1(_1199_),
    .Y(_2978_));
 sky130_fd_sc_hd__or2_1 _6302_ (.A(_1571_),
    .B(_2935_),
    .X(_2979_));
 sky130_fd_sc_hd__mux2_1 _6303_ (.A0(_1535_),
    .A1(_1564_),
    .S(_1203_),
    .X(_2980_));
 sky130_fd_sc_hd__mux2_1 _6304_ (.A0(_1543_),
    .A1(_1586_),
    .S(_1566_),
    .X(_2981_));
 sky130_fd_sc_hd__mux2_1 _6305_ (.A0(_2980_),
    .A1(_2981_),
    .S(_1603_),
    .X(_2982_));
 sky130_fd_sc_hd__or2_1 _6306_ (.A(_2875_),
    .B(_2982_),
    .X(_2983_));
 sky130_fd_sc_hd__and4_1 _6307_ (.A(\core_1.execute.alu_mul_div.mul_res[11] ),
    .B(_2978_),
    .C(_2979_),
    .D(_2983_),
    .X(_2984_));
 sky130_fd_sc_hd__a31o_1 _6308_ (.A1(_2978_),
    .A2(_2979_),
    .A3(_2983_),
    .B1(\core_1.execute.alu_mul_div.mul_res[11] ),
    .X(_2985_));
 sky130_fd_sc_hd__or2b_1 _6309_ (.A(_2984_),
    .B_N(_2985_),
    .X(_2986_));
 sky130_fd_sc_hd__xnor2_1 _6310_ (.A(_2977_),
    .B(_2986_),
    .Y(_2987_));
 sky130_fd_sc_hd__nor2_1 _6311_ (.A(_2886_),
    .B(_2083_),
    .Y(_2988_));
 sky130_fd_sc_hd__a221o_1 _6312_ (.A1(\core_1.execute.alu_mul_div.mul_res[11] ),
    .A2(_2871_),
    .B1(_2874_),
    .B2(_2987_),
    .C1(_2988_),
    .X(_0414_));
 sky130_fd_sc_hd__nand2_1 _6313_ (.A(_1204_),
    .B(_1545_),
    .Y(_2989_));
 sky130_fd_sc_hd__o211a_1 _6314_ (.A1(_1204_),
    .A2(_1587_),
    .B1(_1607_),
    .C1(_2989_),
    .X(_2990_));
 sky130_fd_sc_hd__a221o_1 _6315_ (.A1(_1199_),
    .A2(_2908_),
    .B1(_2945_),
    .B2(_1572_),
    .C1(_2990_),
    .X(_2991_));
 sky130_fd_sc_hd__and2_1 _6316_ (.A(\core_1.execute.alu_mul_div.mul_res[12] ),
    .B(_2991_),
    .X(_2992_));
 sky130_fd_sc_hd__nor2_1 _6317_ (.A(\core_1.execute.alu_mul_div.mul_res[12] ),
    .B(_2991_),
    .Y(_2993_));
 sky130_fd_sc_hd__nor2_1 _6318_ (.A(_2992_),
    .B(_2993_),
    .Y(_2994_));
 sky130_fd_sc_hd__o311ai_2 _6319_ (.A1(_2970_),
    .A2(_2974_),
    .A3(_2984_),
    .B1(_2985_),
    .C1(_2994_),
    .Y(_2995_));
 sky130_fd_sc_hd__inv_2 _6320_ (.A(_2994_),
    .Y(_2996_));
 sky130_fd_sc_hd__o21ai_1 _6321_ (.A1(_2977_),
    .A2(_2984_),
    .B1(_2985_),
    .Y(_2997_));
 sky130_fd_sc_hd__nand2_1 _6322_ (.A(_2996_),
    .B(_2997_),
    .Y(_2998_));
 sky130_fd_sc_hd__a32o_1 _6323_ (.A1(_2886_),
    .A2(_2995_),
    .A3(_2998_),
    .B1(_1580_),
    .B2(_2873_),
    .X(_2999_));
 sky130_fd_sc_hd__mux2_1 _6324_ (.A0(_2999_),
    .A1(\core_1.execute.alu_mul_div.mul_res[12] ),
    .S(_2870_),
    .X(_3000_));
 sky130_fd_sc_hd__clkbuf_1 _6325_ (.A(_3000_),
    .X(_0415_));
 sky130_fd_sc_hd__nor2_1 _6326_ (.A(_2996_),
    .B(_2997_),
    .Y(_3001_));
 sky130_fd_sc_hd__nor2_1 _6327_ (.A(_1608_),
    .B(_2920_),
    .Y(_3002_));
 sky130_fd_sc_hd__mux2_1 _6328_ (.A0(_1580_),
    .A1(_1854_),
    .S(_1566_),
    .X(_3003_));
 sky130_fd_sc_hd__or2_1 _6329_ (.A(_1603_),
    .B(_2981_),
    .X(_3004_));
 sky130_fd_sc_hd__o211a_1 _6330_ (.A1(_1204_),
    .A2(_3003_),
    .B1(_3004_),
    .C1(_1607_),
    .X(_3005_));
 sky130_fd_sc_hd__a211o_1 _6331_ (.A1(_1572_),
    .A2(_2956_),
    .B1(_3002_),
    .C1(_3005_),
    .X(_3006_));
 sky130_fd_sc_hd__nand2_1 _6332_ (.A(\core_1.execute.alu_mul_div.mul_res[13] ),
    .B(_3006_),
    .Y(_3007_));
 sky130_fd_sc_hd__or2_1 _6333_ (.A(\core_1.execute.alu_mul_div.mul_res[13] ),
    .B(_3006_),
    .X(_3008_));
 sky130_fd_sc_hd__and2_1 _6334_ (.A(_3007_),
    .B(_3008_),
    .X(_3009_));
 sky130_fd_sc_hd__or3_1 _6335_ (.A(_2992_),
    .B(_3001_),
    .C(_3009_),
    .X(_3010_));
 sky130_fd_sc_hd__inv_2 _6336_ (.A(_2992_),
    .Y(_3011_));
 sky130_fd_sc_hd__a21bo_1 _6337_ (.A1(_3011_),
    .A2(_2995_),
    .B1_N(_3009_),
    .X(_3012_));
 sky130_fd_sc_hd__a32o_1 _6338_ (.A1(_2886_),
    .A2(_3010_),
    .A3(_3012_),
    .B1(_1854_),
    .B2(_2873_),
    .X(_3013_));
 sky130_fd_sc_hd__mux2_1 _6339_ (.A0(_3013_),
    .A1(\core_1.execute.alu_mul_div.mul_res[13] ),
    .S(_2870_),
    .X(_3014_));
 sky130_fd_sc_hd__clkbuf_1 _6340_ (.A(_3014_),
    .X(_0416_));
 sky130_fd_sc_hd__and2_1 _6341_ (.A(\core_1.execute.alu_mul_div.mul_res[14] ),
    .B(_1671_),
    .X(_3015_));
 sky130_fd_sc_hd__nor2_1 _6342_ (.A(\core_1.execute.alu_mul_div.mul_res[14] ),
    .B(_1671_),
    .Y(_3016_));
 sky130_fd_sc_hd__nor2_1 _6343_ (.A(_3015_),
    .B(_3016_),
    .Y(_3017_));
 sky130_fd_sc_hd__nand2_1 _6344_ (.A(_3007_),
    .B(_3012_),
    .Y(_3018_));
 sky130_fd_sc_hd__xor2_1 _6345_ (.A(_3017_),
    .B(_3018_),
    .X(_3019_));
 sky130_fd_sc_hd__a22o_1 _6346_ (.A1(_1594_),
    .A2(_2872_),
    .B1(_3019_),
    .B2(_2886_),
    .X(_3020_));
 sky130_fd_sc_hd__mux2_1 _6347_ (.A0(_3020_),
    .A1(\core_1.execute.alu_mul_div.mul_res[14] ),
    .S(_2870_),
    .X(_3021_));
 sky130_fd_sc_hd__clkbuf_1 _6348_ (.A(_3021_),
    .X(_0417_));
 sky130_fd_sc_hd__a21boi_1 _6349_ (.A1(_3007_),
    .A2(_3012_),
    .B1_N(_3017_),
    .Y(_3022_));
 sky130_fd_sc_hd__nor2_2 _6350_ (.A(_1566_),
    .B(_1204_),
    .Y(_3023_));
 sky130_fd_sc_hd__a22o_1 _6351_ (.A1(_3023_),
    .A2(_1594_),
    .B1(_3003_),
    .B2(_1204_),
    .X(_3024_));
 sky130_fd_sc_hd__a32o_1 _6352_ (.A1(_1608_),
    .A2(_2877_),
    .A3(_1529_),
    .B1(_1607_),
    .B2(_3024_),
    .X(_3025_));
 sky130_fd_sc_hd__a221o_1 _6353_ (.A1(_1200_),
    .A2(_2936_),
    .B1(_2982_),
    .B2(_1572_),
    .C1(_3025_),
    .X(_3026_));
 sky130_fd_sc_hd__xor2_1 _6354_ (.A(\core_1.execute.alu_mul_div.mul_res[15] ),
    .B(_3026_),
    .X(_3027_));
 sky130_fd_sc_hd__o21ai_1 _6355_ (.A1(_3015_),
    .A2(_3022_),
    .B1(_3027_),
    .Y(_3028_));
 sky130_fd_sc_hd__or3_1 _6356_ (.A(_3015_),
    .B(_3022_),
    .C(_3027_),
    .X(_3029_));
 sky130_fd_sc_hd__a32o_1 _6357_ (.A1(_2886_),
    .A2(_3028_),
    .A3(_3029_),
    .B1(_1529_),
    .B2(_2872_),
    .X(_3030_));
 sky130_fd_sc_hd__mux2_1 _6358_ (.A0(_3030_),
    .A1(\core_1.execute.alu_mul_div.mul_res[15] ),
    .S(_2870_),
    .X(_3031_));
 sky130_fd_sc_hd__clkbuf_1 _6359_ (.A(_3031_),
    .X(_0418_));
 sky130_fd_sc_hd__nor2_1 _6360_ (.A(_1128_),
    .B(_0731_),
    .Y(_0419_));
 sky130_fd_sc_hd__and2_1 _6361_ (.A(_1406_),
    .B(_1408_),
    .X(_3032_));
 sky130_fd_sc_hd__a21oi_1 _6362_ (.A1(_1416_),
    .A2(_3032_),
    .B1(\core_1.execute.alu_mul_div.div_res[0] ),
    .Y(_3033_));
 sky130_fd_sc_hd__nor2_1 _6363_ (.A(_1511_),
    .B(_3033_),
    .Y(_0420_));
 sky130_fd_sc_hd__nor2_2 _6364_ (.A(_1203_),
    .B(_1603_),
    .Y(_3034_));
 sky130_fd_sc_hd__nand2_1 _6365_ (.A(_1406_),
    .B(_1408_),
    .Y(_3035_));
 sky130_fd_sc_hd__nor2_2 _6366_ (.A(_1608_),
    .B(_3035_),
    .Y(_3036_));
 sky130_fd_sc_hd__a31o_1 _6367_ (.A1(_1810_),
    .A2(_3034_),
    .A3(_3036_),
    .B1(\core_1.execute.alu_mul_div.div_res[1] ),
    .X(_3037_));
 sky130_fd_sc_hd__and2_1 _6368_ (.A(_1477_),
    .B(_3037_),
    .X(_3038_));
 sky130_fd_sc_hd__clkbuf_1 _6369_ (.A(_3038_),
    .X(_0421_));
 sky130_fd_sc_hd__a31o_1 _6370_ (.A1(_1810_),
    .A2(_3023_),
    .A3(_3036_),
    .B1(\core_1.execute.alu_mul_div.div_res[2] ),
    .X(_3039_));
 sky130_fd_sc_hd__and2_1 _6371_ (.A(_1477_),
    .B(_3039_),
    .X(_3040_));
 sky130_fd_sc_hd__clkbuf_1 _6372_ (.A(_3040_),
    .X(_0422_));
 sky130_fd_sc_hd__a31o_1 _6373_ (.A1(_1810_),
    .A2(_1595_),
    .A3(_3036_),
    .B1(\core_1.execute.alu_mul_div.div_res[3] ),
    .X(_3041_));
 sky130_fd_sc_hd__and2_1 _6374_ (.A(_1477_),
    .B(_3041_),
    .X(_3042_));
 sky130_fd_sc_hd__clkbuf_1 _6375_ (.A(_3042_),
    .X(_0423_));
 sky130_fd_sc_hd__nor2_1 _6376_ (.A(_1810_),
    .B(_1205_),
    .Y(_3043_));
 sky130_fd_sc_hd__a21oi_1 _6377_ (.A1(_3036_),
    .A2(_3043_),
    .B1(\core_1.execute.alu_mul_div.div_res[4] ),
    .Y(_3044_));
 sky130_fd_sc_hd__nor2_1 _6378_ (.A(_1511_),
    .B(_3044_),
    .Y(_0424_));
 sky130_fd_sc_hd__a31o_1 _6379_ (.A1(_1202_),
    .A2(_3034_),
    .A3(_3036_),
    .B1(\core_1.execute.alu_mul_div.div_res[5] ),
    .X(_3045_));
 sky130_fd_sc_hd__and2_1 _6380_ (.A(_1428_),
    .B(_3045_),
    .X(_3046_));
 sky130_fd_sc_hd__clkbuf_1 _6381_ (.A(_3046_),
    .X(_0425_));
 sky130_fd_sc_hd__and3_1 _6382_ (.A(_1202_),
    .B(_3023_),
    .C(_3036_),
    .X(_3047_));
 sky130_fd_sc_hd__o21a_1 _6383_ (.A1(\core_1.execute.alu_mul_div.div_res[6] ),
    .A2(_3047_),
    .B1(_1429_),
    .X(_0426_));
 sky130_fd_sc_hd__a31o_1 _6384_ (.A1(_1200_),
    .A2(_2877_),
    .A3(_3032_),
    .B1(\core_1.execute.alu_mul_div.div_res[7] ),
    .X(_3048_));
 sky130_fd_sc_hd__and2_1 _6385_ (.A(_1428_),
    .B(_3048_),
    .X(_3049_));
 sky130_fd_sc_hd__clkbuf_1 _6386_ (.A(_3049_),
    .X(_0427_));
 sky130_fd_sc_hd__nor2_2 _6387_ (.A(_1200_),
    .B(_3035_),
    .Y(_3050_));
 sky130_fd_sc_hd__a21oi_1 _6388_ (.A1(_1206_),
    .A2(_3050_),
    .B1(\core_1.execute.alu_mul_div.div_res[8] ),
    .Y(_3051_));
 sky130_fd_sc_hd__nor2_1 _6389_ (.A(_1511_),
    .B(_3051_),
    .Y(_0428_));
 sky130_fd_sc_hd__a31o_1 _6390_ (.A1(_1810_),
    .A2(_3034_),
    .A3(_3050_),
    .B1(\core_1.execute.alu_mul_div.div_res[9] ),
    .X(_3052_));
 sky130_fd_sc_hd__and2_1 _6391_ (.A(_1428_),
    .B(_3052_),
    .X(_3053_));
 sky130_fd_sc_hd__clkbuf_1 _6392_ (.A(_3053_),
    .X(_0429_));
 sky130_fd_sc_hd__a31o_1 _6393_ (.A1(_1810_),
    .A2(_3023_),
    .A3(_3050_),
    .B1(\core_1.execute.alu_mul_div.div_res[10] ),
    .X(_3054_));
 sky130_fd_sc_hd__and2_1 _6394_ (.A(_1428_),
    .B(_3054_),
    .X(_3055_));
 sky130_fd_sc_hd__clkbuf_1 _6395_ (.A(_3055_),
    .X(_0430_));
 sky130_fd_sc_hd__a31o_1 _6396_ (.A1(_1810_),
    .A2(_1595_),
    .A3(_3050_),
    .B1(\core_1.execute.alu_mul_div.div_res[11] ),
    .X(_3056_));
 sky130_fd_sc_hd__and2_1 _6397_ (.A(_1428_),
    .B(_3056_),
    .X(_3057_));
 sky130_fd_sc_hd__clkbuf_1 _6398_ (.A(_3057_),
    .X(_0431_));
 sky130_fd_sc_hd__a21oi_1 _6399_ (.A1(_3043_),
    .A2(_3050_),
    .B1(\core_1.execute.alu_mul_div.div_res[12] ),
    .Y(_3058_));
 sky130_fd_sc_hd__nor2_1 _6400_ (.A(_1511_),
    .B(_3058_),
    .Y(_0432_));
 sky130_fd_sc_hd__a31o_1 _6401_ (.A1(_1202_),
    .A2(_3034_),
    .A3(_3050_),
    .B1(\core_1.execute.alu_mul_div.div_res[13] ),
    .X(_3059_));
 sky130_fd_sc_hd__and2_1 _6402_ (.A(_1428_),
    .B(_3059_),
    .X(_3060_));
 sky130_fd_sc_hd__clkbuf_1 _6403_ (.A(_3060_),
    .X(_0433_));
 sky130_fd_sc_hd__and3_1 _6404_ (.A(_1202_),
    .B(_3023_),
    .C(_3050_),
    .X(_3061_));
 sky130_fd_sc_hd__o21a_1 _6405_ (.A1(\core_1.execute.alu_mul_div.div_res[14] ),
    .A2(_3061_),
    .B1(_1429_),
    .X(_0434_));
 sky130_fd_sc_hd__a21oi_1 _6406_ (.A1(_2877_),
    .A2(_3050_),
    .B1(\core_1.execute.alu_mul_div.div_res[15] ),
    .Y(_3062_));
 sky130_fd_sc_hd__nor2_1 _6407_ (.A(_1511_),
    .B(_3062_),
    .Y(_0435_));
 sky130_fd_sc_hd__clkbuf_4 _6408_ (.A(_1678_),
    .X(_3063_));
 sky130_fd_sc_hd__buf_2 _6409_ (.A(_3063_),
    .X(_3064_));
 sky130_fd_sc_hd__nand2_4 _6410_ (.A(_1799_),
    .B(_1153_),
    .Y(_3065_));
 sky130_fd_sc_hd__or2_2 _6411_ (.A(_1057_),
    .B(_1153_),
    .X(_3066_));
 sky130_fd_sc_hd__o221a_1 _6412_ (.A1(net194),
    .A2(_3065_),
    .B1(_2114_),
    .B2(_3066_),
    .C1(_2053_),
    .X(_3067_));
 sky130_fd_sc_hd__xnor2_1 _6413_ (.A(net211),
    .B(_1681_),
    .Y(_3068_));
 sky130_fd_sc_hd__nand2_1 _6414_ (.A(_3064_),
    .B(_3068_),
    .Y(_3069_));
 sky130_fd_sc_hd__nor2_8 _6415_ (.A(net71),
    .B(_0670_),
    .Y(_3070_));
 sky130_fd_sc_hd__clkbuf_4 _6416_ (.A(_3070_),
    .X(_3071_));
 sky130_fd_sc_hd__o211a_1 _6417_ (.A1(_3064_),
    .A2(_3067_),
    .B1(_3069_),
    .C1(_3071_),
    .X(_0436_));
 sky130_fd_sc_hd__a31o_1 _6418_ (.A1(net211),
    .A2(net79),
    .A3(_1681_),
    .B1(net80),
    .X(_3072_));
 sky130_fd_sc_hd__and3_1 _6419_ (.A(net80),
    .B(net211),
    .C(net79),
    .X(_3073_));
 sky130_fd_sc_hd__nand2_1 _6420_ (.A(_1681_),
    .B(_3073_),
    .Y(_3074_));
 sky130_fd_sc_hd__and3_1 _6421_ (.A(_1679_),
    .B(_3072_),
    .C(_3074_),
    .X(_3075_));
 sky130_fd_sc_hd__inv_2 _6422_ (.A(\core_1.execute.sreg_irq_pc.o_d[2] ),
    .Y(_3076_));
 sky130_fd_sc_hd__a221o_1 _6423_ (.A1(_3076_),
    .A2(_1155_),
    .B1(_0647_),
    .B2(_1801_),
    .C1(_1678_),
    .X(_3077_));
 sky130_fd_sc_hd__o21ba_1 _6424_ (.A1(_3066_),
    .A2(_2182_),
    .B1_N(_3077_),
    .X(_3078_));
 sky130_fd_sc_hd__o21a_1 _6425_ (.A1(_3075_),
    .A2(_3078_),
    .B1(_3071_),
    .X(_0437_));
 sky130_fd_sc_hd__and2_1 _6426_ (.A(_1824_),
    .B(_3074_),
    .X(_3079_));
 sky130_fd_sc_hd__nor2_1 _6427_ (.A(_1824_),
    .B(_3074_),
    .Y(_3080_));
 sky130_fd_sc_hd__o21ai_1 _6428_ (.A1(_3079_),
    .A2(_3080_),
    .B1(_1679_),
    .Y(_3081_));
 sky130_fd_sc_hd__clkbuf_4 _6429_ (.A(_1684_),
    .X(_3082_));
 sky130_fd_sc_hd__a22o_1 _6430_ (.A1(\core_1.execute.sreg_irq_pc.o_d[3] ),
    .A2(_1155_),
    .B1(net203),
    .B2(_1801_),
    .X(_3083_));
 sky130_fd_sc_hd__a211o_1 _6431_ (.A1(_3082_),
    .A2(_2219_),
    .B1(_3083_),
    .C1(_3063_),
    .X(_3084_));
 sky130_fd_sc_hd__and3_1 _6432_ (.A(_3070_),
    .B(_3081_),
    .C(_3084_),
    .X(_3085_));
 sky130_fd_sc_hd__clkbuf_1 _6433_ (.A(_3085_),
    .X(_0438_));
 sky130_fd_sc_hd__nor2_1 _6434_ (.A(_3066_),
    .B(_2245_),
    .Y(_3086_));
 sky130_fd_sc_hd__a221o_1 _6435_ (.A1(\core_1.execute.sreg_irq_pc.o_d[4] ),
    .A2(_1155_),
    .B1(net204),
    .B2(_1801_),
    .C1(_1679_),
    .X(_3087_));
 sky130_fd_sc_hd__o21ai_1 _6436_ (.A1(_1827_),
    .A2(_3080_),
    .B1(_1679_),
    .Y(_3088_));
 sky130_fd_sc_hd__a21o_1 _6437_ (.A1(_1827_),
    .A2(_3080_),
    .B1(_3088_),
    .X(_3089_));
 sky130_fd_sc_hd__o211a_1 _6438_ (.A1(_3086_),
    .A2(_3087_),
    .B1(_3089_),
    .C1(_3071_),
    .X(_0439_));
 sky130_fd_sc_hd__nor2_1 _6439_ (.A(_0627_),
    .B(_3065_),
    .Y(_3090_));
 sky130_fd_sc_hd__a221o_1 _6440_ (.A1(\core_1.execute.sreg_irq_pc.o_d[5] ),
    .A2(_1155_),
    .B1(_3082_),
    .B2(_2292_),
    .C1(_3090_),
    .X(_3091_));
 sky130_fd_sc_hd__and3_1 _6441_ (.A(net82),
    .B(net81),
    .C(_3073_),
    .X(_3092_));
 sky130_fd_sc_hd__a21oi_1 _6442_ (.A1(_1681_),
    .A2(_3092_),
    .B1(net83),
    .Y(_3093_));
 sky130_fd_sc_hd__and3_1 _6443_ (.A(net83),
    .B(net82),
    .C(_3080_),
    .X(_3094_));
 sky130_fd_sc_hd__o21ai_1 _6444_ (.A1(_3093_),
    .A2(_3094_),
    .B1(_3064_),
    .Y(_3095_));
 sky130_fd_sc_hd__o211a_1 _6445_ (.A1(_3064_),
    .A2(_3091_),
    .B1(_3095_),
    .C1(_3071_),
    .X(_0440_));
 sky130_fd_sc_hd__nor2_1 _6446_ (.A(_0621_),
    .B(_3065_),
    .Y(_3096_));
 sky130_fd_sc_hd__a221o_1 _6447_ (.A1(\core_1.execute.sreg_irq_pc.o_d[6] ),
    .A2(_1155_),
    .B1(_3082_),
    .B2(_2326_),
    .C1(_3096_),
    .X(_3097_));
 sky130_fd_sc_hd__xnor2_1 _6448_ (.A(net84),
    .B(_3094_),
    .Y(_3098_));
 sky130_fd_sc_hd__nand2_1 _6449_ (.A(_3064_),
    .B(_3098_),
    .Y(_3099_));
 sky130_fd_sc_hd__o211a_1 _6450_ (.A1(_3064_),
    .A2(_3097_),
    .B1(_3099_),
    .C1(_3071_),
    .X(_0441_));
 sky130_fd_sc_hd__a221o_1 _6451_ (.A1(net207),
    .A2(_1801_),
    .B1(_2363_),
    .B2(_3082_),
    .C1(_2337_),
    .X(_3100_));
 sky130_fd_sc_hd__a21oi_1 _6452_ (.A1(net84),
    .A2(_3094_),
    .B1(net85),
    .Y(_3101_));
 sky130_fd_sc_hd__and3_1 _6453_ (.A(net85),
    .B(net84),
    .C(_3094_),
    .X(_3102_));
 sky130_fd_sc_hd__o21ai_1 _6454_ (.A1(_3101_),
    .A2(_3102_),
    .B1(_1679_),
    .Y(_3103_));
 sky130_fd_sc_hd__o211a_1 _6455_ (.A1(_3064_),
    .A2(_3100_),
    .B1(_3103_),
    .C1(_3071_),
    .X(_0442_));
 sky130_fd_sc_hd__nor2_1 _6456_ (.A(net86),
    .B(_3102_),
    .Y(_3104_));
 sky130_fd_sc_hd__and2_1 _6457_ (.A(net86),
    .B(_3102_),
    .X(_3105_));
 sky130_fd_sc_hd__o21ai_1 _6458_ (.A1(_3104_),
    .A2(_3105_),
    .B1(_1679_),
    .Y(_3106_));
 sky130_fd_sc_hd__a22o_1 _6459_ (.A1(\core_1.execute.sreg_irq_pc.o_d[8] ),
    .A2(_1155_),
    .B1(net208),
    .B2(_1801_),
    .X(_3107_));
 sky130_fd_sc_hd__a211o_1 _6460_ (.A1(_3082_),
    .A2(_2383_),
    .B1(_3107_),
    .C1(_3063_),
    .X(_3108_));
 sky130_fd_sc_hd__and3_1 _6461_ (.A(_3070_),
    .B(_3106_),
    .C(_3108_),
    .X(_3109_));
 sky130_fd_sc_hd__clkbuf_1 _6462_ (.A(_3109_),
    .X(_0443_));
 sky130_fd_sc_hd__xnor2_1 _6463_ (.A(net87),
    .B(_3105_),
    .Y(_3110_));
 sky130_fd_sc_hd__nand2_1 _6464_ (.A(_1679_),
    .B(_3110_),
    .Y(_3111_));
 sky130_fd_sc_hd__o21ai_1 _6465_ (.A1(_0600_),
    .A2(_3065_),
    .B1(_2398_),
    .Y(_3112_));
 sky130_fd_sc_hd__a211o_1 _6466_ (.A1(_3082_),
    .A2(_2423_),
    .B1(_3112_),
    .C1(_3063_),
    .X(_3113_));
 sky130_fd_sc_hd__and3_1 _6467_ (.A(_3070_),
    .B(_3111_),
    .C(_3113_),
    .X(_3114_));
 sky130_fd_sc_hd__clkbuf_1 _6468_ (.A(_3114_),
    .X(_0444_));
 sky130_fd_sc_hd__a21oi_1 _6469_ (.A1(net87),
    .A2(_3105_),
    .B1(net73),
    .Y(_3115_));
 sky130_fd_sc_hd__and3_1 _6470_ (.A(net73),
    .B(net87),
    .C(_3105_),
    .X(_3116_));
 sky130_fd_sc_hd__o21ai_1 _6471_ (.A1(_3115_),
    .A2(_3116_),
    .B1(_1679_),
    .Y(_3117_));
 sky130_fd_sc_hd__a21o_1 _6472_ (.A1(net195),
    .A2(_1801_),
    .B1(_2431_),
    .X(_3118_));
 sky130_fd_sc_hd__a211o_1 _6473_ (.A1(_3082_),
    .A2(_2454_),
    .B1(_3118_),
    .C1(_3063_),
    .X(_3119_));
 sky130_fd_sc_hd__and3_1 _6474_ (.A(_3070_),
    .B(_3117_),
    .C(_3119_),
    .X(_3120_));
 sky130_fd_sc_hd__clkbuf_1 _6475_ (.A(_3120_),
    .X(_0445_));
 sky130_fd_sc_hd__or2_1 _6476_ (.A(net74),
    .B(_3116_),
    .X(_3121_));
 sky130_fd_sc_hd__nand2_1 _6477_ (.A(net74),
    .B(_3116_),
    .Y(_3122_));
 sky130_fd_sc_hd__a21bo_1 _6478_ (.A1(_3121_),
    .A2(_3122_),
    .B1_N(_3063_),
    .X(_3123_));
 sky130_fd_sc_hd__a22o_1 _6479_ (.A1(\core_1.execute.sreg_irq_pc.o_d[11] ),
    .A2(_1155_),
    .B1(net196),
    .B2(_1801_),
    .X(_3124_));
 sky130_fd_sc_hd__a211o_1 _6480_ (.A1(_3082_),
    .A2(_2479_),
    .B1(_3124_),
    .C1(_3063_),
    .X(_3125_));
 sky130_fd_sc_hd__and3_1 _6481_ (.A(_3070_),
    .B(_3123_),
    .C(_3125_),
    .X(_3126_));
 sky130_fd_sc_hd__clkbuf_1 _6482_ (.A(_3126_),
    .X(_0446_));
 sky130_fd_sc_hd__o221ai_1 _6483_ (.A1(_0577_),
    .A2(_3065_),
    .B1(_2512_),
    .B2(_3066_),
    .C1(_2492_),
    .Y(_3127_));
 sky130_fd_sc_hd__o21ai_1 _6484_ (.A1(net75),
    .A2(_3122_),
    .B1(_3063_),
    .Y(_3128_));
 sky130_fd_sc_hd__a21o_1 _6485_ (.A1(net75),
    .A2(_3122_),
    .B1(_3128_),
    .X(_3129_));
 sky130_fd_sc_hd__o211a_1 _6486_ (.A1(_3064_),
    .A2(_3127_),
    .B1(_3129_),
    .C1(_3071_),
    .X(_0447_));
 sky130_fd_sc_hd__a221o_1 _6487_ (.A1(net198),
    .A2(_1801_),
    .B1(_2542_),
    .B2(_3082_),
    .C1(_2521_),
    .X(_3130_));
 sky130_fd_sc_hd__and3_1 _6488_ (.A(net86),
    .B(net85),
    .C(net84),
    .X(_3131_));
 sky130_fd_sc_hd__and4_1 _6489_ (.A(net75),
    .B(net74),
    .C(net73),
    .D(net87),
    .X(_3132_));
 sky130_fd_sc_hd__and3_1 _6490_ (.A(net83),
    .B(_3131_),
    .C(_3132_),
    .X(_3133_));
 sky130_fd_sc_hd__and3_1 _6491_ (.A(_1681_),
    .B(_3092_),
    .C(_3133_),
    .X(_3134_));
 sky130_fd_sc_hd__xnor2_1 _6492_ (.A(net76),
    .B(_3134_),
    .Y(_3135_));
 sky130_fd_sc_hd__nand2_1 _6493_ (.A(_3064_),
    .B(_3135_),
    .Y(_3136_));
 sky130_fd_sc_hd__o211a_1 _6494_ (.A1(_3064_),
    .A2(_3130_),
    .B1(_3136_),
    .C1(_3071_),
    .X(_0448_));
 sky130_fd_sc_hd__o221a_1 _6495_ (.A1(_0556_),
    .A2(_3065_),
    .B1(_2570_),
    .B2(_3066_),
    .C1(_2550_),
    .X(_3137_));
 sky130_fd_sc_hd__and4_1 _6496_ (.A(net83),
    .B(_3092_),
    .C(_3131_),
    .D(_3132_),
    .X(_3138_));
 sky130_fd_sc_hd__and3_1 _6497_ (.A(net76),
    .B(_1681_),
    .C(_3138_),
    .X(_3139_));
 sky130_fd_sc_hd__or2_1 _6498_ (.A(net77),
    .B(_3139_),
    .X(_3140_));
 sky130_fd_sc_hd__nand2_1 _6499_ (.A(net77),
    .B(_3139_),
    .Y(_3141_));
 sky130_fd_sc_hd__nand2_1 _6500_ (.A(_3140_),
    .B(_3141_),
    .Y(_3142_));
 sky130_fd_sc_hd__mux2_1 _6501_ (.A0(_3137_),
    .A1(_3142_),
    .S(_3063_),
    .X(_3143_));
 sky130_fd_sc_hd__nor2_1 _6502_ (.A(_1168_),
    .B(_3143_),
    .Y(_0449_));
 sky130_fd_sc_hd__xor2_1 _6503_ (.A(net78),
    .B(_3141_),
    .X(_3144_));
 sky130_fd_sc_hd__nand2_1 _6504_ (.A(_1679_),
    .B(_3144_),
    .Y(_3145_));
 sky130_fd_sc_hd__a22o_1 _6505_ (.A1(\core_1.execute.sreg_irq_pc.o_d[15] ),
    .A2(_1057_),
    .B1(net200),
    .B2(_1801_),
    .X(_3146_));
 sky130_fd_sc_hd__a211o_1 _6506_ (.A1(_3082_),
    .A2(_2600_),
    .B1(_3146_),
    .C1(_3063_),
    .X(_3147_));
 sky130_fd_sc_hd__and3_1 _6507_ (.A(_3070_),
    .B(_3145_),
    .C(_3147_),
    .X(_3148_));
 sky130_fd_sc_hd__clkbuf_1 _6508_ (.A(_3148_),
    .X(_0450_));
 sky130_fd_sc_hd__and3_1 _6509_ (.A(\core_1.dec_sreg_store ),
    .B(_1056_),
    .C(_2066_),
    .X(_3149_));
 sky130_fd_sc_hd__clkbuf_4 _6510_ (.A(_3149_),
    .X(_3150_));
 sky130_fd_sc_hd__o21a_2 _6511_ (.A1(\core_1.dec_alu_flags_ie ),
    .A2(_3150_),
    .B1(_1029_),
    .X(_3151_));
 sky130_fd_sc_hd__nand2_1 _6512_ (.A(_2380_),
    .B(_2420_),
    .Y(_3152_));
 sky130_fd_sc_hd__or2_1 _6513_ (.A(_2323_),
    .B(_2360_),
    .X(_3153_));
 sky130_fd_sc_hd__or2_1 _6514_ (.A(_2242_),
    .B(_2289_),
    .X(_3154_));
 sky130_fd_sc_hd__nand2_1 _6515_ (.A(_1794_),
    .B(_2110_),
    .Y(_3155_));
 sky130_fd_sc_hd__or4bb_1 _6516_ (.A(_3150_),
    .B(_3155_),
    .C_N(_2179_),
    .D_N(_2216_),
    .X(_3156_));
 sky130_fd_sc_hd__or4_1 _6517_ (.A(_3152_),
    .B(_3153_),
    .C(_3154_),
    .D(_3156_),
    .X(_3157_));
 sky130_fd_sc_hd__and4b_1 _6518_ (.A_N(_2451_),
    .B(_2476_),
    .C(_2509_),
    .D(_2539_),
    .X(_3158_));
 sky130_fd_sc_hd__or4b_1 _6519_ (.A(_2566_),
    .B(_2596_),
    .C(_3157_),
    .D_N(_3158_),
    .X(_3159_));
 sky130_fd_sc_hd__nand2_1 _6520_ (.A(net194),
    .B(_3150_),
    .Y(_3160_));
 sky130_fd_sc_hd__nand3_1 _6521_ (.A(_3159_),
    .B(_3160_),
    .C(_3151_),
    .Y(_3161_));
 sky130_fd_sc_hd__o211a_1 _6522_ (.A1(\core_1.execute.alu_flag_reg.o_d[0] ),
    .A2(_3151_),
    .B1(_3161_),
    .C1(_2842_),
    .X(_0451_));
 sky130_fd_sc_hd__mux2_1 _6523_ (.A0(_2005_),
    .A1(net201),
    .S(_3150_),
    .X(_3162_));
 sky130_fd_sc_hd__mux2_1 _6524_ (.A0(\core_1.execute.alu_flag_reg.o_d[1] ),
    .A1(_3162_),
    .S(_3151_),
    .X(_3163_));
 sky130_fd_sc_hd__and2_1 _6525_ (.A(_1184_),
    .B(_3163_),
    .X(_3164_));
 sky130_fd_sc_hd__clkbuf_1 _6526_ (.A(_3164_),
    .X(_0452_));
 sky130_fd_sc_hd__mux2_1 _6527_ (.A0(_2596_),
    .A1(net202),
    .S(_3150_),
    .X(_3165_));
 sky130_fd_sc_hd__mux2_1 _6528_ (.A0(\core_1.execute.alu_flag_reg.o_d[2] ),
    .A1(_3165_),
    .S(_3151_),
    .X(_3166_));
 sky130_fd_sc_hd__and2_1 _6529_ (.A(_1184_),
    .B(_3166_),
    .X(_3167_));
 sky130_fd_sc_hd__clkbuf_1 _6530_ (.A(_3167_),
    .X(_0453_));
 sky130_fd_sc_hd__nor2_1 _6531_ (.A(_0981_),
    .B(_1852_),
    .Y(_3168_));
 sky130_fd_sc_hd__a21o_1 _6532_ (.A1(_0981_),
    .A2(_1852_),
    .B1(_3150_),
    .X(_3169_));
 sky130_fd_sc_hd__mux2_1 _6533_ (.A0(_2595_),
    .A1(_2596_),
    .S(_1529_),
    .X(_3170_));
 sky130_fd_sc_hd__or3_1 _6534_ (.A(_3168_),
    .B(_3169_),
    .C(_3170_),
    .X(_3171_));
 sky130_fd_sc_hd__nand2_1 _6535_ (.A(net203),
    .B(_3150_),
    .Y(_3172_));
 sky130_fd_sc_hd__a31o_1 _6536_ (.A1(_3151_),
    .A2(_3171_),
    .A3(_3172_),
    .B1(_1121_),
    .X(_3173_));
 sky130_fd_sc_hd__o21ba_1 _6537_ (.A1(\core_1.execute.alu_flag_reg.o_d[3] ),
    .A2(_3151_),
    .B1_N(_3173_),
    .X(_0454_));
 sky130_fd_sc_hd__nor2_1 _6538_ (.A(\core_1.execute.alu_flag_reg.o_d[4] ),
    .B(_3151_),
    .Y(_3174_));
 sky130_fd_sc_hd__xnor2_1 _6539_ (.A(_2179_),
    .B(_2216_),
    .Y(_3175_));
 sky130_fd_sc_hd__xor2_1 _6540_ (.A(_2242_),
    .B(_2289_),
    .X(_3176_));
 sky130_fd_sc_hd__or2_1 _6541_ (.A(_1794_),
    .B(_2110_),
    .X(_3177_));
 sky130_fd_sc_hd__and2_1 _6542_ (.A(_3155_),
    .B(_3177_),
    .X(_3178_));
 sky130_fd_sc_hd__xnor2_1 _6543_ (.A(_3176_),
    .B(_3178_),
    .Y(_3179_));
 sky130_fd_sc_hd__xnor2_1 _6544_ (.A(_3175_),
    .B(_3179_),
    .Y(_3180_));
 sky130_fd_sc_hd__xor2_1 _6545_ (.A(_2380_),
    .B(_2420_),
    .X(_3181_));
 sky130_fd_sc_hd__xor2_1 _6546_ (.A(_2509_),
    .B(_2539_),
    .X(_3182_));
 sky130_fd_sc_hd__xnor2_1 _6547_ (.A(_2451_),
    .B(_2476_),
    .Y(_3183_));
 sky130_fd_sc_hd__xnor2_1 _6548_ (.A(_3182_),
    .B(_3183_),
    .Y(_3184_));
 sky130_fd_sc_hd__xnor2_1 _6549_ (.A(_3181_),
    .B(_3184_),
    .Y(_3185_));
 sky130_fd_sc_hd__xnor2_1 _6550_ (.A(_3180_),
    .B(_3185_),
    .Y(_3186_));
 sky130_fd_sc_hd__xnor2_1 _6551_ (.A(_2566_),
    .B(_2596_),
    .Y(_3187_));
 sky130_fd_sc_hd__nand2_1 _6552_ (.A(_2323_),
    .B(_2360_),
    .Y(_3188_));
 sky130_fd_sc_hd__and2_1 _6553_ (.A(_3153_),
    .B(_3188_),
    .X(_3189_));
 sky130_fd_sc_hd__xnor2_1 _6554_ (.A(_3187_),
    .B(_3189_),
    .Y(_3190_));
 sky130_fd_sc_hd__xnor2_1 _6555_ (.A(_3186_),
    .B(_3190_),
    .Y(_3191_));
 sky130_fd_sc_hd__nand2_1 _6556_ (.A(net204),
    .B(_3150_),
    .Y(_3192_));
 sky130_fd_sc_hd__o211a_1 _6557_ (.A1(_3150_),
    .A2(_3191_),
    .B1(_3192_),
    .C1(_3151_),
    .X(_3193_));
 sky130_fd_sc_hd__nor3_1 _6558_ (.A(_1122_),
    .B(_3174_),
    .C(_3193_),
    .Y(_0455_));
 sky130_fd_sc_hd__nand2_1 _6559_ (.A(_1153_),
    .B(_2332_),
    .Y(_3194_));
 sky130_fd_sc_hd__inv_2 _6560_ (.A(_3194_),
    .Y(_3195_));
 sky130_fd_sc_hd__a21o_2 _6561_ (.A1(_1071_),
    .A2(_3195_),
    .B1(_0670_),
    .X(_3196_));
 sky130_fd_sc_hd__clkbuf_4 _6562_ (.A(_3196_),
    .X(_3197_));
 sky130_fd_sc_hd__a21oi_4 _6563_ (.A1(_1071_),
    .A2(_3195_),
    .B1(_0670_),
    .Y(_3198_));
 sky130_fd_sc_hd__mux2_1 _6564_ (.A0(net211),
    .A1(\core_1.execute.mem_stage_pc[0] ),
    .S(net37),
    .X(_3199_));
 sky130_fd_sc_hd__buf_4 _6565_ (.A(_3194_),
    .X(_3200_));
 sky130_fd_sc_hd__mux2_1 _6566_ (.A0(net194),
    .A1(_3199_),
    .S(_3200_),
    .X(_3201_));
 sky130_fd_sc_hd__or2_1 _6567_ (.A(_3198_),
    .B(_3201_),
    .X(_3202_));
 sky130_fd_sc_hd__o211a_1 _6568_ (.A1(\core_1.execute.sreg_irq_pc.o_d[0] ),
    .A2(_3197_),
    .B1(_3202_),
    .C1(_2842_),
    .X(_0456_));
 sky130_fd_sc_hd__mux2_1 _6569_ (.A0(net79),
    .A1(\core_1.execute.mem_stage_pc[1] ),
    .S(net37),
    .X(_3203_));
 sky130_fd_sc_hd__mux2_1 _6570_ (.A0(net201),
    .A1(_3203_),
    .S(_3200_),
    .X(_3204_));
 sky130_fd_sc_hd__or2_1 _6571_ (.A(_3198_),
    .B(_3204_),
    .X(_3205_));
 sky130_fd_sc_hd__o211a_1 _6572_ (.A1(\core_1.execute.sreg_irq_pc.o_d[1] ),
    .A2(_3197_),
    .B1(_3205_),
    .C1(_2842_),
    .X(_0457_));
 sky130_fd_sc_hd__clkbuf_4 _6573_ (.A(_3200_),
    .X(_3206_));
 sky130_fd_sc_hd__buf_4 _6574_ (.A(net37),
    .X(_3207_));
 sky130_fd_sc_hd__mux2_1 _6575_ (.A0(net80),
    .A1(\core_1.execute.mem_stage_pc[2] ),
    .S(_3207_),
    .X(_3208_));
 sky130_fd_sc_hd__clkbuf_4 _6576_ (.A(_3200_),
    .X(_3209_));
 sky130_fd_sc_hd__nor2_1 _6577_ (.A(_0647_),
    .B(_3209_),
    .Y(_3210_));
 sky130_fd_sc_hd__clkbuf_4 _6578_ (.A(_3198_),
    .X(_3211_));
 sky130_fd_sc_hd__a211o_1 _6579_ (.A1(_3206_),
    .A2(_3208_),
    .B1(_3210_),
    .C1(_3211_),
    .X(_3212_));
 sky130_fd_sc_hd__clkbuf_4 _6580_ (.A(_0998_),
    .X(_3213_));
 sky130_fd_sc_hd__o211a_1 _6581_ (.A1(\core_1.execute.sreg_irq_pc.o_d[2] ),
    .A2(_3197_),
    .B1(_3212_),
    .C1(_3213_),
    .X(_0458_));
 sky130_fd_sc_hd__mux2_1 _6582_ (.A0(net81),
    .A1(\core_1.execute.mem_stage_pc[3] ),
    .S(net37),
    .X(_3214_));
 sky130_fd_sc_hd__mux2_1 _6583_ (.A0(net203),
    .A1(_3214_),
    .S(_3194_),
    .X(_3215_));
 sky130_fd_sc_hd__or2_1 _6584_ (.A(_3198_),
    .B(_3215_),
    .X(_3216_));
 sky130_fd_sc_hd__o211a_1 _6585_ (.A1(\core_1.execute.sreg_irq_pc.o_d[3] ),
    .A2(_3197_),
    .B1(_3216_),
    .C1(_3213_),
    .X(_0459_));
 sky130_fd_sc_hd__mux2_1 _6586_ (.A0(net82),
    .A1(\core_1.execute.mem_stage_pc[4] ),
    .S(_3207_),
    .X(_3217_));
 sky130_fd_sc_hd__nor2_1 _6587_ (.A(_0633_),
    .B(_3209_),
    .Y(_3218_));
 sky130_fd_sc_hd__a211o_1 _6588_ (.A1(_3206_),
    .A2(_3217_),
    .B1(_3218_),
    .C1(_3211_),
    .X(_3219_));
 sky130_fd_sc_hd__o211a_1 _6589_ (.A1(\core_1.execute.sreg_irq_pc.o_d[4] ),
    .A2(_3197_),
    .B1(_3219_),
    .C1(_3213_),
    .X(_0460_));
 sky130_fd_sc_hd__mux2_1 _6590_ (.A0(net83),
    .A1(\core_1.execute.mem_stage_pc[5] ),
    .S(_3207_),
    .X(_3220_));
 sky130_fd_sc_hd__nor2_1 _6591_ (.A(_0627_),
    .B(_3209_),
    .Y(_3221_));
 sky130_fd_sc_hd__a211o_1 _6592_ (.A1(_3206_),
    .A2(_3220_),
    .B1(_3221_),
    .C1(_3211_),
    .X(_3222_));
 sky130_fd_sc_hd__o211a_1 _6593_ (.A1(\core_1.execute.sreg_irq_pc.o_d[5] ),
    .A2(_3197_),
    .B1(_3222_),
    .C1(_3213_),
    .X(_0461_));
 sky130_fd_sc_hd__mux2_1 _6594_ (.A0(net84),
    .A1(\core_1.execute.mem_stage_pc[6] ),
    .S(_3207_),
    .X(_3223_));
 sky130_fd_sc_hd__nor2_1 _6595_ (.A(_0621_),
    .B(_3209_),
    .Y(_3224_));
 sky130_fd_sc_hd__a211o_1 _6596_ (.A1(_3206_),
    .A2(_3223_),
    .B1(_3224_),
    .C1(_3211_),
    .X(_3225_));
 sky130_fd_sc_hd__o211a_1 _6597_ (.A1(\core_1.execute.sreg_irq_pc.o_d[6] ),
    .A2(_3197_),
    .B1(_3225_),
    .C1(_3213_),
    .X(_0462_));
 sky130_fd_sc_hd__mux2_1 _6598_ (.A0(net85),
    .A1(\core_1.execute.mem_stage_pc[7] ),
    .S(_3207_),
    .X(_3226_));
 sky130_fd_sc_hd__nor2_1 _6599_ (.A(_0614_),
    .B(_3209_),
    .Y(_3227_));
 sky130_fd_sc_hd__a211o_1 _6600_ (.A1(_3206_),
    .A2(_3226_),
    .B1(_3227_),
    .C1(_3211_),
    .X(_3228_));
 sky130_fd_sc_hd__o211a_1 _6601_ (.A1(\core_1.execute.sreg_irq_pc.o_d[7] ),
    .A2(_3197_),
    .B1(_3228_),
    .C1(_3213_),
    .X(_0463_));
 sky130_fd_sc_hd__mux2_1 _6602_ (.A0(net86),
    .A1(\core_1.execute.mem_stage_pc[8] ),
    .S(_3207_),
    .X(_3229_));
 sky130_fd_sc_hd__nor2_1 _6603_ (.A(_0606_),
    .B(_3209_),
    .Y(_3230_));
 sky130_fd_sc_hd__a211o_1 _6604_ (.A1(_3206_),
    .A2(_3229_),
    .B1(_3230_),
    .C1(_3211_),
    .X(_3231_));
 sky130_fd_sc_hd__o211a_1 _6605_ (.A1(\core_1.execute.sreg_irq_pc.o_d[8] ),
    .A2(_3197_),
    .B1(_3231_),
    .C1(_3213_),
    .X(_0464_));
 sky130_fd_sc_hd__mux2_1 _6606_ (.A0(net87),
    .A1(\core_1.execute.mem_stage_pc[9] ),
    .S(_3207_),
    .X(_3232_));
 sky130_fd_sc_hd__nor2_1 _6607_ (.A(_0600_),
    .B(_3209_),
    .Y(_3233_));
 sky130_fd_sc_hd__a211o_1 _6608_ (.A1(_3206_),
    .A2(_3232_),
    .B1(_3233_),
    .C1(_3211_),
    .X(_3234_));
 sky130_fd_sc_hd__o211a_1 _6609_ (.A1(\core_1.execute.sreg_irq_pc.o_d[9] ),
    .A2(_3197_),
    .B1(_3234_),
    .C1(_3213_),
    .X(_0465_));
 sky130_fd_sc_hd__mux2_1 _6610_ (.A0(net73),
    .A1(\core_1.execute.mem_stage_pc[10] ),
    .S(_3207_),
    .X(_3235_));
 sky130_fd_sc_hd__nor2_1 _6611_ (.A(_0593_),
    .B(_3200_),
    .Y(_3236_));
 sky130_fd_sc_hd__a211o_1 _6612_ (.A1(_3206_),
    .A2(_3235_),
    .B1(_3236_),
    .C1(_3211_),
    .X(_3237_));
 sky130_fd_sc_hd__o211a_1 _6613_ (.A1(\core_1.execute.sreg_irq_pc.o_d[10] ),
    .A2(_3196_),
    .B1(_3237_),
    .C1(_3213_),
    .X(_0466_));
 sky130_fd_sc_hd__mux2_1 _6614_ (.A0(net74),
    .A1(\core_1.execute.mem_stage_pc[11] ),
    .S(_3207_),
    .X(_3238_));
 sky130_fd_sc_hd__nor2_1 _6615_ (.A(_0585_),
    .B(_3200_),
    .Y(_3239_));
 sky130_fd_sc_hd__a211o_1 _6616_ (.A1(_3206_),
    .A2(_3238_),
    .B1(_3239_),
    .C1(_3211_),
    .X(_3240_));
 sky130_fd_sc_hd__o211a_1 _6617_ (.A1(\core_1.execute.sreg_irq_pc.o_d[11] ),
    .A2(_3196_),
    .B1(_3240_),
    .C1(_3213_),
    .X(_0467_));
 sky130_fd_sc_hd__mux2_1 _6618_ (.A0(net75),
    .A1(\core_1.execute.mem_stage_pc[12] ),
    .S(net37),
    .X(_3241_));
 sky130_fd_sc_hd__nor2_1 _6619_ (.A(_0577_),
    .B(_3200_),
    .Y(_3242_));
 sky130_fd_sc_hd__a211o_1 _6620_ (.A1(_3206_),
    .A2(_3241_),
    .B1(_3242_),
    .C1(_3211_),
    .X(_3243_));
 sky130_fd_sc_hd__buf_6 _6621_ (.A(_0998_),
    .X(_3244_));
 sky130_fd_sc_hd__o211a_1 _6622_ (.A1(\core_1.execute.sreg_irq_pc.o_d[12] ),
    .A2(_3196_),
    .B1(_3243_),
    .C1(_3244_),
    .X(_0468_));
 sky130_fd_sc_hd__mux2_1 _6623_ (.A0(net76),
    .A1(\core_1.execute.mem_stage_pc[13] ),
    .S(net37),
    .X(_3245_));
 sky130_fd_sc_hd__nor2_1 _6624_ (.A(_0571_),
    .B(_3200_),
    .Y(_3246_));
 sky130_fd_sc_hd__a211o_1 _6625_ (.A1(_3209_),
    .A2(_3245_),
    .B1(_3246_),
    .C1(_3198_),
    .X(_3247_));
 sky130_fd_sc_hd__o211a_1 _6626_ (.A1(\core_1.execute.sreg_irq_pc.o_d[13] ),
    .A2(_3196_),
    .B1(_3247_),
    .C1(_3244_),
    .X(_0469_));
 sky130_fd_sc_hd__mux2_1 _6627_ (.A0(net77),
    .A1(\core_1.execute.mem_stage_pc[14] ),
    .S(net37),
    .X(_3248_));
 sky130_fd_sc_hd__nor2_1 _6628_ (.A(_0556_),
    .B(_3200_),
    .Y(_3249_));
 sky130_fd_sc_hd__a211o_1 _6629_ (.A1(_3209_),
    .A2(_3248_),
    .B1(_3249_),
    .C1(_3198_),
    .X(_3250_));
 sky130_fd_sc_hd__o211a_1 _6630_ (.A1(\core_1.execute.sreg_irq_pc.o_d[14] ),
    .A2(_3196_),
    .B1(_3250_),
    .C1(_3244_),
    .X(_0470_));
 sky130_fd_sc_hd__mux2_1 _6631_ (.A0(net78),
    .A1(\core_1.execute.mem_stage_pc[15] ),
    .S(net37),
    .X(_3251_));
 sky130_fd_sc_hd__nor2_1 _6632_ (.A(_0545_),
    .B(_3200_),
    .Y(_3252_));
 sky130_fd_sc_hd__a211o_1 _6633_ (.A1(_3209_),
    .A2(_3251_),
    .B1(_3252_),
    .C1(_3198_),
    .X(_3253_));
 sky130_fd_sc_hd__o211a_1 _6634_ (.A1(\core_1.execute.sreg_irq_pc.o_d[15] ),
    .A2(_3196_),
    .B1(_3253_),
    .C1(_3244_),
    .X(_0471_));
 sky130_fd_sc_hd__and4_2 _6635_ (.A(\core_1.execute.sreg_priv_control.o_d[0] ),
    .B(_1153_),
    .C(_0737_),
    .D(_2127_),
    .X(_3254_));
 sky130_fd_sc_hd__nor2_1 _6636_ (.A(_0670_),
    .B(_3254_),
    .Y(_3255_));
 sky130_fd_sc_hd__a22o_1 _6637_ (.A1(net194),
    .A2(_3254_),
    .B1(_3255_),
    .B2(\core_1.execute.sreg_jtr_buff.o_d[0] ),
    .X(_3256_));
 sky130_fd_sc_hd__and2_1 _6638_ (.A(_1307_),
    .B(_3256_),
    .X(_3257_));
 sky130_fd_sc_hd__clkbuf_1 _6639_ (.A(_3257_),
    .X(_0472_));
 sky130_fd_sc_hd__a22o_1 _6640_ (.A1(net201),
    .A2(_3254_),
    .B1(_3255_),
    .B2(\core_1.execute.sreg_jtr_buff.o_d[1] ),
    .X(_3258_));
 sky130_fd_sc_hd__and2_1 _6641_ (.A(_1307_),
    .B(_3258_),
    .X(_3259_));
 sky130_fd_sc_hd__clkbuf_1 _6642_ (.A(_3259_),
    .X(_0473_));
 sky130_fd_sc_hd__a22o_1 _6643_ (.A1(net202),
    .A2(_3254_),
    .B1(_3255_),
    .B2(\core_1.execute.sreg_jtr_buff.o_d[2] ),
    .X(_3260_));
 sky130_fd_sc_hd__and2_1 _6644_ (.A(_1307_),
    .B(_3260_),
    .X(_3261_));
 sky130_fd_sc_hd__clkbuf_1 _6645_ (.A(_3261_),
    .X(_0474_));
 sky130_fd_sc_hd__nor2_1 _6646_ (.A(_0670_),
    .B(_1059_),
    .Y(_3262_));
 sky130_fd_sc_hd__nand2_1 _6647_ (.A(net106),
    .B(_3262_),
    .Y(_3263_));
 sky130_fd_sc_hd__a21oi_1 _6648_ (.A1(_1064_),
    .A2(_3263_),
    .B1(_1122_),
    .Y(_0475_));
 sky130_fd_sc_hd__a22o_1 _6649_ (.A1(\core_1.execute.sreg_jtr_buff.o_d[1] ),
    .A2(_1059_),
    .B1(_3262_),
    .B2(\core_1.execute.trap_flag ),
    .X(_3264_));
 sky130_fd_sc_hd__and2_1 _6650_ (.A(_1307_),
    .B(_3264_),
    .X(_3265_));
 sky130_fd_sc_hd__clkbuf_1 _6651_ (.A(_3265_),
    .X(_0476_));
 sky130_fd_sc_hd__a22o_1 _6652_ (.A1(\core_1.execute.sreg_jtr_buff.o_d[2] ),
    .A2(_1059_),
    .B1(_3262_),
    .B2(_0671_),
    .X(_3266_));
 sky130_fd_sc_hd__and2_1 _6653_ (.A(_1307_),
    .B(_3266_),
    .X(_3267_));
 sky130_fd_sc_hd__clkbuf_1 _6654_ (.A(_3267_),
    .X(_0477_));
 sky130_fd_sc_hd__and3_4 _6655_ (.A(_1153_),
    .B(_1071_),
    .C(_2331_),
    .X(_3268_));
 sky130_fd_sc_hd__clkinv_2 _6656_ (.A(_3268_),
    .Y(_3269_));
 sky130_fd_sc_hd__buf_4 _6657_ (.A(_3269_),
    .X(_3270_));
 sky130_fd_sc_hd__clkbuf_4 _6658_ (.A(_3268_),
    .X(_3271_));
 sky130_fd_sc_hd__or2_1 _6659_ (.A(\core_1.execute.sreg_scratch.o_d[0] ),
    .B(_3271_),
    .X(_3272_));
 sky130_fd_sc_hd__o211a_1 _6660_ (.A1(net194),
    .A2(_3270_),
    .B1(_3272_),
    .C1(_3244_),
    .X(_0478_));
 sky130_fd_sc_hd__or2_1 _6661_ (.A(\core_1.execute.sreg_scratch.o_d[1] ),
    .B(_3271_),
    .X(_3273_));
 sky130_fd_sc_hd__o211a_1 _6662_ (.A1(net201),
    .A2(_3270_),
    .B1(_3273_),
    .C1(_3244_),
    .X(_0479_));
 sky130_fd_sc_hd__or2_1 _6663_ (.A(\core_1.execute.sreg_scratch.o_d[2] ),
    .B(_3271_),
    .X(_3274_));
 sky130_fd_sc_hd__o211a_1 _6664_ (.A1(net202),
    .A2(_3270_),
    .B1(_3274_),
    .C1(_3244_),
    .X(_0480_));
 sky130_fd_sc_hd__or2_1 _6665_ (.A(\core_1.execute.sreg_scratch.o_d[3] ),
    .B(_3271_),
    .X(_3275_));
 sky130_fd_sc_hd__o211a_1 _6666_ (.A1(net203),
    .A2(_3270_),
    .B1(_3275_),
    .C1(_3244_),
    .X(_0481_));
 sky130_fd_sc_hd__or2_1 _6667_ (.A(\core_1.execute.sreg_scratch.o_d[4] ),
    .B(_3271_),
    .X(_3276_));
 sky130_fd_sc_hd__o211a_1 _6668_ (.A1(net204),
    .A2(_3270_),
    .B1(_3276_),
    .C1(_3244_),
    .X(_0482_));
 sky130_fd_sc_hd__or2_1 _6669_ (.A(\core_1.execute.sreg_scratch.o_d[5] ),
    .B(_3271_),
    .X(_3277_));
 sky130_fd_sc_hd__o211a_1 _6670_ (.A1(net205),
    .A2(_3270_),
    .B1(_3277_),
    .C1(_3244_),
    .X(_0483_));
 sky130_fd_sc_hd__or2_1 _6671_ (.A(\core_1.execute.sreg_scratch.o_d[6] ),
    .B(_3271_),
    .X(_3278_));
 sky130_fd_sc_hd__buf_4 _6672_ (.A(_0998_),
    .X(_3279_));
 sky130_fd_sc_hd__o211a_1 _6673_ (.A1(net206),
    .A2(_3270_),
    .B1(_3278_),
    .C1(_3279_),
    .X(_0484_));
 sky130_fd_sc_hd__or2_1 _6674_ (.A(\core_1.execute.sreg_scratch.o_d[7] ),
    .B(_3271_),
    .X(_3280_));
 sky130_fd_sc_hd__o211a_1 _6675_ (.A1(net207),
    .A2(_3270_),
    .B1(_3280_),
    .C1(_3279_),
    .X(_0485_));
 sky130_fd_sc_hd__or2_1 _6676_ (.A(\core_1.execute.sreg_scratch.o_d[8] ),
    .B(_3271_),
    .X(_3281_));
 sky130_fd_sc_hd__o211a_1 _6677_ (.A1(net208),
    .A2(_3270_),
    .B1(_3281_),
    .C1(_3279_),
    .X(_0486_));
 sky130_fd_sc_hd__or2_1 _6678_ (.A(\core_1.execute.sreg_scratch.o_d[9] ),
    .B(_3271_),
    .X(_3282_));
 sky130_fd_sc_hd__o211a_1 _6679_ (.A1(net209),
    .A2(_3270_),
    .B1(_3282_),
    .C1(_3279_),
    .X(_0487_));
 sky130_fd_sc_hd__or2_1 _6680_ (.A(\core_1.execute.sreg_scratch.o_d[10] ),
    .B(_3268_),
    .X(_3283_));
 sky130_fd_sc_hd__o211a_1 _6681_ (.A1(net195),
    .A2(_3269_),
    .B1(_3283_),
    .C1(_3279_),
    .X(_0488_));
 sky130_fd_sc_hd__or2_1 _6682_ (.A(\core_1.execute.sreg_scratch.o_d[11] ),
    .B(_3268_),
    .X(_3284_));
 sky130_fd_sc_hd__o211a_1 _6683_ (.A1(net196),
    .A2(_3269_),
    .B1(_3284_),
    .C1(_3279_),
    .X(_0489_));
 sky130_fd_sc_hd__or2_1 _6684_ (.A(\core_1.execute.sreg_scratch.o_d[12] ),
    .B(_3268_),
    .X(_3285_));
 sky130_fd_sc_hd__o211a_1 _6685_ (.A1(net197),
    .A2(_3269_),
    .B1(_3285_),
    .C1(_3279_),
    .X(_0490_));
 sky130_fd_sc_hd__or2_1 _6686_ (.A(\core_1.execute.sreg_scratch.o_d[13] ),
    .B(_3268_),
    .X(_3286_));
 sky130_fd_sc_hd__o211a_1 _6687_ (.A1(net198),
    .A2(_3269_),
    .B1(_3286_),
    .C1(_3279_),
    .X(_0491_));
 sky130_fd_sc_hd__or2_1 _6688_ (.A(\core_1.execute.sreg_scratch.o_d[14] ),
    .B(_3268_),
    .X(_3287_));
 sky130_fd_sc_hd__o211a_1 _6689_ (.A1(net199),
    .A2(_3269_),
    .B1(_3287_),
    .C1(_3279_),
    .X(_0492_));
 sky130_fd_sc_hd__or2_1 _6690_ (.A(\core_1.execute.sreg_scratch.o_d[15] ),
    .B(_3268_),
    .X(_3288_));
 sky130_fd_sc_hd__o211a_1 _6691_ (.A1(net200),
    .A2(_3269_),
    .B1(_3288_),
    .C1(_3279_),
    .X(_0493_));
 sky130_fd_sc_hd__a32o_1 _6692_ (.A1(\core_1.execute.irq_en ),
    .A2(net18),
    .A3(_1075_),
    .B1(_3070_),
    .B2(\core_1.execute.sreg_irq_flags.o_d[0] ),
    .X(_0494_));
 sky130_fd_sc_hd__inv_2 _6693_ (.A(\core_1.execute.sreg_irq_flags.o_d[1] ),
    .Y(_3289_));
 sky130_fd_sc_hd__nor2_1 _6694_ (.A(_3289_),
    .B(_0668_),
    .Y(_3290_));
 sky130_fd_sc_hd__o21a_1 _6695_ (.A1(\core_1.execute.prev_sys ),
    .A2(_3290_),
    .B1(_0999_),
    .X(_0495_));
 sky130_fd_sc_hd__a22o_1 _6696_ (.A1(\core_1.execute.sreg_irq_flags.i_d[2] ),
    .A2(_1075_),
    .B1(_3071_),
    .B2(\core_1.execute.sreg_irq_flags.o_d[2] ),
    .X(_0496_));
 sky130_fd_sc_hd__a22o_1 _6697_ (.A1(_3207_),
    .A2(_1075_),
    .B1(_3071_),
    .B2(\core_1.execute.sreg_irq_flags.o_d[3] ),
    .X(_0497_));
 sky130_fd_sc_hd__a32o_1 _6698_ (.A1(\core_1.execute.irq_en ),
    .A2(net19),
    .A3(_1068_),
    .B1(_3070_),
    .B2(\core_1.execute.sreg_irq_flags.o_d[4] ),
    .X(_0498_));
 sky130_fd_sc_hd__and2_1 _6699_ (.A(_0671_),
    .B(_1059_),
    .X(_3291_));
 sky130_fd_sc_hd__and3_2 _6700_ (.A(\core_1.dec_sreg_store ),
    .B(_1056_),
    .C(_2064_),
    .X(_3292_));
 sky130_fd_sc_hd__a311o_1 _6701_ (.A1(_0671_),
    .A2(net77),
    .A3(_1681_),
    .B1(_3291_),
    .C1(_3292_),
    .X(_3293_));
 sky130_fd_sc_hd__and2_1 _6702_ (.A(_1029_),
    .B(_3293_),
    .X(_3294_));
 sky130_fd_sc_hd__buf_2 _6703_ (.A(_3294_),
    .X(_3295_));
 sky130_fd_sc_hd__nand2_2 _6704_ (.A(_0671_),
    .B(_1059_),
    .Y(_3296_));
 sky130_fd_sc_hd__buf_2 _6705_ (.A(_3296_),
    .X(_3297_));
 sky130_fd_sc_hd__nand2_1 _6706_ (.A(\core_1.execute.pc_high_out[0] ),
    .B(_3297_),
    .Y(_3298_));
 sky130_fd_sc_hd__nand2_4 _6707_ (.A(_1153_),
    .B(_2129_),
    .Y(_3299_));
 sky130_fd_sc_hd__o211a_1 _6708_ (.A1(\core_1.execute.pc_high_buff_out[0] ),
    .A2(_3297_),
    .B1(_3298_),
    .C1(_3299_),
    .X(_3300_));
 sky130_fd_sc_hd__nand2_4 _6709_ (.A(_1029_),
    .B(_3293_),
    .Y(_3301_));
 sky130_fd_sc_hd__a211o_1 _6710_ (.A1(net194),
    .A2(_3292_),
    .B1(_3300_),
    .C1(_3301_),
    .X(_3302_));
 sky130_fd_sc_hd__clkbuf_4 _6711_ (.A(_0998_),
    .X(_3303_));
 sky130_fd_sc_hd__o211a_1 _6712_ (.A1(\core_1.execute.pc_high_out[0] ),
    .A2(_3295_),
    .B1(_3302_),
    .C1(_3303_),
    .X(_0499_));
 sky130_fd_sc_hd__nand2_1 _6713_ (.A(\core_1.execute.pc_high_out[1] ),
    .B(\core_1.execute.pc_high_out[0] ),
    .Y(_3304_));
 sky130_fd_sc_hd__o21a_1 _6714_ (.A1(\core_1.execute.pc_high_out[1] ),
    .A2(\core_1.execute.pc_high_out[0] ),
    .B1(_3296_),
    .X(_3305_));
 sky130_fd_sc_hd__a22o_1 _6715_ (.A1(\core_1.execute.pc_high_buff_out[1] ),
    .A2(_3291_),
    .B1(_3304_),
    .B2(_3305_),
    .X(_3306_));
 sky130_fd_sc_hd__mux2_1 _6716_ (.A0(net201),
    .A1(_3306_),
    .S(_3299_),
    .X(_3307_));
 sky130_fd_sc_hd__or2_1 _6717_ (.A(\core_1.execute.pc_high_out[1] ),
    .B(_3295_),
    .X(_3308_));
 sky130_fd_sc_hd__o211a_1 _6718_ (.A1(_3301_),
    .A2(_3307_),
    .B1(_3308_),
    .C1(_3303_),
    .X(_0500_));
 sky130_fd_sc_hd__xor2_1 _6719_ (.A(\core_1.execute.pc_high_out[2] ),
    .B(_3304_),
    .X(_3309_));
 sky130_fd_sc_hd__a21oi_1 _6720_ (.A1(_3297_),
    .A2(_3309_),
    .B1(_3292_),
    .Y(_3310_));
 sky130_fd_sc_hd__or2_1 _6721_ (.A(\core_1.execute.pc_high_buff_out[2] ),
    .B(_3297_),
    .X(_3311_));
 sky130_fd_sc_hd__a221o_1 _6722_ (.A1(net202),
    .A2(_3292_),
    .B1(_3310_),
    .B2(_3311_),
    .C1(_3301_),
    .X(_3312_));
 sky130_fd_sc_hd__o211a_1 _6723_ (.A1(\core_1.execute.pc_high_out[2] ),
    .A2(_3295_),
    .B1(_3312_),
    .C1(_3303_),
    .X(_0501_));
 sky130_fd_sc_hd__and4_1 _6724_ (.A(\core_1.execute.pc_high_out[3] ),
    .B(\core_1.execute.pc_high_out[2] ),
    .C(\core_1.execute.pc_high_out[1] ),
    .D(\core_1.execute.pc_high_out[0] ),
    .X(_3313_));
 sky130_fd_sc_hd__a31oi_1 _6725_ (.A1(\core_1.execute.pc_high_out[2] ),
    .A2(\core_1.execute.pc_high_out[1] ),
    .A3(\core_1.execute.pc_high_out[0] ),
    .B1(\core_1.execute.pc_high_out[3] ),
    .Y(_3314_));
 sky130_fd_sc_hd__o21ai_1 _6726_ (.A1(_3313_),
    .A2(_3314_),
    .B1(_3297_),
    .Y(_3315_));
 sky130_fd_sc_hd__o211a_1 _6727_ (.A1(\core_1.execute.pc_high_buff_out[3] ),
    .A2(_3297_),
    .B1(_3299_),
    .C1(_3315_),
    .X(_3316_));
 sky130_fd_sc_hd__a211o_1 _6728_ (.A1(net203),
    .A2(_3292_),
    .B1(_3301_),
    .C1(_3316_),
    .X(_3317_));
 sky130_fd_sc_hd__o211a_1 _6729_ (.A1(\core_1.execute.pc_high_out[3] ),
    .A2(_3295_),
    .B1(_3317_),
    .C1(_3303_),
    .X(_0502_));
 sky130_fd_sc_hd__nand2_1 _6730_ (.A(\core_1.execute.pc_high_out[4] ),
    .B(_3313_),
    .Y(_3318_));
 sky130_fd_sc_hd__o21a_1 _6731_ (.A1(\core_1.execute.pc_high_out[4] ),
    .A2(_3313_),
    .B1(_3296_),
    .X(_3319_));
 sky130_fd_sc_hd__a22o_1 _6732_ (.A1(\core_1.execute.pc_high_buff_out[4] ),
    .A2(_3291_),
    .B1(_3318_),
    .B2(_3319_),
    .X(_3320_));
 sky130_fd_sc_hd__nor2_1 _6733_ (.A(_0633_),
    .B(_3299_),
    .Y(_3321_));
 sky130_fd_sc_hd__a211o_1 _6734_ (.A1(_3299_),
    .A2(_3320_),
    .B1(_3321_),
    .C1(_3301_),
    .X(_3322_));
 sky130_fd_sc_hd__o211a_1 _6735_ (.A1(\core_1.execute.pc_high_out[4] ),
    .A2(_3295_),
    .B1(_3322_),
    .C1(_3303_),
    .X(_0503_));
 sky130_fd_sc_hd__and3_1 _6736_ (.A(\core_1.execute.pc_high_out[5] ),
    .B(\core_1.execute.pc_high_out[4] ),
    .C(_3313_),
    .X(_3323_));
 sky130_fd_sc_hd__a21oi_1 _6737_ (.A1(\core_1.execute.pc_high_out[4] ),
    .A2(_3313_),
    .B1(\core_1.execute.pc_high_out[5] ),
    .Y(_3324_));
 sky130_fd_sc_hd__o21ai_1 _6738_ (.A1(_3323_),
    .A2(_3324_),
    .B1(_3297_),
    .Y(_3325_));
 sky130_fd_sc_hd__o211a_1 _6739_ (.A1(\core_1.execute.pc_high_buff_out[5] ),
    .A2(_3297_),
    .B1(_3299_),
    .C1(_3325_),
    .X(_3326_));
 sky130_fd_sc_hd__a211o_1 _6740_ (.A1(net205),
    .A2(_3292_),
    .B1(_3301_),
    .C1(_3326_),
    .X(_3327_));
 sky130_fd_sc_hd__o211a_1 _6741_ (.A1(\core_1.execute.pc_high_out[5] ),
    .A2(_3295_),
    .B1(_3327_),
    .C1(_3303_),
    .X(_0504_));
 sky130_fd_sc_hd__and2_1 _6742_ (.A(\core_1.execute.pc_high_out[6] ),
    .B(_3323_),
    .X(_3328_));
 sky130_fd_sc_hd__nor2_1 _6743_ (.A(\core_1.execute.pc_high_out[6] ),
    .B(_3323_),
    .Y(_3329_));
 sky130_fd_sc_hd__o21ai_1 _6744_ (.A1(_3328_),
    .A2(_3329_),
    .B1(_3297_),
    .Y(_3330_));
 sky130_fd_sc_hd__o211a_1 _6745_ (.A1(\core_1.execute.pc_high_buff_out[6] ),
    .A2(_3297_),
    .B1(_3299_),
    .C1(_3330_),
    .X(_3331_));
 sky130_fd_sc_hd__a211o_1 _6746_ (.A1(net206),
    .A2(_3292_),
    .B1(_3301_),
    .C1(_3331_),
    .X(_3332_));
 sky130_fd_sc_hd__o211a_1 _6747_ (.A1(\core_1.execute.pc_high_out[6] ),
    .A2(_3295_),
    .B1(_3332_),
    .C1(_3303_),
    .X(_0505_));
 sky130_fd_sc_hd__inv_2 _6748_ (.A(\core_1.execute.pc_high_buff_out[7] ),
    .Y(_3333_));
 sky130_fd_sc_hd__xnor2_1 _6749_ (.A(\core_1.execute.pc_high_out[7] ),
    .B(_3328_),
    .Y(_3334_));
 sky130_fd_sc_hd__mux2_1 _6750_ (.A0(_3333_),
    .A1(_3334_),
    .S(_3296_),
    .X(_3335_));
 sky130_fd_sc_hd__nand2_1 _6751_ (.A(_3299_),
    .B(_3335_),
    .Y(_3336_));
 sky130_fd_sc_hd__o211a_1 _6752_ (.A1(net207),
    .A2(_3299_),
    .B1(_3295_),
    .C1(_3336_),
    .X(_3337_));
 sky130_fd_sc_hd__a211o_1 _6753_ (.A1(\core_1.execute.pc_high_out[7] ),
    .A2(_3301_),
    .B1(_3337_),
    .C1(_1122_),
    .X(_0506_));
 sky130_fd_sc_hd__and3_1 _6754_ (.A(_1153_),
    .B(_1160_),
    .C(_2064_),
    .X(_3338_));
 sky130_fd_sc_hd__a21o_1 _6755_ (.A1(_0671_),
    .A2(\core_1.dec_sreg_jal_over ),
    .B1(_3338_),
    .X(_3339_));
 sky130_fd_sc_hd__and2_1 _6756_ (.A(_0737_),
    .B(_3339_),
    .X(_3340_));
 sky130_fd_sc_hd__buf_2 _6757_ (.A(_3340_),
    .X(_3341_));
 sky130_fd_sc_hd__clkbuf_4 _6758_ (.A(_3341_),
    .X(_3342_));
 sky130_fd_sc_hd__buf_4 _6759_ (.A(_3338_),
    .X(_3343_));
 sky130_fd_sc_hd__mux2_1 _6760_ (.A0(_0685_),
    .A1(_0661_),
    .S(_3343_),
    .X(_3344_));
 sky130_fd_sc_hd__nand2_1 _6761_ (.A(_3342_),
    .B(_3344_),
    .Y(_3345_));
 sky130_fd_sc_hd__o211a_1 _6762_ (.A1(\core_1.execute.pc_high_buff_out[0] ),
    .A2(_3342_),
    .B1(_3345_),
    .C1(_3303_),
    .X(_0507_));
 sky130_fd_sc_hd__nand2_1 _6763_ (.A(net201),
    .B(_3343_),
    .Y(_3346_));
 sky130_fd_sc_hd__o211ai_1 _6764_ (.A1(_0683_),
    .A2(_3343_),
    .B1(_3341_),
    .C1(_3346_),
    .Y(_3347_));
 sky130_fd_sc_hd__o211a_1 _6765_ (.A1(\core_1.execute.pc_high_buff_out[1] ),
    .A2(_3342_),
    .B1(_3347_),
    .C1(_3303_),
    .X(_0508_));
 sky130_fd_sc_hd__mux2_1 _6766_ (.A0(_0672_),
    .A1(_0647_),
    .S(_3343_),
    .X(_3348_));
 sky130_fd_sc_hd__nand2_1 _6767_ (.A(_3342_),
    .B(_3348_),
    .Y(_3349_));
 sky130_fd_sc_hd__o211a_1 _6768_ (.A1(\core_1.execute.pc_high_buff_out[2] ),
    .A2(_3342_),
    .B1(_3349_),
    .C1(_3303_),
    .X(_0509_));
 sky130_fd_sc_hd__nand2_1 _6769_ (.A(net203),
    .B(_3343_),
    .Y(_3350_));
 sky130_fd_sc_hd__o211ai_1 _6770_ (.A1(_0674_),
    .A2(_3343_),
    .B1(_3341_),
    .C1(_3350_),
    .Y(_3351_));
 sky130_fd_sc_hd__o211a_1 _6771_ (.A1(\core_1.execute.pc_high_buff_out[3] ),
    .A2(_3342_),
    .B1(_3351_),
    .C1(_1075_),
    .X(_0510_));
 sky130_fd_sc_hd__mux2_1 _6772_ (.A0(_0678_),
    .A1(_0633_),
    .S(_3343_),
    .X(_3352_));
 sky130_fd_sc_hd__nand2_1 _6773_ (.A(_3342_),
    .B(_3352_),
    .Y(_3353_));
 sky130_fd_sc_hd__o211a_1 _6774_ (.A1(\core_1.execute.pc_high_buff_out[4] ),
    .A2(_3342_),
    .B1(_3353_),
    .C1(_1075_),
    .X(_0511_));
 sky130_fd_sc_hd__mux2_1 _6775_ (.A0(_0681_),
    .A1(_0627_),
    .S(_3343_),
    .X(_3354_));
 sky130_fd_sc_hd__nand2_1 _6776_ (.A(_3341_),
    .B(_3354_),
    .Y(_3355_));
 sky130_fd_sc_hd__o211a_1 _6777_ (.A1(\core_1.execute.pc_high_buff_out[5] ),
    .A2(_3342_),
    .B1(_3355_),
    .C1(_1075_),
    .X(_0512_));
 sky130_fd_sc_hd__mux2_1 _6778_ (.A0(_0677_),
    .A1(_0621_),
    .S(_3343_),
    .X(_3356_));
 sky130_fd_sc_hd__nand2_1 _6779_ (.A(_3341_),
    .B(_3356_),
    .Y(_3357_));
 sky130_fd_sc_hd__o211a_1 _6780_ (.A1(\core_1.execute.pc_high_buff_out[6] ),
    .A2(_3342_),
    .B1(_3357_),
    .C1(_1075_),
    .X(_0513_));
 sky130_fd_sc_hd__mux2_1 _6781_ (.A0(_0673_),
    .A1(_0614_),
    .S(_3343_),
    .X(_3358_));
 sky130_fd_sc_hd__mux2_1 _6782_ (.A0(_3333_),
    .A1(_3358_),
    .S(_3341_),
    .X(_3359_));
 sky130_fd_sc_hd__nand2_1 _6783_ (.A(_0999_),
    .B(_3359_),
    .Y(_0514_));
 sky130_fd_sc_hd__dfxtp_4 _6784_ (.CLK(clknet_leaf_45_i_clk),
    .D(_0015_),
    .Q(\core_1.decode.o_submit ));
 sky130_fd_sc_hd__dfxtp_1 _6785_ (.CLK(clknet_leaf_45_i_clk),
    .D(_0016_),
    .Q(\core_1.dec_pc_inc ));
 sky130_fd_sc_hd__dfxtp_4 _6786_ (.CLK(clknet_leaf_45_i_clk),
    .D(_0017_),
    .Q(\core_1.dec_r_bus_imm ));
 sky130_fd_sc_hd__dfxtp_1 _6787_ (.CLK(clknet_leaf_45_i_clk),
    .D(_0018_),
    .Q(\core_1.dec_alu_flags_ie ));
 sky130_fd_sc_hd__dfxtp_1 _6788_ (.CLK(clknet_leaf_45_i_clk),
    .D(_0019_),
    .Q(\core_1.dec_alu_carry_en ));
 sky130_fd_sc_hd__dfxtp_4 _6789_ (.CLK(clknet_leaf_4_i_clk),
    .D(_0020_),
    .Q(\core_1.dec_l_reg_sel[0] ));
 sky130_fd_sc_hd__dfxtp_1 _6790_ (.CLK(clknet_leaf_4_i_clk),
    .D(_0021_),
    .Q(\core_1.dec_l_reg_sel[1] ));
 sky130_fd_sc_hd__dfxtp_1 _6791_ (.CLK(clknet_leaf_31_i_clk),
    .D(_0022_),
    .Q(\core_1.dec_l_reg_sel[2] ));
 sky130_fd_sc_hd__dfxtp_1 _6792_ (.CLK(clknet_leaf_16_i_clk),
    .D(_0023_),
    .Q(\core_1.dec_r_reg_sel[0] ));
 sky130_fd_sc_hd__dfxtp_1 _6793_ (.CLK(clknet_leaf_16_i_clk),
    .D(_0024_),
    .Q(\core_1.dec_r_reg_sel[1] ));
 sky130_fd_sc_hd__dfxtp_1 _6794_ (.CLK(clknet_leaf_16_i_clk),
    .D(_0025_),
    .Q(\core_1.dec_r_reg_sel[2] ));
 sky130_fd_sc_hd__dfxtp_1 _6795_ (.CLK(clknet_leaf_47_i_clk),
    .D(_0026_),
    .Q(\core_1.dec_rf_ie[0] ));
 sky130_fd_sc_hd__dfxtp_1 _6796_ (.CLK(clknet_leaf_31_i_clk),
    .D(_0027_),
    .Q(\core_1.dec_rf_ie[1] ));
 sky130_fd_sc_hd__dfxtp_1 _6797_ (.CLK(clknet_leaf_47_i_clk),
    .D(_0028_),
    .Q(\core_1.dec_rf_ie[2] ));
 sky130_fd_sc_hd__dfxtp_1 _6798_ (.CLK(clknet_leaf_47_i_clk),
    .D(_0029_),
    .Q(\core_1.dec_rf_ie[3] ));
 sky130_fd_sc_hd__dfxtp_1 _6799_ (.CLK(clknet_leaf_47_i_clk),
    .D(_0030_),
    .Q(\core_1.dec_rf_ie[4] ));
 sky130_fd_sc_hd__dfxtp_1 _6800_ (.CLK(clknet_leaf_31_i_clk),
    .D(_0031_),
    .Q(\core_1.dec_rf_ie[5] ));
 sky130_fd_sc_hd__dfxtp_1 _6801_ (.CLK(clknet_leaf_47_i_clk),
    .D(_0032_),
    .Q(\core_1.dec_rf_ie[6] ));
 sky130_fd_sc_hd__dfxtp_1 _6802_ (.CLK(clknet_leaf_46_i_clk),
    .D(_0033_),
    .Q(\core_1.dec_rf_ie[7] ));
 sky130_fd_sc_hd__dfxtp_1 _6803_ (.CLK(clknet_leaf_45_i_clk),
    .D(_0034_),
    .Q(\core_1.dec_jump_cond_code[0] ));
 sky130_fd_sc_hd__dfxtp_2 _6804_ (.CLK(clknet_leaf_46_i_clk),
    .D(_0035_),
    .Q(\core_1.dec_jump_cond_code[1] ));
 sky130_fd_sc_hd__dfxtp_1 _6805_ (.CLK(clknet_leaf_46_i_clk),
    .D(_0036_),
    .Q(\core_1.dec_jump_cond_code[2] ));
 sky130_fd_sc_hd__dfxtp_1 _6806_ (.CLK(clknet_leaf_46_i_clk),
    .D(_0037_),
    .Q(\core_1.dec_jump_cond_code[3] ));
 sky130_fd_sc_hd__dfxtp_1 _6807_ (.CLK(clknet_leaf_45_i_clk),
    .D(_0038_),
    .Q(\core_1.dec_jump_cond_code[4] ));
 sky130_fd_sc_hd__dfxtp_4 _6808_ (.CLK(clknet_leaf_46_i_clk),
    .D(_0039_),
    .Q(net178));
 sky130_fd_sc_hd__dfxtp_2 _6809_ (.CLK(clknet_leaf_46_i_clk),
    .D(_0040_),
    .Q(net185));
 sky130_fd_sc_hd__dfxtp_2 _6810_ (.CLK(clknet_leaf_46_i_clk),
    .D(_0041_),
    .Q(net186));
 sky130_fd_sc_hd__dfxtp_2 _6811_ (.CLK(clknet_leaf_46_i_clk),
    .D(_0042_),
    .Q(net187));
 sky130_fd_sc_hd__dfxtp_4 _6812_ (.CLK(clknet_leaf_19_i_clk),
    .D(_0043_),
    .Q(net188));
 sky130_fd_sc_hd__dfxtp_4 _6813_ (.CLK(clknet_leaf_20_i_clk),
    .D(_0044_),
    .Q(net189));
 sky130_fd_sc_hd__dfxtp_4 _6814_ (.CLK(clknet_leaf_20_i_clk),
    .D(_0045_),
    .Q(net190));
 sky130_fd_sc_hd__dfxtp_4 _6815_ (.CLK(clknet_leaf_19_i_clk),
    .D(_0046_),
    .Q(net191));
 sky130_fd_sc_hd__dfxtp_4 _6816_ (.CLK(clknet_leaf_20_i_clk),
    .D(_0047_),
    .Q(net192));
 sky130_fd_sc_hd__dfxtp_4 _6817_ (.CLK(clknet_leaf_20_i_clk),
    .D(_0048_),
    .Q(net193));
 sky130_fd_sc_hd__dfxtp_4 _6818_ (.CLK(clknet_leaf_19_i_clk),
    .D(_0049_),
    .Q(net179));
 sky130_fd_sc_hd__dfxtp_4 _6819_ (.CLK(clknet_leaf_22_i_clk),
    .D(_0050_),
    .Q(net180));
 sky130_fd_sc_hd__dfxtp_4 _6820_ (.CLK(clknet_leaf_20_i_clk),
    .D(_0051_),
    .Q(net181));
 sky130_fd_sc_hd__dfxtp_4 _6821_ (.CLK(clknet_leaf_23_i_clk),
    .D(_0052_),
    .Q(net182));
 sky130_fd_sc_hd__dfxtp_4 _6822_ (.CLK(clknet_leaf_19_i_clk),
    .D(_0053_),
    .Q(net183));
 sky130_fd_sc_hd__dfxtp_4 _6823_ (.CLK(clknet_leaf_19_i_clk),
    .D(_0054_),
    .Q(net184));
 sky130_fd_sc_hd__dfxtp_1 _6824_ (.CLK(clknet_leaf_46_i_clk),
    .D(_0055_),
    .Q(\core_1.dec_mem_access ));
 sky130_fd_sc_hd__dfxtp_1 _6825_ (.CLK(clknet_leaf_42_i_clk),
    .D(_0056_),
    .Q(\core_1.dec_mem_we ));
 sky130_fd_sc_hd__dfxtp_2 _6826_ (.CLK(clknet_leaf_45_i_clk),
    .D(_0057_),
    .Q(\core_1.dec_used_operands[0] ));
 sky130_fd_sc_hd__dfxtp_2 _6827_ (.CLK(clknet_leaf_45_i_clk),
    .D(_0058_),
    .Q(\core_1.dec_used_operands[1] ));
 sky130_fd_sc_hd__dfxtp_1 _6828_ (.CLK(clknet_leaf_42_i_clk),
    .D(_0059_),
    .Q(\core_1.dec_sreg_load ));
 sky130_fd_sc_hd__dfxtp_2 _6829_ (.CLK(clknet_leaf_42_i_clk),
    .D(_0060_),
    .Q(\core_1.dec_sreg_store ));
 sky130_fd_sc_hd__dfxtp_4 _6830_ (.CLK(clknet_leaf_45_i_clk),
    .D(_0061_),
    .Q(\core_1.dec_sreg_jal_over ));
 sky130_fd_sc_hd__dfxtp_4 _6831_ (.CLK(clknet_leaf_42_i_clk),
    .D(_0062_),
    .Q(\core_1.dec_sreg_irt ));
 sky130_fd_sc_hd__dfxtp_1 _6832_ (.CLK(clknet_leaf_43_i_clk),
    .D(_0063_),
    .Q(\core_1.dec_sys ));
 sky130_fd_sc_hd__dfxtp_1 _6833_ (.CLK(clknet_leaf_45_i_clk),
    .D(_0064_),
    .Q(\core_1.dec_mem_width ));
 sky130_fd_sc_hd__dfxtp_2 _6834_ (.CLK(clknet_leaf_43_i_clk),
    .D(_0065_),
    .Q(\core_1.dec_mem_long ));
 sky130_fd_sc_hd__dfxtp_1 _6835_ (.CLK(clknet_leaf_32_i_clk),
    .D(_0066_),
    .Q(\core_1.decode.input_valid ));
 sky130_fd_sc_hd__dfxtp_1 _6836_ (.CLK(clknet_leaf_42_i_clk),
    .D(_0067_),
    .Q(\core_1.execute.sreg_priv_control.o_d[0] ));
 sky130_fd_sc_hd__dfxtp_1 _6837_ (.CLK(clknet_leaf_39_i_clk),
    .D(_0068_),
    .Q(\core_1.execute.sreg_data_page ));
 sky130_fd_sc_hd__dfxtp_2 _6838_ (.CLK(clknet_leaf_39_i_clk),
    .D(_0069_),
    .Q(\core_1.execute.sreg_long_ptr_en ));
 sky130_fd_sc_hd__dfxtp_1 _6839_ (.CLK(clknet_leaf_37_i_clk),
    .D(_0070_),
    .Q(\core_1.execute.sreg_priv_control.o_d[4] ));
 sky130_fd_sc_hd__dfxtp_1 _6840_ (.CLK(clknet_leaf_39_i_clk),
    .D(_0071_),
    .Q(\core_1.execute.sreg_priv_control.o_d[5] ));
 sky130_fd_sc_hd__dfxtp_1 _6841_ (.CLK(clknet_leaf_37_i_clk),
    .D(_0072_),
    .Q(\core_1.execute.sreg_priv_control.o_d[6] ));
 sky130_fd_sc_hd__dfxtp_1 _6842_ (.CLK(clknet_leaf_35_i_clk),
    .D(_0073_),
    .Q(\core_1.execute.sreg_priv_control.o_d[7] ));
 sky130_fd_sc_hd__dfxtp_1 _6843_ (.CLK(clknet_leaf_35_i_clk),
    .D(_0074_),
    .Q(\core_1.execute.sreg_priv_control.o_d[8] ));
 sky130_fd_sc_hd__dfxtp_1 _6844_ (.CLK(clknet_leaf_27_i_clk),
    .D(_0075_),
    .Q(\core_1.execute.sreg_priv_control.o_d[9] ));
 sky130_fd_sc_hd__dfxtp_1 _6845_ (.CLK(clknet_leaf_27_i_clk),
    .D(_0076_),
    .Q(\core_1.execute.sreg_priv_control.o_d[10] ));
 sky130_fd_sc_hd__dfxtp_1 _6846_ (.CLK(clknet_leaf_25_i_clk),
    .D(_0077_),
    .Q(\core_1.execute.sreg_priv_control.o_d[11] ));
 sky130_fd_sc_hd__dfxtp_1 _6847_ (.CLK(clknet_leaf_29_i_clk),
    .D(_0078_),
    .Q(\core_1.execute.sreg_priv_control.o_d[12] ));
 sky130_fd_sc_hd__dfxtp_1 _6848_ (.CLK(clknet_leaf_28_i_clk),
    .D(_0079_),
    .Q(\core_1.execute.sreg_priv_control.o_d[13] ));
 sky130_fd_sc_hd__dfxtp_1 _6849_ (.CLK(clknet_leaf_25_i_clk),
    .D(_0080_),
    .Q(\core_1.execute.sreg_priv_control.o_d[14] ));
 sky130_fd_sc_hd__dfxtp_1 _6850_ (.CLK(clknet_leaf_28_i_clk),
    .D(_0081_),
    .Q(\core_1.execute.sreg_priv_control.o_d[15] ));
 sky130_fd_sc_hd__dfxtp_2 _6851_ (.CLK(clknet_leaf_3_i_clk),
    .D(_0082_),
    .Q(\core_1.execute.alu_mul_div.comp ));
 sky130_fd_sc_hd__dfxtp_1 _6852_ (.CLK(clknet_leaf_39_i_clk),
    .D(_0083_),
    .Q(\core_1.fetch.out_buffer_data_instr[0] ));
 sky130_fd_sc_hd__dfxtp_1 _6853_ (.CLK(clknet_leaf_39_i_clk),
    .D(_0084_),
    .Q(\core_1.fetch.out_buffer_data_instr[1] ));
 sky130_fd_sc_hd__dfxtp_1 _6854_ (.CLK(clknet_leaf_39_i_clk),
    .D(_0085_),
    .Q(\core_1.fetch.out_buffer_data_instr[2] ));
 sky130_fd_sc_hd__dfxtp_1 _6855_ (.CLK(clknet_leaf_37_i_clk),
    .D(_0086_),
    .Q(\core_1.fetch.out_buffer_data_instr[3] ));
 sky130_fd_sc_hd__dfxtp_1 _6856_ (.CLK(clknet_leaf_36_i_clk),
    .D(_0087_),
    .Q(\core_1.fetch.out_buffer_data_instr[4] ));
 sky130_fd_sc_hd__dfxtp_1 _6857_ (.CLK(clknet_leaf_36_i_clk),
    .D(_0088_),
    .Q(\core_1.fetch.out_buffer_data_instr[5] ));
 sky130_fd_sc_hd__dfxtp_1 _6858_ (.CLK(clknet_leaf_36_i_clk),
    .D(_0089_),
    .Q(\core_1.fetch.out_buffer_data_instr[6] ));
 sky130_fd_sc_hd__dfxtp_1 _6859_ (.CLK(clknet_leaf_36_i_clk),
    .D(_0090_),
    .Q(\core_1.fetch.out_buffer_data_instr[7] ));
 sky130_fd_sc_hd__dfxtp_1 _6860_ (.CLK(clknet_leaf_26_i_clk),
    .D(_0091_),
    .Q(\core_1.fetch.out_buffer_data_instr[8] ));
 sky130_fd_sc_hd__dfxtp_1 _6861_ (.CLK(clknet_leaf_25_i_clk),
    .D(_0092_),
    .Q(\core_1.fetch.out_buffer_data_instr[9] ));
 sky130_fd_sc_hd__dfxtp_1 _6862_ (.CLK(clknet_leaf_26_i_clk),
    .D(_0093_),
    .Q(\core_1.fetch.out_buffer_data_instr[10] ));
 sky130_fd_sc_hd__dfxtp_1 _6863_ (.CLK(clknet_leaf_16_i_clk),
    .D(_0094_),
    .Q(\core_1.fetch.out_buffer_data_instr[11] ));
 sky130_fd_sc_hd__dfxtp_1 _6864_ (.CLK(clknet_leaf_16_i_clk),
    .D(_0095_),
    .Q(\core_1.fetch.out_buffer_data_instr[12] ));
 sky130_fd_sc_hd__dfxtp_1 _6865_ (.CLK(clknet_leaf_17_i_clk),
    .D(_0096_),
    .Q(\core_1.fetch.out_buffer_data_instr[13] ));
 sky130_fd_sc_hd__dfxtp_1 _6866_ (.CLK(clknet_leaf_17_i_clk),
    .D(_0097_),
    .Q(\core_1.fetch.out_buffer_data_instr[14] ));
 sky130_fd_sc_hd__dfxtp_1 _6867_ (.CLK(clknet_leaf_20_i_clk),
    .D(_0098_),
    .Q(\core_1.fetch.out_buffer_data_instr[15] ));
 sky130_fd_sc_hd__dfxtp_1 _6868_ (.CLK(clknet_leaf_22_i_clk),
    .D(_0099_),
    .Q(\core_1.fetch.out_buffer_data_instr[16] ));
 sky130_fd_sc_hd__dfxtp_1 _6869_ (.CLK(clknet_leaf_24_i_clk),
    .D(_0100_),
    .Q(\core_1.fetch.out_buffer_data_instr[17] ));
 sky130_fd_sc_hd__dfxtp_1 _6870_ (.CLK(clknet_leaf_23_i_clk),
    .D(_0101_),
    .Q(\core_1.fetch.out_buffer_data_instr[18] ));
 sky130_fd_sc_hd__dfxtp_1 _6871_ (.CLK(clknet_leaf_23_i_clk),
    .D(_0102_),
    .Q(\core_1.fetch.out_buffer_data_instr[19] ));
 sky130_fd_sc_hd__dfxtp_1 _6872_ (.CLK(clknet_leaf_24_i_clk),
    .D(_0103_),
    .Q(\core_1.fetch.out_buffer_data_instr[20] ));
 sky130_fd_sc_hd__dfxtp_1 _6873_ (.CLK(clknet_leaf_23_i_clk),
    .D(_0104_),
    .Q(\core_1.fetch.out_buffer_data_instr[21] ));
 sky130_fd_sc_hd__dfxtp_1 _6874_ (.CLK(clknet_leaf_24_i_clk),
    .D(_0105_),
    .Q(\core_1.fetch.out_buffer_data_instr[22] ));
 sky130_fd_sc_hd__dfxtp_1 _6875_ (.CLK(clknet_leaf_23_i_clk),
    .D(_0106_),
    .Q(\core_1.fetch.out_buffer_data_instr[23] ));
 sky130_fd_sc_hd__dfxtp_1 _6876_ (.CLK(clknet_leaf_23_i_clk),
    .D(_0107_),
    .Q(\core_1.fetch.out_buffer_data_instr[24] ));
 sky130_fd_sc_hd__dfxtp_1 _6877_ (.CLK(clknet_leaf_23_i_clk),
    .D(_0108_),
    .Q(\core_1.fetch.out_buffer_data_instr[25] ));
 sky130_fd_sc_hd__dfxtp_1 _6878_ (.CLK(clknet_leaf_23_i_clk),
    .D(_0109_),
    .Q(\core_1.fetch.out_buffer_data_instr[26] ));
 sky130_fd_sc_hd__dfxtp_1 _6879_ (.CLK(clknet_leaf_23_i_clk),
    .D(_0110_),
    .Q(\core_1.fetch.out_buffer_data_instr[27] ));
 sky130_fd_sc_hd__dfxtp_1 _6880_ (.CLK(clknet_leaf_23_i_clk),
    .D(_0111_),
    .Q(\core_1.fetch.out_buffer_data_instr[28] ));
 sky130_fd_sc_hd__dfxtp_1 _6881_ (.CLK(clknet_leaf_23_i_clk),
    .D(_0112_),
    .Q(\core_1.fetch.out_buffer_data_instr[29] ));
 sky130_fd_sc_hd__dfxtp_1 _6882_ (.CLK(clknet_leaf_23_i_clk),
    .D(_0113_),
    .Q(\core_1.fetch.out_buffer_data_instr[30] ));
 sky130_fd_sc_hd__dfxtp_1 _6883_ (.CLK(clknet_leaf_23_i_clk),
    .D(_0114_),
    .Q(\core_1.fetch.out_buffer_data_instr[31] ));
 sky130_fd_sc_hd__dfxtp_4 _6884_ (.CLK(clknet_leaf_20_i_clk),
    .D(_0115_),
    .Q(\core_1.fetch.out_buffer_valid ));
 sky130_fd_sc_hd__dfxtp_1 _6885_ (.CLK(clknet_leaf_16_i_clk),
    .D(\core_1.fetch.current_req_branch_pred ),
    .Q(\core_1.fetch.prev_req_branch_pred ));
 sky130_fd_sc_hd__dfxtp_1 _6886_ (.CLK(clknet_leaf_21_i_clk),
    .D(_0116_),
    .Q(\core_1.fetch.prev_request_pc[0] ));
 sky130_fd_sc_hd__dfxtp_1 _6887_ (.CLK(clknet_leaf_21_i_clk),
    .D(_0117_),
    .Q(\core_1.fetch.prev_request_pc[1] ));
 sky130_fd_sc_hd__dfxtp_1 _6888_ (.CLK(clknet_leaf_21_i_clk),
    .D(_0118_),
    .Q(\core_1.fetch.prev_request_pc[2] ));
 sky130_fd_sc_hd__dfxtp_1 _6889_ (.CLK(clknet_leaf_21_i_clk),
    .D(_0119_),
    .Q(\core_1.fetch.prev_request_pc[3] ));
 sky130_fd_sc_hd__dfxtp_1 _6890_ (.CLK(clknet_leaf_22_i_clk),
    .D(_0120_),
    .Q(\core_1.fetch.prev_request_pc[4] ));
 sky130_fd_sc_hd__dfxtp_1 _6891_ (.CLK(clknet_leaf_25_i_clk),
    .D(_0121_),
    .Q(\core_1.fetch.prev_request_pc[5] ));
 sky130_fd_sc_hd__dfxtp_1 _6892_ (.CLK(clknet_leaf_22_i_clk),
    .D(_0122_),
    .Q(\core_1.fetch.prev_request_pc[6] ));
 sky130_fd_sc_hd__dfxtp_1 _6893_ (.CLK(clknet_leaf_22_i_clk),
    .D(_0123_),
    .Q(\core_1.fetch.prev_request_pc[7] ));
 sky130_fd_sc_hd__dfxtp_2 _6894_ (.CLK(clknet_leaf_24_i_clk),
    .D(_0124_),
    .Q(\core_1.fetch.prev_request_pc[8] ));
 sky130_fd_sc_hd__dfxtp_1 _6895_ (.CLK(clknet_leaf_24_i_clk),
    .D(_0125_),
    .Q(\core_1.fetch.prev_request_pc[9] ));
 sky130_fd_sc_hd__dfxtp_1 _6896_ (.CLK(clknet_leaf_24_i_clk),
    .D(_0126_),
    .Q(\core_1.fetch.prev_request_pc[10] ));
 sky130_fd_sc_hd__dfxtp_1 _6897_ (.CLK(clknet_leaf_24_i_clk),
    .D(_0127_),
    .Q(\core_1.fetch.prev_request_pc[11] ));
 sky130_fd_sc_hd__dfxtp_1 _6898_ (.CLK(clknet_leaf_24_i_clk),
    .D(_0128_),
    .Q(\core_1.fetch.prev_request_pc[12] ));
 sky130_fd_sc_hd__dfxtp_1 _6899_ (.CLK(clknet_leaf_24_i_clk),
    .D(_0129_),
    .Q(\core_1.fetch.prev_request_pc[13] ));
 sky130_fd_sc_hd__dfxtp_1 _6900_ (.CLK(clknet_leaf_24_i_clk),
    .D(_0130_),
    .Q(\core_1.fetch.prev_request_pc[14] ));
 sky130_fd_sc_hd__dfxtp_1 _6901_ (.CLK(clknet_leaf_24_i_clk),
    .D(_0131_),
    .Q(\core_1.fetch.prev_request_pc[15] ));
 sky130_fd_sc_hd__dfxtp_1 _6902_ (.CLK(clknet_leaf_32_i_clk),
    .D(\core_1.fetch.submitable ),
    .Q(\core_1.decode.i_submit ));
 sky130_fd_sc_hd__dfxtp_1 _6903_ (.CLK(clknet_leaf_17_i_clk),
    .D(_0132_),
    .Q(\core_1.fetch.out_buffer_data_pred ));
 sky130_fd_sc_hd__dfxtp_4 _6904_ (.CLK(clknet_leaf_42_i_clk),
    .D(_0133_),
    .Q(\core_1.decode.i_instr_l[0] ));
 sky130_fd_sc_hd__dfxtp_2 _6905_ (.CLK(clknet_leaf_42_i_clk),
    .D(_0134_),
    .Q(\core_1.decode.i_instr_l[1] ));
 sky130_fd_sc_hd__dfxtp_1 _6906_ (.CLK(clknet_leaf_43_i_clk),
    .D(_0135_),
    .Q(\core_1.decode.i_instr_l[2] ));
 sky130_fd_sc_hd__dfxtp_1 _6907_ (.CLK(clknet_leaf_43_i_clk),
    .D(_0136_),
    .Q(\core_1.decode.i_instr_l[3] ));
 sky130_fd_sc_hd__dfxtp_1 _6908_ (.CLK(clknet_leaf_42_i_clk),
    .D(_0137_),
    .Q(\core_1.decode.i_instr_l[4] ));
 sky130_fd_sc_hd__dfxtp_1 _6909_ (.CLK(clknet_leaf_42_i_clk),
    .D(_0138_),
    .Q(\core_1.decode.i_instr_l[5] ));
 sky130_fd_sc_hd__dfxtp_1 _6910_ (.CLK(clknet_leaf_42_i_clk),
    .D(_0139_),
    .Q(\core_1.decode.i_instr_l[6] ));
 sky130_fd_sc_hd__dfxtp_1 _6911_ (.CLK(clknet_leaf_47_i_clk),
    .D(_0140_),
    .Q(\core_1.decode.i_instr_l[7] ));
 sky130_fd_sc_hd__dfxtp_1 _6912_ (.CLK(clknet_leaf_46_i_clk),
    .D(_0141_),
    .Q(\core_1.decode.i_instr_l[8] ));
 sky130_fd_sc_hd__dfxtp_1 _6913_ (.CLK(clknet_leaf_46_i_clk),
    .D(_0142_),
    .Q(\core_1.decode.i_instr_l[9] ));
 sky130_fd_sc_hd__dfxtp_2 _6914_ (.CLK(clknet_leaf_16_i_clk),
    .D(_0143_),
    .Q(\core_1.decode.i_instr_l[10] ));
 sky130_fd_sc_hd__dfxtp_1 _6915_ (.CLK(clknet_leaf_16_i_clk),
    .D(_0144_),
    .Q(\core_1.decode.i_instr_l[11] ));
 sky130_fd_sc_hd__dfxtp_1 _6916_ (.CLK(clknet_leaf_16_i_clk),
    .D(_0145_),
    .Q(\core_1.decode.i_instr_l[12] ));
 sky130_fd_sc_hd__dfxtp_2 _6917_ (.CLK(clknet_leaf_17_i_clk),
    .D(_0146_),
    .Q(\core_1.decode.i_instr_l[13] ));
 sky130_fd_sc_hd__dfxtp_2 _6918_ (.CLK(clknet_leaf_17_i_clk),
    .D(_0147_),
    .Q(\core_1.decode.i_instr_l[14] ));
 sky130_fd_sc_hd__dfxtp_2 _6919_ (.CLK(clknet_leaf_21_i_clk),
    .D(_0148_),
    .Q(\core_1.decode.i_instr_l[15] ));
 sky130_fd_sc_hd__dfxtp_4 _6920_ (.CLK(clknet_leaf_21_i_clk),
    .D(_0149_),
    .Q(\core_1.decode.i_imm_pass[0] ));
 sky130_fd_sc_hd__dfxtp_4 _6921_ (.CLK(clknet_leaf_21_i_clk),
    .D(_0150_),
    .Q(\core_1.decode.i_imm_pass[1] ));
 sky130_fd_sc_hd__dfxtp_4 _6922_ (.CLK(clknet_leaf_21_i_clk),
    .D(_0151_),
    .Q(\core_1.decode.i_imm_pass[2] ));
 sky130_fd_sc_hd__dfxtp_2 _6923_ (.CLK(clknet_leaf_17_i_clk),
    .D(_0152_),
    .Q(\core_1.decode.i_imm_pass[3] ));
 sky130_fd_sc_hd__dfxtp_1 _6924_ (.CLK(clknet_leaf_20_i_clk),
    .D(_0153_),
    .Q(\core_1.decode.i_imm_pass[4] ));
 sky130_fd_sc_hd__dfxtp_1 _6925_ (.CLK(clknet_leaf_20_i_clk),
    .D(_0154_),
    .Q(\core_1.decode.i_imm_pass[5] ));
 sky130_fd_sc_hd__dfxtp_1 _6926_ (.CLK(clknet_leaf_22_i_clk),
    .D(_0155_),
    .Q(\core_1.decode.i_imm_pass[6] ));
 sky130_fd_sc_hd__dfxtp_1 _6927_ (.CLK(clknet_leaf_20_i_clk),
    .D(_0156_),
    .Q(\core_1.decode.i_imm_pass[7] ));
 sky130_fd_sc_hd__dfxtp_1 _6928_ (.CLK(clknet_leaf_20_i_clk),
    .D(_0157_),
    .Q(\core_1.decode.i_imm_pass[8] ));
 sky130_fd_sc_hd__dfxtp_1 _6929_ (.CLK(clknet_leaf_22_i_clk),
    .D(_0158_),
    .Q(\core_1.decode.i_imm_pass[9] ));
 sky130_fd_sc_hd__dfxtp_1 _6930_ (.CLK(clknet_leaf_20_i_clk),
    .D(_0159_),
    .Q(\core_1.decode.i_imm_pass[10] ));
 sky130_fd_sc_hd__dfxtp_1 _6931_ (.CLK(clknet_leaf_22_i_clk),
    .D(_0160_),
    .Q(\core_1.decode.i_imm_pass[11] ));
 sky130_fd_sc_hd__dfxtp_1 _6932_ (.CLK(clknet_leaf_20_i_clk),
    .D(_0161_),
    .Q(\core_1.decode.i_imm_pass[12] ));
 sky130_fd_sc_hd__dfxtp_1 _6933_ (.CLK(clknet_leaf_23_i_clk),
    .D(_0162_),
    .Q(\core_1.decode.i_imm_pass[13] ));
 sky130_fd_sc_hd__dfxtp_1 _6934_ (.CLK(clknet_leaf_19_i_clk),
    .D(_0163_),
    .Q(\core_1.decode.i_imm_pass[14] ));
 sky130_fd_sc_hd__dfxtp_1 _6935_ (.CLK(clknet_leaf_19_i_clk),
    .D(_0164_),
    .Q(\core_1.decode.i_imm_pass[15] ));
 sky130_fd_sc_hd__dfxtp_1 _6936_ (.CLK(clknet_leaf_21_i_clk),
    .D(_0165_),
    .Q(\core_1.fetch.dbg_out ));
 sky130_fd_sc_hd__dfxtp_1 _6937_ (.CLK(clknet_leaf_17_i_clk),
    .D(_0166_),
    .Q(\core_1.fetch.flush_event_invalidate ));
 sky130_fd_sc_hd__dfxtp_1 _6938_ (.CLK(clknet_leaf_21_i_clk),
    .D(_0167_),
    .Q(\core_1.fetch.pc_flush_override ));
 sky130_fd_sc_hd__dfxtp_1 _6939_ (.CLK(clknet_leaf_17_i_clk),
    .D(_0168_),
    .Q(\core_1.fetch.pc_reset_override ));
 sky130_fd_sc_hd__dfxtp_2 _6940_ (.CLK(clknet_leaf_32_i_clk),
    .D(_0169_),
    .Q(net156));
 sky130_fd_sc_hd__dfxtp_1 _6941_ (.CLK(clknet_leaf_32_i_clk),
    .D(_0170_),
    .Q(\core_1.decode.i_jmp_pred_pass ));
 sky130_fd_sc_hd__dfxtp_1 _6942_ (.CLK(clknet_leaf_43_i_clk),
    .D(_0004_),
    .Q(\core_1.decode.oc_alu_mode[1] ));
 sky130_fd_sc_hd__dfxtp_4 _6943_ (.CLK(clknet_leaf_45_i_clk),
    .D(_0005_),
    .Q(\core_1.decode.oc_alu_mode[2] ));
 sky130_fd_sc_hd__dfxtp_2 _6944_ (.CLK(clknet_leaf_45_i_clk),
    .D(_0006_),
    .Q(\core_1.decode.oc_alu_mode[3] ));
 sky130_fd_sc_hd__dfxtp_1 _6945_ (.CLK(clknet_leaf_48_i_clk),
    .D(_0007_),
    .Q(\core_1.decode.oc_alu_mode[4] ));
 sky130_fd_sc_hd__dfxtp_4 _6946_ (.CLK(clknet_leaf_45_i_clk),
    .D(_0008_),
    .Q(\core_1.execute.alu_mul_div.i_div ));
 sky130_fd_sc_hd__dfxtp_4 _6947_ (.CLK(clknet_leaf_48_i_clk),
    .D(_0009_),
    .Q(\core_1.decode.oc_alu_mode[6] ));
 sky130_fd_sc_hd__dfxtp_4 _6948_ (.CLK(clknet_leaf_45_i_clk),
    .D(_0010_),
    .Q(\core_1.decode.oc_alu_mode[7] ));
 sky130_fd_sc_hd__dfxtp_1 _6949_ (.CLK(clknet_leaf_49_i_clk),
    .D(_0011_),
    .Q(\core_1.execute.alu_mul_div.i_mul ));
 sky130_fd_sc_hd__dfxtp_4 _6950_ (.CLK(clknet_leaf_44_i_clk),
    .D(_0012_),
    .Q(\core_1.decode.oc_alu_mode[9] ));
 sky130_fd_sc_hd__dfxtp_4 _6951_ (.CLK(clknet_leaf_47_i_clk),
    .D(_0000_),
    .Q(\core_1.execute.alu_mul_div.i_mod ));
 sky130_fd_sc_hd__dfxtp_1 _6952_ (.CLK(clknet_leaf_44_i_clk),
    .D(_0001_),
    .Q(\core_1.decode.oc_alu_mode[11] ));
 sky130_fd_sc_hd__dfxtp_4 _6953_ (.CLK(clknet_leaf_44_i_clk),
    .D(_0002_),
    .Q(\core_1.decode.oc_alu_mode[12] ));
 sky130_fd_sc_hd__dfxtp_1 _6954_ (.CLK(clknet_leaf_44_i_clk),
    .D(_0003_),
    .Q(\core_1.decode.oc_alu_mode[13] ));
 sky130_fd_sc_hd__dfxtp_1 _6955_ (.CLK(clknet_leaf_3_i_clk),
    .D(_0171_),
    .Q(\core_1.execute.alu_mul_div.div_cur[1] ));
 sky130_fd_sc_hd__dfxtp_1 _6956_ (.CLK(clknet_leaf_3_i_clk),
    .D(_0172_),
    .Q(\core_1.execute.alu_mul_div.div_cur[2] ));
 sky130_fd_sc_hd__dfxtp_1 _6957_ (.CLK(clknet_leaf_3_i_clk),
    .D(_0173_),
    .Q(\core_1.execute.alu_mul_div.div_cur[3] ));
 sky130_fd_sc_hd__dfxtp_1 _6958_ (.CLK(clknet_leaf_3_i_clk),
    .D(_0174_),
    .Q(\core_1.execute.alu_mul_div.div_cur[4] ));
 sky130_fd_sc_hd__dfxtp_1 _6959_ (.CLK(clknet_leaf_7_i_clk),
    .D(_0175_),
    .Q(\core_1.execute.alu_mul_div.div_cur[5] ));
 sky130_fd_sc_hd__dfxtp_1 _6960_ (.CLK(clknet_leaf_7_i_clk),
    .D(_0176_),
    .Q(\core_1.execute.alu_mul_div.div_cur[6] ));
 sky130_fd_sc_hd__dfxtp_2 _6961_ (.CLK(clknet_leaf_7_i_clk),
    .D(_0177_),
    .Q(\core_1.execute.alu_mul_div.div_cur[7] ));
 sky130_fd_sc_hd__dfxtp_2 _6962_ (.CLK(clknet_leaf_7_i_clk),
    .D(_0178_),
    .Q(\core_1.execute.alu_mul_div.div_cur[8] ));
 sky130_fd_sc_hd__dfxtp_1 _6963_ (.CLK(clknet_leaf_7_i_clk),
    .D(_0179_),
    .Q(\core_1.execute.alu_mul_div.div_cur[9] ));
 sky130_fd_sc_hd__dfxtp_2 _6964_ (.CLK(clknet_leaf_7_i_clk),
    .D(_0180_),
    .Q(\core_1.execute.alu_mul_div.div_cur[10] ));
 sky130_fd_sc_hd__dfxtp_1 _6965_ (.CLK(clknet_leaf_7_i_clk),
    .D(_0181_),
    .Q(\core_1.execute.alu_mul_div.div_cur[11] ));
 sky130_fd_sc_hd__dfxtp_1 _6966_ (.CLK(clknet_leaf_7_i_clk),
    .D(_0182_),
    .Q(\core_1.execute.alu_mul_div.div_cur[12] ));
 sky130_fd_sc_hd__dfxtp_1 _6967_ (.CLK(clknet_leaf_4_i_clk),
    .D(_0183_),
    .Q(\core_1.execute.alu_mul_div.div_cur[13] ));
 sky130_fd_sc_hd__dfxtp_1 _6968_ (.CLK(clknet_leaf_4_i_clk),
    .D(_0184_),
    .Q(\core_1.execute.alu_mul_div.div_cur[14] ));
 sky130_fd_sc_hd__dfxtp_1 _6969_ (.CLK(clknet_leaf_3_i_clk),
    .D(_0185_),
    .Q(\core_1.execute.alu_mul_div.div_cur[15] ));
 sky130_fd_sc_hd__dfxtp_1 _6970_ (.CLK(clknet_leaf_2_i_clk),
    .D(_0186_),
    .Q(\core_1.execute.alu_mul_div.div_cur[0] ));
 sky130_fd_sc_hd__dfxtp_4 _6971_ (.CLK(clknet_leaf_34_i_clk),
    .D(_0187_),
    .Q(net79));
 sky130_fd_sc_hd__dfxtp_2 _6972_ (.CLK(clknet_leaf_0_i_clk),
    .D(_0188_),
    .Q(\core_1.execute.alu_mul_div.cbit[1] ));
 sky130_fd_sc_hd__dfxtp_2 _6973_ (.CLK(clknet_leaf_1_i_clk),
    .D(_0189_),
    .Q(\core_1.execute.alu_mul_div.cbit[2] ));
 sky130_fd_sc_hd__dfxtp_2 _6974_ (.CLK(clknet_leaf_1_i_clk),
    .D(_0190_),
    .Q(\core_1.execute.alu_mul_div.cbit[3] ));
 sky130_fd_sc_hd__dfxtp_1 _6975_ (.CLK(clknet_leaf_46_i_clk),
    .D(_0191_),
    .Q(\core_1.de_jmp_pred ));
 sky130_fd_sc_hd__dfxtp_1 _6976_ (.CLK(clknet_leaf_39_i_clk),
    .D(_0192_),
    .Q(net104));
 sky130_fd_sc_hd__dfxtp_1 _6977_ (.CLK(clknet_leaf_40_i_clk),
    .D(_0014_),
    .Q(net107));
 sky130_fd_sc_hd__dfxtp_1 _6978_ (.CLK(clknet_leaf_33_i_clk),
    .D(_0193_),
    .Q(\core_1.execute.mem_stage_pc[0] ));
 sky130_fd_sc_hd__dfxtp_1 _6979_ (.CLK(clknet_leaf_33_i_clk),
    .D(_0194_),
    .Q(\core_1.execute.mem_stage_pc[1] ));
 sky130_fd_sc_hd__dfxtp_1 _6980_ (.CLK(clknet_leaf_32_i_clk),
    .D(_0195_),
    .Q(\core_1.execute.mem_stage_pc[2] ));
 sky130_fd_sc_hd__dfxtp_1 _6981_ (.CLK(clknet_leaf_34_i_clk),
    .D(_0196_),
    .Q(\core_1.execute.mem_stage_pc[3] ));
 sky130_fd_sc_hd__dfxtp_1 _6982_ (.CLK(clknet_leaf_35_i_clk),
    .D(_0197_),
    .Q(\core_1.execute.mem_stage_pc[4] ));
 sky130_fd_sc_hd__dfxtp_1 _6983_ (.CLK(clknet_leaf_32_i_clk),
    .D(_0198_),
    .Q(\core_1.execute.mem_stage_pc[5] ));
 sky130_fd_sc_hd__dfxtp_1 _6984_ (.CLK(clknet_leaf_33_i_clk),
    .D(_0199_),
    .Q(\core_1.execute.mem_stage_pc[6] ));
 sky130_fd_sc_hd__dfxtp_1 _6985_ (.CLK(clknet_leaf_32_i_clk),
    .D(_0200_),
    .Q(\core_1.execute.mem_stage_pc[7] ));
 sky130_fd_sc_hd__dfxtp_1 _6986_ (.CLK(clknet_leaf_30_i_clk),
    .D(_0201_),
    .Q(\core_1.execute.mem_stage_pc[8] ));
 sky130_fd_sc_hd__dfxtp_1 _6987_ (.CLK(clknet_leaf_30_i_clk),
    .D(_0202_),
    .Q(\core_1.execute.mem_stage_pc[9] ));
 sky130_fd_sc_hd__dfxtp_1 _6988_ (.CLK(clknet_leaf_30_i_clk),
    .D(_0203_),
    .Q(\core_1.execute.mem_stage_pc[10] ));
 sky130_fd_sc_hd__dfxtp_1 _6989_ (.CLK(clknet_leaf_30_i_clk),
    .D(_0204_),
    .Q(\core_1.execute.mem_stage_pc[11] ));
 sky130_fd_sc_hd__dfxtp_1 _6990_ (.CLK(clknet_leaf_29_i_clk),
    .D(_0205_),
    .Q(\core_1.execute.mem_stage_pc[12] ));
 sky130_fd_sc_hd__dfxtp_1 _6991_ (.CLK(clknet_leaf_29_i_clk),
    .D(_0206_),
    .Q(\core_1.execute.mem_stage_pc[13] ));
 sky130_fd_sc_hd__dfxtp_1 _6992_ (.CLK(clknet_leaf_30_i_clk),
    .D(_0207_),
    .Q(\core_1.execute.mem_stage_pc[14] ));
 sky130_fd_sc_hd__dfxtp_1 _6993_ (.CLK(clknet_leaf_30_i_clk),
    .D(_0208_),
    .Q(\core_1.execute.mem_stage_pc[15] ));
 sky130_fd_sc_hd__dfxtp_1 _6994_ (.CLK(clknet_leaf_39_i_clk),
    .D(_0209_),
    .Q(\core_1.execute.prev_pc_high[0] ));
 sky130_fd_sc_hd__dfxtp_1 _6995_ (.CLK(clknet_leaf_40_i_clk),
    .D(_0210_),
    .Q(\core_1.execute.prev_pc_high[1] ));
 sky130_fd_sc_hd__dfxtp_1 _6996_ (.CLK(clknet_leaf_40_i_clk),
    .D(_0211_),
    .Q(\core_1.execute.prev_pc_high[2] ));
 sky130_fd_sc_hd__dfxtp_1 _6997_ (.CLK(clknet_leaf_40_i_clk),
    .D(_0212_),
    .Q(\core_1.execute.prev_pc_high[3] ));
 sky130_fd_sc_hd__dfxtp_1 _6998_ (.CLK(clknet_leaf_40_i_clk),
    .D(_0213_),
    .Q(\core_1.execute.prev_pc_high[4] ));
 sky130_fd_sc_hd__dfxtp_1 _6999_ (.CLK(clknet_leaf_39_i_clk),
    .D(_0214_),
    .Q(\core_1.execute.prev_pc_high[5] ));
 sky130_fd_sc_hd__dfxtp_1 _7000_ (.CLK(clknet_leaf_40_i_clk),
    .D(_0215_),
    .Q(\core_1.execute.prev_pc_high[6] ));
 sky130_fd_sc_hd__dfxtp_1 _7001_ (.CLK(clknet_leaf_40_i_clk),
    .D(_0216_),
    .Q(\core_1.execute.prev_pc_high[7] ));
 sky130_fd_sc_hd__dfxtp_1 _7002_ (.CLK(clknet_leaf_41_i_clk),
    .D(_0217_),
    .Q(\core_1.execute.sreg_irq_flags.i_d[2] ));
 sky130_fd_sc_hd__dfxtp_1 _7003_ (.CLK(clknet_leaf_43_i_clk),
    .D(_0218_),
    .Q(\core_1.execute.prev_sys ));
 sky130_fd_sc_hd__dfxtp_1 _7004_ (.CLK(clknet_leaf_42_i_clk),
    .D(_0219_),
    .Q(net159));
 sky130_fd_sc_hd__dfxtp_1 _7005_ (.CLK(clknet_leaf_31_i_clk),
    .D(_0220_),
    .Q(\core_1.ew_addr_high[0] ));
 sky130_fd_sc_hd__dfxtp_2 _7006_ (.CLK(clknet_leaf_47_i_clk),
    .D(_0221_),
    .Q(net132));
 sky130_fd_sc_hd__dfxtp_2 _7007_ (.CLK(clknet_leaf_47_i_clk),
    .D(_0222_),
    .Q(net133));
 sky130_fd_sc_hd__dfxtp_1 _7008_ (.CLK(clknet_leaf_47_i_clk),
    .D(_0223_),
    .Q(net134));
 sky130_fd_sc_hd__dfxtp_1 _7009_ (.CLK(clknet_leaf_47_i_clk),
    .D(_0224_),
    .Q(net135));
 sky130_fd_sc_hd__dfxtp_1 _7010_ (.CLK(clknet_leaf_47_i_clk),
    .D(_0225_),
    .Q(net136));
 sky130_fd_sc_hd__dfxtp_1 _7011_ (.CLK(clknet_leaf_47_i_clk),
    .D(_0226_),
    .Q(net137));
 sky130_fd_sc_hd__dfxtp_1 _7012_ (.CLK(clknet_leaf_47_i_clk),
    .D(_0227_),
    .Q(net138));
 sky130_fd_sc_hd__dfxtp_1 _7013_ (.CLK(clknet_leaf_30_i_clk),
    .D(_0228_),
    .Q(\core_1.ew_submit ));
 sky130_fd_sc_hd__dfxtp_2 _7014_ (.CLK(clknet_leaf_36_i_clk),
    .D(_0229_),
    .Q(\core_1.ew_data[0] ));
 sky130_fd_sc_hd__dfxtp_2 _7015_ (.CLK(clknet_leaf_36_i_clk),
    .D(_0230_),
    .Q(\core_1.ew_data[1] ));
 sky130_fd_sc_hd__dfxtp_2 _7016_ (.CLK(clknet_leaf_37_i_clk),
    .D(_0231_),
    .Q(\core_1.ew_data[2] ));
 sky130_fd_sc_hd__dfxtp_2 _7017_ (.CLK(clknet_leaf_37_i_clk),
    .D(_0232_),
    .Q(\core_1.ew_data[3] ));
 sky130_fd_sc_hd__dfxtp_2 _7018_ (.CLK(clknet_leaf_36_i_clk),
    .D(_0233_),
    .Q(\core_1.ew_data[4] ));
 sky130_fd_sc_hd__dfxtp_2 _7019_ (.CLK(clknet_leaf_36_i_clk),
    .D(_0234_),
    .Q(\core_1.ew_data[5] ));
 sky130_fd_sc_hd__dfxtp_2 _7020_ (.CLK(clknet_leaf_36_i_clk),
    .D(_0235_),
    .Q(\core_1.ew_data[6] ));
 sky130_fd_sc_hd__dfxtp_1 _7021_ (.CLK(clknet_leaf_36_i_clk),
    .D(_0236_),
    .Q(\core_1.ew_data[7] ));
 sky130_fd_sc_hd__dfxtp_1 _7022_ (.CLK(clknet_leaf_27_i_clk),
    .D(_0237_),
    .Q(\core_1.ew_data[8] ));
 sky130_fd_sc_hd__dfxtp_1 _7023_ (.CLK(clknet_leaf_27_i_clk),
    .D(_0238_),
    .Q(\core_1.ew_data[9] ));
 sky130_fd_sc_hd__dfxtp_1 _7024_ (.CLK(clknet_leaf_26_i_clk),
    .D(_0239_),
    .Q(\core_1.ew_data[10] ));
 sky130_fd_sc_hd__dfxtp_1 _7025_ (.CLK(clknet_leaf_26_i_clk),
    .D(_0240_),
    .Q(\core_1.ew_data[11] ));
 sky130_fd_sc_hd__dfxtp_1 _7026_ (.CLK(clknet_leaf_28_i_clk),
    .D(_0241_),
    .Q(\core_1.ew_data[12] ));
 sky130_fd_sc_hd__dfxtp_1 _7027_ (.CLK(clknet_leaf_25_i_clk),
    .D(_0242_),
    .Q(\core_1.ew_data[13] ));
 sky130_fd_sc_hd__dfxtp_1 _7028_ (.CLK(clknet_leaf_25_i_clk),
    .D(_0243_),
    .Q(\core_1.ew_data[14] ));
 sky130_fd_sc_hd__dfxtp_1 _7029_ (.CLK(clknet_leaf_25_i_clk),
    .D(_0244_),
    .Q(\core_1.ew_data[15] ));
 sky130_fd_sc_hd__dfxtp_1 _7030_ (.CLK(clknet_leaf_36_i_clk),
    .D(_0245_),
    .Q(\core_1.ew_addr[0] ));
 sky130_fd_sc_hd__dfxtp_1 _7031_ (.CLK(clknet_leaf_39_i_clk),
    .D(_0246_),
    .Q(net116));
 sky130_fd_sc_hd__dfxtp_1 _7032_ (.CLK(clknet_leaf_39_i_clk),
    .D(_0247_),
    .Q(net123));
 sky130_fd_sc_hd__dfxtp_1 _7033_ (.CLK(clknet_leaf_37_i_clk),
    .D(_0248_),
    .Q(net124));
 sky130_fd_sc_hd__dfxtp_1 _7034_ (.CLK(clknet_leaf_37_i_clk),
    .D(_0249_),
    .Q(net125));
 sky130_fd_sc_hd__dfxtp_1 _7035_ (.CLK(clknet_leaf_36_i_clk),
    .D(_0250_),
    .Q(net126));
 sky130_fd_sc_hd__dfxtp_1 _7036_ (.CLK(clknet_leaf_36_i_clk),
    .D(_0251_),
    .Q(net127));
 sky130_fd_sc_hd__dfxtp_1 _7037_ (.CLK(clknet_leaf_36_i_clk),
    .D(_0252_),
    .Q(net128));
 sky130_fd_sc_hd__dfxtp_1 _7038_ (.CLK(clknet_leaf_36_i_clk),
    .D(_0253_),
    .Q(net129));
 sky130_fd_sc_hd__dfxtp_1 _7039_ (.CLK(clknet_leaf_27_i_clk),
    .D(_0254_),
    .Q(net130));
 sky130_fd_sc_hd__dfxtp_1 _7040_ (.CLK(clknet_leaf_26_i_clk),
    .D(_0255_),
    .Q(net131));
 sky130_fd_sc_hd__dfxtp_1 _7041_ (.CLK(clknet_leaf_26_i_clk),
    .D(_0256_),
    .Q(net117));
 sky130_fd_sc_hd__dfxtp_1 _7042_ (.CLK(clknet_leaf_26_i_clk),
    .D(_0257_),
    .Q(net118));
 sky130_fd_sc_hd__dfxtp_1 _7043_ (.CLK(clknet_leaf_26_i_clk),
    .D(_0258_),
    .Q(net119));
 sky130_fd_sc_hd__dfxtp_1 _7044_ (.CLK(clknet_leaf_24_i_clk),
    .D(_0259_),
    .Q(net120));
 sky130_fd_sc_hd__dfxtp_1 _7045_ (.CLK(clknet_leaf_24_i_clk),
    .D(_0260_),
    .Q(net121));
 sky130_fd_sc_hd__dfxtp_1 _7046_ (.CLK(clknet_leaf_31_i_clk),
    .D(_0261_),
    .Q(\core_1.ew_reg_ie[0] ));
 sky130_fd_sc_hd__dfxtp_2 _7047_ (.CLK(clknet_leaf_47_i_clk),
    .D(_0262_),
    .Q(\core_1.ew_reg_ie[1] ));
 sky130_fd_sc_hd__dfxtp_2 _7048_ (.CLK(clknet_leaf_47_i_clk),
    .D(_0263_),
    .Q(\core_1.ew_reg_ie[2] ));
 sky130_fd_sc_hd__dfxtp_2 _7049_ (.CLK(clknet_leaf_47_i_clk),
    .D(_0264_),
    .Q(\core_1.ew_reg_ie[3] ));
 sky130_fd_sc_hd__dfxtp_2 _7050_ (.CLK(clknet_leaf_31_i_clk),
    .D(_0265_),
    .Q(\core_1.ew_reg_ie[4] ));
 sky130_fd_sc_hd__dfxtp_2 _7051_ (.CLK(clknet_leaf_31_i_clk),
    .D(_0266_),
    .Q(\core_1.ew_reg_ie[5] ));
 sky130_fd_sc_hd__dfxtp_2 _7052_ (.CLK(clknet_leaf_47_i_clk),
    .D(_0267_),
    .Q(\core_1.ew_reg_ie[6] ));
 sky130_fd_sc_hd__dfxtp_2 _7053_ (.CLK(clknet_leaf_47_i_clk),
    .D(_0268_),
    .Q(\core_1.ew_reg_ie[7] ));
 sky130_fd_sc_hd__dfxtp_1 _7054_ (.CLK(clknet_leaf_32_i_clk),
    .D(_0269_),
    .Q(\core_1.ew_mem_access ));
 sky130_fd_sc_hd__dfxtp_2 _7055_ (.CLK(clknet_leaf_46_i_clk),
    .D(_0270_),
    .Q(\core_1.ew_mem_width ));
 sky130_fd_sc_hd__dfxtp_1 _7056_ (.CLK(clknet_leaf_46_i_clk),
    .D(_0013_),
    .Q(\core_1.decode.i_flush ));
 sky130_fd_sc_hd__dfxtp_2 _7057_ (.CLK(clknet_leaf_46_i_clk),
    .D(_0271_),
    .Q(net155));
 sky130_fd_sc_hd__dfxtp_1 _7058_ (.CLK(clknet_leaf_47_i_clk),
    .D(_0272_),
    .Q(\core_1.execute.hold_valid ));
 sky130_fd_sc_hd__dfxtp_1 _7059_ (.CLK(clknet_leaf_4_i_clk),
    .D(_0273_),
    .Q(\core_1.execute.rf.reg_outputs[7][0] ));
 sky130_fd_sc_hd__dfxtp_1 _7060_ (.CLK(clknet_leaf_5_i_clk),
    .D(_0274_),
    .Q(\core_1.execute.rf.reg_outputs[7][1] ));
 sky130_fd_sc_hd__dfxtp_1 _7061_ (.CLK(clknet_leaf_13_i_clk),
    .D(_0275_),
    .Q(\core_1.execute.rf.reg_outputs[7][2] ));
 sky130_fd_sc_hd__dfxtp_1 _7062_ (.CLK(clknet_leaf_6_i_clk),
    .D(_0276_),
    .Q(\core_1.execute.rf.reg_outputs[7][3] ));
 sky130_fd_sc_hd__dfxtp_1 _7063_ (.CLK(clknet_leaf_15_i_clk),
    .D(_0277_),
    .Q(\core_1.execute.rf.reg_outputs[7][4] ));
 sky130_fd_sc_hd__dfxtp_1 _7064_ (.CLK(clknet_leaf_5_i_clk),
    .D(_0278_),
    .Q(\core_1.execute.rf.reg_outputs[7][5] ));
 sky130_fd_sc_hd__dfxtp_1 _7065_ (.CLK(clknet_leaf_5_i_clk),
    .D(_0279_),
    .Q(\core_1.execute.rf.reg_outputs[7][6] ));
 sky130_fd_sc_hd__dfxtp_1 _7066_ (.CLK(clknet_leaf_14_i_clk),
    .D(_0280_),
    .Q(\core_1.execute.rf.reg_outputs[7][7] ));
 sky130_fd_sc_hd__dfxtp_1 _7067_ (.CLK(clknet_leaf_18_i_clk),
    .D(_0281_),
    .Q(\core_1.execute.rf.reg_outputs[7][8] ));
 sky130_fd_sc_hd__dfxtp_1 _7068_ (.CLK(clknet_leaf_9_i_clk),
    .D(_0282_),
    .Q(\core_1.execute.rf.reg_outputs[7][9] ));
 sky130_fd_sc_hd__dfxtp_1 _7069_ (.CLK(clknet_leaf_9_i_clk),
    .D(_0283_),
    .Q(\core_1.execute.rf.reg_outputs[7][10] ));
 sky130_fd_sc_hd__dfxtp_1 _7070_ (.CLK(clknet_leaf_9_i_clk),
    .D(_0284_),
    .Q(\core_1.execute.rf.reg_outputs[7][11] ));
 sky130_fd_sc_hd__dfxtp_1 _7071_ (.CLK(clknet_leaf_11_i_clk),
    .D(_0285_),
    .Q(\core_1.execute.rf.reg_outputs[7][12] ));
 sky130_fd_sc_hd__dfxtp_1 _7072_ (.CLK(clknet_leaf_11_i_clk),
    .D(_0286_),
    .Q(\core_1.execute.rf.reg_outputs[7][13] ));
 sky130_fd_sc_hd__dfxtp_1 _7073_ (.CLK(clknet_leaf_10_i_clk),
    .D(_0287_),
    .Q(\core_1.execute.rf.reg_outputs[7][14] ));
 sky130_fd_sc_hd__dfxtp_1 _7074_ (.CLK(clknet_leaf_13_i_clk),
    .D(_0288_),
    .Q(\core_1.execute.rf.reg_outputs[7][15] ));
 sky130_fd_sc_hd__dfxtp_1 _7075_ (.CLK(clknet_leaf_6_i_clk),
    .D(_0289_),
    .Q(\core_1.execute.rf.reg_outputs[6][0] ));
 sky130_fd_sc_hd__dfxtp_1 _7076_ (.CLK(clknet_leaf_6_i_clk),
    .D(_0290_),
    .Q(\core_1.execute.rf.reg_outputs[6][1] ));
 sky130_fd_sc_hd__dfxtp_1 _7077_ (.CLK(clknet_leaf_6_i_clk),
    .D(_0291_),
    .Q(\core_1.execute.rf.reg_outputs[6][2] ));
 sky130_fd_sc_hd__dfxtp_1 _7078_ (.CLK(clknet_leaf_6_i_clk),
    .D(_0292_),
    .Q(\core_1.execute.rf.reg_outputs[6][3] ));
 sky130_fd_sc_hd__dfxtp_1 _7079_ (.CLK(clknet_leaf_15_i_clk),
    .D(_0293_),
    .Q(\core_1.execute.rf.reg_outputs[6][4] ));
 sky130_fd_sc_hd__dfxtp_1 _7080_ (.CLK(clknet_leaf_14_i_clk),
    .D(_0294_),
    .Q(\core_1.execute.rf.reg_outputs[6][5] ));
 sky130_fd_sc_hd__dfxtp_1 _7081_ (.CLK(clknet_leaf_14_i_clk),
    .D(_0295_),
    .Q(\core_1.execute.rf.reg_outputs[6][6] ));
 sky130_fd_sc_hd__dfxtp_1 _7082_ (.CLK(clknet_leaf_13_i_clk),
    .D(_0296_),
    .Q(\core_1.execute.rf.reg_outputs[6][7] ));
 sky130_fd_sc_hd__dfxtp_1 _7083_ (.CLK(clknet_leaf_11_i_clk),
    .D(_0297_),
    .Q(\core_1.execute.rf.reg_outputs[6][8] ));
 sky130_fd_sc_hd__dfxtp_2 _7084_ (.CLK(clknet_leaf_11_i_clk),
    .D(_0298_),
    .Q(\core_1.execute.rf.reg_outputs[6][9] ));
 sky130_fd_sc_hd__dfxtp_1 _7085_ (.CLK(clknet_leaf_10_i_clk),
    .D(_0299_),
    .Q(\core_1.execute.rf.reg_outputs[6][10] ));
 sky130_fd_sc_hd__dfxtp_1 _7086_ (.CLK(clknet_leaf_10_i_clk),
    .D(_0300_),
    .Q(\core_1.execute.rf.reg_outputs[6][11] ));
 sky130_fd_sc_hd__dfxtp_1 _7087_ (.CLK(clknet_leaf_11_i_clk),
    .D(_0301_),
    .Q(\core_1.execute.rf.reg_outputs[6][12] ));
 sky130_fd_sc_hd__dfxtp_1 _7088_ (.CLK(clknet_leaf_11_i_clk),
    .D(_0302_),
    .Q(\core_1.execute.rf.reg_outputs[6][13] ));
 sky130_fd_sc_hd__dfxtp_1 _7089_ (.CLK(clknet_leaf_10_i_clk),
    .D(_0303_),
    .Q(\core_1.execute.rf.reg_outputs[6][14] ));
 sky130_fd_sc_hd__dfxtp_1 _7090_ (.CLK(clknet_leaf_13_i_clk),
    .D(_0304_),
    .Q(\core_1.execute.rf.reg_outputs[6][15] ));
 sky130_fd_sc_hd__dfxtp_1 _7091_ (.CLK(clknet_leaf_6_i_clk),
    .D(_0305_),
    .Q(\core_1.execute.rf.reg_outputs[5][0] ));
 sky130_fd_sc_hd__dfxtp_1 _7092_ (.CLK(clknet_leaf_6_i_clk),
    .D(_0306_),
    .Q(\core_1.execute.rf.reg_outputs[5][1] ));
 sky130_fd_sc_hd__dfxtp_1 _7093_ (.CLK(clknet_leaf_6_i_clk),
    .D(_0307_),
    .Q(\core_1.execute.rf.reg_outputs[5][2] ));
 sky130_fd_sc_hd__dfxtp_1 _7094_ (.CLK(clknet_leaf_6_i_clk),
    .D(_0308_),
    .Q(\core_1.execute.rf.reg_outputs[5][3] ));
 sky130_fd_sc_hd__dfxtp_1 _7095_ (.CLK(clknet_leaf_15_i_clk),
    .D(_0309_),
    .Q(\core_1.execute.rf.reg_outputs[5][4] ));
 sky130_fd_sc_hd__dfxtp_1 _7096_ (.CLK(clknet_leaf_15_i_clk),
    .D(_0310_),
    .Q(\core_1.execute.rf.reg_outputs[5][5] ));
 sky130_fd_sc_hd__dfxtp_1 _7097_ (.CLK(clknet_leaf_31_i_clk),
    .D(_0311_),
    .Q(\core_1.execute.rf.reg_outputs[5][6] ));
 sky130_fd_sc_hd__dfxtp_1 _7098_ (.CLK(clknet_leaf_14_i_clk),
    .D(_0312_),
    .Q(\core_1.execute.rf.reg_outputs[5][7] ));
 sky130_fd_sc_hd__dfxtp_1 _7099_ (.CLK(clknet_leaf_18_i_clk),
    .D(_0313_),
    .Q(\core_1.execute.rf.reg_outputs[5][8] ));
 sky130_fd_sc_hd__dfxtp_1 _7100_ (.CLK(clknet_leaf_11_i_clk),
    .D(_0314_),
    .Q(\core_1.execute.rf.reg_outputs[5][9] ));
 sky130_fd_sc_hd__dfxtp_1 _7101_ (.CLK(clknet_leaf_10_i_clk),
    .D(_0315_),
    .Q(\core_1.execute.rf.reg_outputs[5][10] ));
 sky130_fd_sc_hd__dfxtp_1 _7102_ (.CLK(clknet_leaf_10_i_clk),
    .D(_0316_),
    .Q(\core_1.execute.rf.reg_outputs[5][11] ));
 sky130_fd_sc_hd__dfxtp_1 _7103_ (.CLK(clknet_leaf_11_i_clk),
    .D(_0317_),
    .Q(\core_1.execute.rf.reg_outputs[5][12] ));
 sky130_fd_sc_hd__dfxtp_1 _7104_ (.CLK(clknet_leaf_11_i_clk),
    .D(_0318_),
    .Q(\core_1.execute.rf.reg_outputs[5][13] ));
 sky130_fd_sc_hd__dfxtp_1 _7105_ (.CLK(clknet_leaf_10_i_clk),
    .D(_0319_),
    .Q(\core_1.execute.rf.reg_outputs[5][14] ));
 sky130_fd_sc_hd__dfxtp_1 _7106_ (.CLK(clknet_leaf_12_i_clk),
    .D(_0320_),
    .Q(\core_1.execute.rf.reg_outputs[5][15] ));
 sky130_fd_sc_hd__dfxtp_1 _7107_ (.CLK(clknet_leaf_6_i_clk),
    .D(_0321_),
    .Q(\core_1.execute.rf.reg_outputs[4][0] ));
 sky130_fd_sc_hd__dfxtp_1 _7108_ (.CLK(clknet_leaf_6_i_clk),
    .D(_0322_),
    .Q(\core_1.execute.rf.reg_outputs[4][1] ));
 sky130_fd_sc_hd__dfxtp_1 _7109_ (.CLK(clknet_leaf_13_i_clk),
    .D(_0323_),
    .Q(\core_1.execute.rf.reg_outputs[4][2] ));
 sky130_fd_sc_hd__dfxtp_1 _7110_ (.CLK(clknet_leaf_6_i_clk),
    .D(_0324_),
    .Q(\core_1.execute.rf.reg_outputs[4][3] ));
 sky130_fd_sc_hd__dfxtp_1 _7111_ (.CLK(clknet_leaf_15_i_clk),
    .D(_0325_),
    .Q(\core_1.execute.rf.reg_outputs[4][4] ));
 sky130_fd_sc_hd__dfxtp_1 _7112_ (.CLK(clknet_leaf_31_i_clk),
    .D(_0326_),
    .Q(\core_1.execute.rf.reg_outputs[4][5] ));
 sky130_fd_sc_hd__dfxtp_1 _7113_ (.CLK(clknet_leaf_16_i_clk),
    .D(_0327_),
    .Q(\core_1.execute.rf.reg_outputs[4][6] ));
 sky130_fd_sc_hd__dfxtp_1 _7114_ (.CLK(clknet_leaf_16_i_clk),
    .D(_0328_),
    .Q(\core_1.execute.rf.reg_outputs[4][7] ));
 sky130_fd_sc_hd__dfxtp_1 _7115_ (.CLK(clknet_leaf_19_i_clk),
    .D(_0329_),
    .Q(\core_1.execute.rf.reg_outputs[4][8] ));
 sky130_fd_sc_hd__dfxtp_1 _7116_ (.CLK(clknet_leaf_10_i_clk),
    .D(_0330_),
    .Q(\core_1.execute.rf.reg_outputs[4][9] ));
 sky130_fd_sc_hd__dfxtp_1 _7117_ (.CLK(clknet_leaf_10_i_clk),
    .D(_0331_),
    .Q(\core_1.execute.rf.reg_outputs[4][10] ));
 sky130_fd_sc_hd__dfxtp_1 _7118_ (.CLK(clknet_leaf_10_i_clk),
    .D(_0332_),
    .Q(\core_1.execute.rf.reg_outputs[4][11] ));
 sky130_fd_sc_hd__dfxtp_1 _7119_ (.CLK(clknet_leaf_19_i_clk),
    .D(_0333_),
    .Q(\core_1.execute.rf.reg_outputs[4][12] ));
 sky130_fd_sc_hd__dfxtp_1 _7120_ (.CLK(clknet_leaf_19_i_clk),
    .D(_0334_),
    .Q(\core_1.execute.rf.reg_outputs[4][13] ));
 sky130_fd_sc_hd__dfxtp_1 _7121_ (.CLK(clknet_leaf_10_i_clk),
    .D(_0335_),
    .Q(\core_1.execute.rf.reg_outputs[4][14] ));
 sky130_fd_sc_hd__dfxtp_1 _7122_ (.CLK(clknet_leaf_10_i_clk),
    .D(_0336_),
    .Q(\core_1.execute.rf.reg_outputs[4][15] ));
 sky130_fd_sc_hd__dfxtp_1 _7123_ (.CLK(clknet_leaf_5_i_clk),
    .D(_0337_),
    .Q(\core_1.execute.rf.reg_outputs[3][0] ));
 sky130_fd_sc_hd__dfxtp_1 _7124_ (.CLK(clknet_leaf_5_i_clk),
    .D(_0338_),
    .Q(\core_1.execute.rf.reg_outputs[3][1] ));
 sky130_fd_sc_hd__dfxtp_1 _7125_ (.CLK(clknet_leaf_6_i_clk),
    .D(_0339_),
    .Q(\core_1.execute.rf.reg_outputs[3][2] ));
 sky130_fd_sc_hd__dfxtp_1 _7126_ (.CLK(clknet_leaf_6_i_clk),
    .D(_0340_),
    .Q(\core_1.execute.rf.reg_outputs[3][3] ));
 sky130_fd_sc_hd__dfxtp_1 _7127_ (.CLK(clknet_leaf_16_i_clk),
    .D(_0341_),
    .Q(\core_1.execute.rf.reg_outputs[3][4] ));
 sky130_fd_sc_hd__dfxtp_1 _7128_ (.CLK(clknet_leaf_5_i_clk),
    .D(_0342_),
    .Q(\core_1.execute.rf.reg_outputs[3][5] ));
 sky130_fd_sc_hd__dfxtp_1 _7129_ (.CLK(clknet_leaf_5_i_clk),
    .D(_0343_),
    .Q(\core_1.execute.rf.reg_outputs[3][6] ));
 sky130_fd_sc_hd__dfxtp_1 _7130_ (.CLK(clknet_leaf_14_i_clk),
    .D(_0344_),
    .Q(\core_1.execute.rf.reg_outputs[3][7] ));
 sky130_fd_sc_hd__dfxtp_1 _7131_ (.CLK(clknet_leaf_12_i_clk),
    .D(_0345_),
    .Q(\core_1.execute.rf.reg_outputs[3][8] ));
 sky130_fd_sc_hd__dfxtp_1 _7132_ (.CLK(clknet_leaf_10_i_clk),
    .D(_0346_),
    .Q(\core_1.execute.rf.reg_outputs[3][9] ));
 sky130_fd_sc_hd__dfxtp_1 _7133_ (.CLK(clknet_leaf_10_i_clk),
    .D(_0347_),
    .Q(\core_1.execute.rf.reg_outputs[3][10] ));
 sky130_fd_sc_hd__dfxtp_1 _7134_ (.CLK(clknet_leaf_10_i_clk),
    .D(_0348_),
    .Q(\core_1.execute.rf.reg_outputs[3][11] ));
 sky130_fd_sc_hd__dfxtp_1 _7135_ (.CLK(clknet_leaf_11_i_clk),
    .D(_0349_),
    .Q(\core_1.execute.rf.reg_outputs[3][12] ));
 sky130_fd_sc_hd__dfxtp_1 _7136_ (.CLK(clknet_leaf_11_i_clk),
    .D(_0350_),
    .Q(\core_1.execute.rf.reg_outputs[3][13] ));
 sky130_fd_sc_hd__dfxtp_1 _7137_ (.CLK(clknet_leaf_9_i_clk),
    .D(_0351_),
    .Q(\core_1.execute.rf.reg_outputs[3][14] ));
 sky130_fd_sc_hd__dfxtp_1 _7138_ (.CLK(clknet_leaf_12_i_clk),
    .D(_0352_),
    .Q(\core_1.execute.rf.reg_outputs[3][15] ));
 sky130_fd_sc_hd__dfxtp_1 _7139_ (.CLK(clknet_leaf_6_i_clk),
    .D(_0353_),
    .Q(\core_1.execute.rf.reg_outputs[2][0] ));
 sky130_fd_sc_hd__dfxtp_1 _7140_ (.CLK(clknet_leaf_6_i_clk),
    .D(_0354_),
    .Q(\core_1.execute.rf.reg_outputs[2][1] ));
 sky130_fd_sc_hd__dfxtp_1 _7141_ (.CLK(clknet_leaf_6_i_clk),
    .D(_0355_),
    .Q(\core_1.execute.rf.reg_outputs[2][2] ));
 sky130_fd_sc_hd__dfxtp_1 _7142_ (.CLK(clknet_leaf_6_i_clk),
    .D(_0356_),
    .Q(\core_1.execute.rf.reg_outputs[2][3] ));
 sky130_fd_sc_hd__dfxtp_1 _7143_ (.CLK(clknet_leaf_15_i_clk),
    .D(_0357_),
    .Q(\core_1.execute.rf.reg_outputs[2][4] ));
 sky130_fd_sc_hd__dfxtp_1 _7144_ (.CLK(clknet_leaf_14_i_clk),
    .D(_0358_),
    .Q(\core_1.execute.rf.reg_outputs[2][5] ));
 sky130_fd_sc_hd__dfxtp_1 _7145_ (.CLK(clknet_leaf_14_i_clk),
    .D(_0359_),
    .Q(\core_1.execute.rf.reg_outputs[2][6] ));
 sky130_fd_sc_hd__dfxtp_1 _7146_ (.CLK(clknet_leaf_13_i_clk),
    .D(_0360_),
    .Q(\core_1.execute.rf.reg_outputs[2][7] ));
 sky130_fd_sc_hd__dfxtp_1 _7147_ (.CLK(clknet_leaf_18_i_clk),
    .D(_0361_),
    .Q(\core_1.execute.rf.reg_outputs[2][8] ));
 sky130_fd_sc_hd__dfxtp_1 _7148_ (.CLK(clknet_leaf_9_i_clk),
    .D(_0362_),
    .Q(\core_1.execute.rf.reg_outputs[2][9] ));
 sky130_fd_sc_hd__dfxtp_1 _7149_ (.CLK(clknet_leaf_9_i_clk),
    .D(_0363_),
    .Q(\core_1.execute.rf.reg_outputs[2][10] ));
 sky130_fd_sc_hd__dfxtp_1 _7150_ (.CLK(clknet_leaf_9_i_clk),
    .D(_0364_),
    .Q(\core_1.execute.rf.reg_outputs[2][11] ));
 sky130_fd_sc_hd__dfxtp_1 _7151_ (.CLK(clknet_leaf_11_i_clk),
    .D(_0365_),
    .Q(\core_1.execute.rf.reg_outputs[2][12] ));
 sky130_fd_sc_hd__dfxtp_1 _7152_ (.CLK(clknet_leaf_19_i_clk),
    .D(_0366_),
    .Q(\core_1.execute.rf.reg_outputs[2][13] ));
 sky130_fd_sc_hd__dfxtp_1 _7153_ (.CLK(clknet_leaf_9_i_clk),
    .D(_0367_),
    .Q(\core_1.execute.rf.reg_outputs[2][14] ));
 sky130_fd_sc_hd__dfxtp_1 _7154_ (.CLK(clknet_leaf_12_i_clk),
    .D(_0368_),
    .Q(\core_1.execute.rf.reg_outputs[2][15] ));
 sky130_fd_sc_hd__dfxtp_1 _7155_ (.CLK(clknet_leaf_5_i_clk),
    .D(_0369_),
    .Q(\core_1.execute.rf.reg_outputs[1][0] ));
 sky130_fd_sc_hd__dfxtp_1 _7156_ (.CLK(clknet_leaf_5_i_clk),
    .D(_0370_),
    .Q(\core_1.execute.rf.reg_outputs[1][1] ));
 sky130_fd_sc_hd__dfxtp_1 _7157_ (.CLK(clknet_leaf_6_i_clk),
    .D(_0371_),
    .Q(\core_1.execute.rf.reg_outputs[1][2] ));
 sky130_fd_sc_hd__dfxtp_2 _7158_ (.CLK(clknet_leaf_4_i_clk),
    .D(_0372_),
    .Q(\core_1.execute.rf.reg_outputs[1][3] ));
 sky130_fd_sc_hd__dfxtp_2 _7159_ (.CLK(clknet_leaf_15_i_clk),
    .D(_0373_),
    .Q(\core_1.execute.rf.reg_outputs[1][4] ));
 sky130_fd_sc_hd__dfxtp_1 _7160_ (.CLK(clknet_leaf_15_i_clk),
    .D(_0374_),
    .Q(\core_1.execute.rf.reg_outputs[1][5] ));
 sky130_fd_sc_hd__dfxtp_2 _7161_ (.CLK(clknet_leaf_16_i_clk),
    .D(_0375_),
    .Q(\core_1.execute.rf.reg_outputs[1][6] ));
 sky130_fd_sc_hd__dfxtp_1 _7162_ (.CLK(clknet_leaf_16_i_clk),
    .D(_0376_),
    .Q(\core_1.execute.rf.reg_outputs[1][7] ));
 sky130_fd_sc_hd__dfxtp_1 _7163_ (.CLK(clknet_leaf_18_i_clk),
    .D(_0377_),
    .Q(\core_1.execute.rf.reg_outputs[1][8] ));
 sky130_fd_sc_hd__dfxtp_1 _7164_ (.CLK(clknet_leaf_18_i_clk),
    .D(_0378_),
    .Q(\core_1.execute.rf.reg_outputs[1][9] ));
 sky130_fd_sc_hd__dfxtp_1 _7165_ (.CLK(clknet_leaf_19_i_clk),
    .D(_0379_),
    .Q(\core_1.execute.rf.reg_outputs[1][10] ));
 sky130_fd_sc_hd__dfxtp_1 _7166_ (.CLK(clknet_leaf_18_i_clk),
    .D(_0380_),
    .Q(\core_1.execute.rf.reg_outputs[1][11] ));
 sky130_fd_sc_hd__dfxtp_1 _7167_ (.CLK(clknet_leaf_18_i_clk),
    .D(_0381_),
    .Q(\core_1.execute.rf.reg_outputs[1][12] ));
 sky130_fd_sc_hd__dfxtp_1 _7168_ (.CLK(clknet_leaf_18_i_clk),
    .D(_0382_),
    .Q(\core_1.execute.rf.reg_outputs[1][13] ));
 sky130_fd_sc_hd__dfxtp_1 _7169_ (.CLK(clknet_leaf_19_i_clk),
    .D(_0383_),
    .Q(\core_1.execute.rf.reg_outputs[1][14] ));
 sky130_fd_sc_hd__dfxtp_1 _7170_ (.CLK(clknet_leaf_18_i_clk),
    .D(_0384_),
    .Q(\core_1.execute.rf.reg_outputs[1][15] ));
 sky130_fd_sc_hd__dfxtp_4 _7171_ (.CLK(clknet_leaf_30_i_clk),
    .D(_0385_),
    .Q(net88));
 sky130_fd_sc_hd__dfxtp_4 _7172_ (.CLK(clknet_leaf_30_i_clk),
    .D(_0386_),
    .Q(net95));
 sky130_fd_sc_hd__dfxtp_4 _7173_ (.CLK(clknet_leaf_16_i_clk),
    .D(_0387_),
    .Q(net96));
 sky130_fd_sc_hd__dfxtp_4 _7174_ (.CLK(clknet_leaf_16_i_clk),
    .D(_0388_),
    .Q(net97));
 sky130_fd_sc_hd__dfxtp_4 _7175_ (.CLK(clknet_leaf_16_i_clk),
    .D(_0389_),
    .Q(net98));
 sky130_fd_sc_hd__dfxtp_2 _7176_ (.CLK(clknet_leaf_30_i_clk),
    .D(_0390_),
    .Q(net99));
 sky130_fd_sc_hd__dfxtp_2 _7177_ (.CLK(clknet_leaf_31_i_clk),
    .D(_0391_),
    .Q(net100));
 sky130_fd_sc_hd__dfxtp_2 _7178_ (.CLK(clknet_leaf_16_i_clk),
    .D(_0392_),
    .Q(net101));
 sky130_fd_sc_hd__dfxtp_4 _7179_ (.CLK(clknet_leaf_17_i_clk),
    .D(_0393_),
    .Q(net102));
 sky130_fd_sc_hd__dfxtp_2 _7180_ (.CLK(clknet_leaf_18_i_clk),
    .D(_0394_),
    .Q(net103));
 sky130_fd_sc_hd__dfxtp_4 _7181_ (.CLK(clknet_leaf_19_i_clk),
    .D(_0395_),
    .Q(net89));
 sky130_fd_sc_hd__dfxtp_4 _7182_ (.CLK(clknet_leaf_17_i_clk),
    .D(_0396_),
    .Q(net90));
 sky130_fd_sc_hd__dfxtp_2 _7183_ (.CLK(clknet_leaf_17_i_clk),
    .D(_0397_),
    .Q(net91));
 sky130_fd_sc_hd__dfxtp_2 _7184_ (.CLK(clknet_leaf_18_i_clk),
    .D(_0398_),
    .Q(net92));
 sky130_fd_sc_hd__dfxtp_4 _7185_ (.CLK(clknet_leaf_18_i_clk),
    .D(_0399_),
    .Q(net93));
 sky130_fd_sc_hd__dfxtp_4 _7186_ (.CLK(clknet_leaf_18_i_clk),
    .D(_0400_),
    .Q(net94));
 sky130_fd_sc_hd__dfxtp_2 _7187_ (.CLK(clknet_leaf_37_i_clk),
    .D(_0401_),
    .Q(\core_1.execute.irq_en ));
 sky130_fd_sc_hd__dfxtp_2 _7188_ (.CLK(clknet_leaf_0_i_clk),
    .D(_0402_),
    .Q(\core_1.execute.alu_mul_div.cbit[0] ));
 sky130_fd_sc_hd__dfxtp_1 _7189_ (.CLK(clknet_leaf_50_i_clk),
    .D(_0403_),
    .Q(\core_1.execute.alu_mul_div.mul_res[0] ));
 sky130_fd_sc_hd__dfxtp_1 _7190_ (.CLK(clknet_leaf_0_i_clk),
    .D(_0404_),
    .Q(\core_1.execute.alu_mul_div.mul_res[1] ));
 sky130_fd_sc_hd__dfxtp_1 _7191_ (.CLK(clknet_leaf_49_i_clk),
    .D(_0405_),
    .Q(\core_1.execute.alu_mul_div.mul_res[2] ));
 sky130_fd_sc_hd__dfxtp_1 _7192_ (.CLK(clknet_leaf_49_i_clk),
    .D(_0406_),
    .Q(\core_1.execute.alu_mul_div.mul_res[3] ));
 sky130_fd_sc_hd__dfxtp_1 _7193_ (.CLK(clknet_leaf_49_i_clk),
    .D(_0407_),
    .Q(\core_1.execute.alu_mul_div.mul_res[4] ));
 sky130_fd_sc_hd__dfxtp_1 _7194_ (.CLK(clknet_leaf_49_i_clk),
    .D(_0408_),
    .Q(\core_1.execute.alu_mul_div.mul_res[5] ));
 sky130_fd_sc_hd__dfxtp_1 _7195_ (.CLK(clknet_leaf_50_i_clk),
    .D(_0409_),
    .Q(\core_1.execute.alu_mul_div.mul_res[6] ));
 sky130_fd_sc_hd__dfxtp_1 _7196_ (.CLK(clknet_leaf_50_i_clk),
    .D(_0410_),
    .Q(\core_1.execute.alu_mul_div.mul_res[7] ));
 sky130_fd_sc_hd__dfxtp_1 _7197_ (.CLK(clknet_leaf_50_i_clk),
    .D(_0411_),
    .Q(\core_1.execute.alu_mul_div.mul_res[8] ));
 sky130_fd_sc_hd__dfxtp_1 _7198_ (.CLK(clknet_leaf_50_i_clk),
    .D(_0412_),
    .Q(\core_1.execute.alu_mul_div.mul_res[9] ));
 sky130_fd_sc_hd__dfxtp_1 _7199_ (.CLK(clknet_leaf_50_i_clk),
    .D(_0413_),
    .Q(\core_1.execute.alu_mul_div.mul_res[10] ));
 sky130_fd_sc_hd__dfxtp_1 _7200_ (.CLK(clknet_leaf_50_i_clk),
    .D(_0414_),
    .Q(\core_1.execute.alu_mul_div.mul_res[11] ));
 sky130_fd_sc_hd__dfxtp_1 _7201_ (.CLK(clknet_leaf_1_i_clk),
    .D(_0415_),
    .Q(\core_1.execute.alu_mul_div.mul_res[12] ));
 sky130_fd_sc_hd__dfxtp_1 _7202_ (.CLK(clknet_leaf_1_i_clk),
    .D(_0416_),
    .Q(\core_1.execute.alu_mul_div.mul_res[13] ));
 sky130_fd_sc_hd__dfxtp_1 _7203_ (.CLK(clknet_leaf_2_i_clk),
    .D(_0417_),
    .Q(\core_1.execute.alu_mul_div.mul_res[14] ));
 sky130_fd_sc_hd__dfxtp_1 _7204_ (.CLK(clknet_leaf_1_i_clk),
    .D(_0418_),
    .Q(\core_1.execute.alu_mul_div.mul_res[15] ));
 sky130_fd_sc_hd__dfxtp_1 _7205_ (.CLK(clknet_leaf_31_i_clk),
    .D(_0419_),
    .Q(\core_1.execute.next_ready_delayed ));
 sky130_fd_sc_hd__dfxtp_1 _7206_ (.CLK(clknet_leaf_2_i_clk),
    .D(_0420_),
    .Q(\core_1.execute.alu_mul_div.div_res[0] ));
 sky130_fd_sc_hd__dfxtp_1 _7207_ (.CLK(clknet_leaf_2_i_clk),
    .D(_0421_),
    .Q(\core_1.execute.alu_mul_div.div_res[1] ));
 sky130_fd_sc_hd__dfxtp_1 _7208_ (.CLK(clknet_leaf_2_i_clk),
    .D(_0422_),
    .Q(\core_1.execute.alu_mul_div.div_res[2] ));
 sky130_fd_sc_hd__dfxtp_1 _7209_ (.CLK(clknet_leaf_2_i_clk),
    .D(_0423_),
    .Q(\core_1.execute.alu_mul_div.div_res[3] ));
 sky130_fd_sc_hd__dfxtp_1 _7210_ (.CLK(clknet_leaf_2_i_clk),
    .D(_0424_),
    .Q(\core_1.execute.alu_mul_div.div_res[4] ));
 sky130_fd_sc_hd__dfxtp_1 _7211_ (.CLK(clknet_leaf_8_i_clk),
    .D(_0425_),
    .Q(\core_1.execute.alu_mul_div.div_res[5] ));
 sky130_fd_sc_hd__dfxtp_1 _7212_ (.CLK(clknet_leaf_7_i_clk),
    .D(_0426_),
    .Q(\core_1.execute.alu_mul_div.div_res[6] ));
 sky130_fd_sc_hd__dfxtp_1 _7213_ (.CLK(clknet_leaf_2_i_clk),
    .D(_0427_),
    .Q(\core_1.execute.alu_mul_div.div_res[7] ));
 sky130_fd_sc_hd__dfxtp_1 _7214_ (.CLK(clknet_leaf_2_i_clk),
    .D(_0428_),
    .Q(\core_1.execute.alu_mul_div.div_res[8] ));
 sky130_fd_sc_hd__dfxtp_1 _7215_ (.CLK(clknet_leaf_8_i_clk),
    .D(_0429_),
    .Q(\core_1.execute.alu_mul_div.div_res[9] ));
 sky130_fd_sc_hd__dfxtp_1 _7216_ (.CLK(clknet_leaf_8_i_clk),
    .D(_0430_),
    .Q(\core_1.execute.alu_mul_div.div_res[10] ));
 sky130_fd_sc_hd__dfxtp_1 _7217_ (.CLK(clknet_leaf_2_i_clk),
    .D(_0431_),
    .Q(\core_1.execute.alu_mul_div.div_res[11] ));
 sky130_fd_sc_hd__dfxtp_1 _7218_ (.CLK(clknet_leaf_2_i_clk),
    .D(_0432_),
    .Q(\core_1.execute.alu_mul_div.div_res[12] ));
 sky130_fd_sc_hd__dfxtp_1 _7219_ (.CLK(clknet_leaf_2_i_clk),
    .D(_0433_),
    .Q(\core_1.execute.alu_mul_div.div_res[13] ));
 sky130_fd_sc_hd__dfxtp_1 _7220_ (.CLK(clknet_leaf_8_i_clk),
    .D(_0434_),
    .Q(\core_1.execute.alu_mul_div.div_res[14] ));
 sky130_fd_sc_hd__dfxtp_1 _7221_ (.CLK(clknet_leaf_2_i_clk),
    .D(_0435_),
    .Q(\core_1.execute.alu_mul_div.div_res[15] ));
 sky130_fd_sc_hd__dfxtp_1 _7222_ (.CLK(clknet_leaf_35_i_clk),
    .D(_0436_),
    .Q(net72));
 sky130_fd_sc_hd__dfxtp_4 _7223_ (.CLK(clknet_leaf_34_i_clk),
    .D(_0437_),
    .Q(net80));
 sky130_fd_sc_hd__dfxtp_4 _7224_ (.CLK(clknet_leaf_34_i_clk),
    .D(_0438_),
    .Q(net81));
 sky130_fd_sc_hd__dfxtp_4 _7225_ (.CLK(clknet_leaf_35_i_clk),
    .D(_0439_),
    .Q(net82));
 sky130_fd_sc_hd__dfxtp_4 _7226_ (.CLK(clknet_leaf_35_i_clk),
    .D(_0440_),
    .Q(net83));
 sky130_fd_sc_hd__dfxtp_4 _7227_ (.CLK(clknet_leaf_35_i_clk),
    .D(_0441_),
    .Q(net84));
 sky130_fd_sc_hd__dfxtp_4 _7228_ (.CLK(clknet_leaf_35_i_clk),
    .D(_0442_),
    .Q(net85));
 sky130_fd_sc_hd__dfxtp_4 _7229_ (.CLK(clknet_leaf_35_i_clk),
    .D(_0443_),
    .Q(net86));
 sky130_fd_sc_hd__dfxtp_4 _7230_ (.CLK(clknet_leaf_27_i_clk),
    .D(_0444_),
    .Q(net87));
 sky130_fd_sc_hd__dfxtp_2 _7231_ (.CLK(clknet_leaf_28_i_clk),
    .D(_0445_),
    .Q(net73));
 sky130_fd_sc_hd__dfxtp_2 _7232_ (.CLK(clknet_leaf_28_i_clk),
    .D(_0446_),
    .Q(net74));
 sky130_fd_sc_hd__dfxtp_4 _7233_ (.CLK(clknet_leaf_28_i_clk),
    .D(_0447_),
    .Q(net75));
 sky130_fd_sc_hd__dfxtp_4 _7234_ (.CLK(clknet_leaf_27_i_clk),
    .D(_0448_),
    .Q(net76));
 sky130_fd_sc_hd__dfxtp_4 _7235_ (.CLK(clknet_leaf_34_i_clk),
    .D(_0449_),
    .Q(net77));
 sky130_fd_sc_hd__dfxtp_4 _7236_ (.CLK(clknet_leaf_28_i_clk),
    .D(_0450_),
    .Q(net78));
 sky130_fd_sc_hd__dfxtp_2 _7237_ (.CLK(clknet_leaf_46_i_clk),
    .D(_0451_),
    .Q(\core_1.execute.alu_flag_reg.o_d[0] ));
 sky130_fd_sc_hd__dfxtp_2 _7238_ (.CLK(clknet_leaf_47_i_clk),
    .D(_0452_),
    .Q(\core_1.execute.alu_flag_reg.o_d[1] ));
 sky130_fd_sc_hd__dfxtp_1 _7239_ (.CLK(clknet_leaf_45_i_clk),
    .D(_0453_),
    .Q(\core_1.execute.alu_flag_reg.o_d[2] ));
 sky130_fd_sc_hd__dfxtp_1 _7240_ (.CLK(clknet_leaf_46_i_clk),
    .D(_0454_),
    .Q(\core_1.execute.alu_flag_reg.o_d[3] ));
 sky130_fd_sc_hd__dfxtp_1 _7241_ (.CLK(clknet_leaf_46_i_clk),
    .D(_0455_),
    .Q(\core_1.execute.alu_flag_reg.o_d[4] ));
 sky130_fd_sc_hd__dfxtp_1 _7242_ (.CLK(clknet_leaf_33_i_clk),
    .D(_0456_),
    .Q(\core_1.execute.sreg_irq_pc.o_d[0] ));
 sky130_fd_sc_hd__dfxtp_1 _7243_ (.CLK(clknet_leaf_46_i_clk),
    .D(_0457_),
    .Q(\core_1.execute.sreg_irq_pc.o_d[1] ));
 sky130_fd_sc_hd__dfxtp_2 _7244_ (.CLK(clknet_leaf_33_i_clk),
    .D(_0458_),
    .Q(\core_1.execute.sreg_irq_pc.o_d[2] ));
 sky130_fd_sc_hd__dfxtp_1 _7245_ (.CLK(clknet_leaf_33_i_clk),
    .D(_0459_),
    .Q(\core_1.execute.sreg_irq_pc.o_d[3] ));
 sky130_fd_sc_hd__dfxtp_1 _7246_ (.CLK(clknet_leaf_33_i_clk),
    .D(_0460_),
    .Q(\core_1.execute.sreg_irq_pc.o_d[4] ));
 sky130_fd_sc_hd__dfxtp_2 _7247_ (.CLK(clknet_leaf_35_i_clk),
    .D(_0461_),
    .Q(\core_1.execute.sreg_irq_pc.o_d[5] ));
 sky130_fd_sc_hd__dfxtp_1 _7248_ (.CLK(clknet_leaf_32_i_clk),
    .D(_0462_),
    .Q(\core_1.execute.sreg_irq_pc.o_d[6] ));
 sky130_fd_sc_hd__dfxtp_1 _7249_ (.CLK(clknet_leaf_32_i_clk),
    .D(_0463_),
    .Q(\core_1.execute.sreg_irq_pc.o_d[7] ));
 sky130_fd_sc_hd__dfxtp_1 _7250_ (.CLK(clknet_leaf_30_i_clk),
    .D(_0464_),
    .Q(\core_1.execute.sreg_irq_pc.o_d[8] ));
 sky130_fd_sc_hd__dfxtp_1 _7251_ (.CLK(clknet_leaf_30_i_clk),
    .D(_0465_),
    .Q(\core_1.execute.sreg_irq_pc.o_d[9] ));
 sky130_fd_sc_hd__dfxtp_1 _7252_ (.CLK(clknet_leaf_30_i_clk),
    .D(_0466_),
    .Q(\core_1.execute.sreg_irq_pc.o_d[10] ));
 sky130_fd_sc_hd__dfxtp_1 _7253_ (.CLK(clknet_leaf_29_i_clk),
    .D(_0467_),
    .Q(\core_1.execute.sreg_irq_pc.o_d[11] ));
 sky130_fd_sc_hd__dfxtp_1 _7254_ (.CLK(clknet_leaf_29_i_clk),
    .D(_0468_),
    .Q(\core_1.execute.sreg_irq_pc.o_d[12] ));
 sky130_fd_sc_hd__dfxtp_1 _7255_ (.CLK(clknet_leaf_16_i_clk),
    .D(_0469_),
    .Q(\core_1.execute.sreg_irq_pc.o_d[13] ));
 sky130_fd_sc_hd__dfxtp_1 _7256_ (.CLK(clknet_leaf_29_i_clk),
    .D(_0470_),
    .Q(\core_1.execute.sreg_irq_pc.o_d[14] ));
 sky130_fd_sc_hd__dfxtp_1 _7257_ (.CLK(clknet_leaf_29_i_clk),
    .D(_0471_),
    .Q(\core_1.execute.sreg_irq_pc.o_d[15] ));
 sky130_fd_sc_hd__dfxtp_1 _7258_ (.CLK(clknet_leaf_42_i_clk),
    .D(_0472_),
    .Q(\core_1.execute.sreg_jtr_buff.o_d[0] ));
 sky130_fd_sc_hd__dfxtp_1 _7259_ (.CLK(clknet_leaf_43_i_clk),
    .D(_0473_),
    .Q(\core_1.execute.sreg_jtr_buff.o_d[1] ));
 sky130_fd_sc_hd__dfxtp_1 _7260_ (.CLK(clknet_leaf_43_i_clk),
    .D(_0474_),
    .Q(\core_1.execute.sreg_jtr_buff.o_d[2] ));
 sky130_fd_sc_hd__dfxtp_2 _7261_ (.CLK(clknet_leaf_42_i_clk),
    .D(_0475_),
    .Q(net106));
 sky130_fd_sc_hd__dfxtp_1 _7262_ (.CLK(clknet_leaf_43_i_clk),
    .D(_0476_),
    .Q(\core_1.execute.trap_flag ));
 sky130_fd_sc_hd__dfxtp_2 _7263_ (.CLK(clknet_leaf_41_i_clk),
    .D(_0477_),
    .Q(net105));
 sky130_fd_sc_hd__dfxtp_1 _7264_ (.CLK(clknet_leaf_39_i_clk),
    .D(_0478_),
    .Q(\core_1.execute.sreg_scratch.o_d[0] ));
 sky130_fd_sc_hd__dfxtp_1 _7265_ (.CLK(clknet_leaf_39_i_clk),
    .D(_0479_),
    .Q(\core_1.execute.sreg_scratch.o_d[1] ));
 sky130_fd_sc_hd__dfxtp_1 _7266_ (.CLK(clknet_leaf_39_i_clk),
    .D(_0480_),
    .Q(\core_1.execute.sreg_scratch.o_d[2] ));
 sky130_fd_sc_hd__dfxtp_1 _7267_ (.CLK(clknet_leaf_39_i_clk),
    .D(_0481_),
    .Q(\core_1.execute.sreg_scratch.o_d[3] ));
 sky130_fd_sc_hd__dfxtp_1 _7268_ (.CLK(clknet_leaf_37_i_clk),
    .D(_0482_),
    .Q(\core_1.execute.sreg_scratch.o_d[4] ));
 sky130_fd_sc_hd__dfxtp_1 _7269_ (.CLK(clknet_leaf_39_i_clk),
    .D(_0483_),
    .Q(\core_1.execute.sreg_scratch.o_d[5] ));
 sky130_fd_sc_hd__dfxtp_1 _7270_ (.CLK(clknet_leaf_36_i_clk),
    .D(_0484_),
    .Q(\core_1.execute.sreg_scratch.o_d[6] ));
 sky130_fd_sc_hd__dfxtp_1 _7271_ (.CLK(clknet_leaf_36_i_clk),
    .D(_0485_),
    .Q(\core_1.execute.sreg_scratch.o_d[7] ));
 sky130_fd_sc_hd__dfxtp_1 _7272_ (.CLK(clknet_leaf_27_i_clk),
    .D(_0486_),
    .Q(\core_1.execute.sreg_scratch.o_d[8] ));
 sky130_fd_sc_hd__dfxtp_1 _7273_ (.CLK(clknet_leaf_27_i_clk),
    .D(_0487_),
    .Q(\core_1.execute.sreg_scratch.o_d[9] ));
 sky130_fd_sc_hd__dfxtp_1 _7274_ (.CLK(clknet_leaf_25_i_clk),
    .D(_0488_),
    .Q(\core_1.execute.sreg_scratch.o_d[10] ));
 sky130_fd_sc_hd__dfxtp_1 _7275_ (.CLK(clknet_leaf_25_i_clk),
    .D(_0489_),
    .Q(\core_1.execute.sreg_scratch.o_d[11] ));
 sky130_fd_sc_hd__dfxtp_1 _7276_ (.CLK(clknet_leaf_25_i_clk),
    .D(_0490_),
    .Q(\core_1.execute.sreg_scratch.o_d[12] ));
 sky130_fd_sc_hd__dfxtp_1 _7277_ (.CLK(clknet_leaf_25_i_clk),
    .D(_0491_),
    .Q(\core_1.execute.sreg_scratch.o_d[13] ));
 sky130_fd_sc_hd__dfxtp_1 _7278_ (.CLK(clknet_leaf_25_i_clk),
    .D(_0492_),
    .Q(\core_1.execute.sreg_scratch.o_d[14] ));
 sky130_fd_sc_hd__dfxtp_1 _7279_ (.CLK(clknet_leaf_25_i_clk),
    .D(_0493_),
    .Q(\core_1.execute.sreg_scratch.o_d[15] ));
 sky130_fd_sc_hd__dfxtp_1 _7280_ (.CLK(clknet_leaf_41_i_clk),
    .D(_0494_),
    .Q(\core_1.execute.sreg_irq_flags.o_d[0] ));
 sky130_fd_sc_hd__dfxtp_1 _7281_ (.CLK(clknet_leaf_42_i_clk),
    .D(_0495_),
    .Q(\core_1.execute.sreg_irq_flags.o_d[1] ));
 sky130_fd_sc_hd__dfxtp_1 _7282_ (.CLK(clknet_leaf_38_i_clk),
    .D(_0496_),
    .Q(\core_1.execute.sreg_irq_flags.o_d[2] ));
 sky130_fd_sc_hd__dfxtp_1 _7283_ (.CLK(clknet_leaf_38_i_clk),
    .D(_0497_),
    .Q(\core_1.execute.sreg_irq_flags.o_d[3] ));
 sky130_fd_sc_hd__dfxtp_1 _7284_ (.CLK(clknet_leaf_41_i_clk),
    .D(_0498_),
    .Q(\core_1.execute.sreg_irq_flags.o_d[4] ));
 sky130_fd_sc_hd__dfxtp_2 _7285_ (.CLK(clknet_leaf_40_i_clk),
    .D(_0499_),
    .Q(\core_1.execute.pc_high_out[0] ));
 sky130_fd_sc_hd__dfxtp_2 _7286_ (.CLK(clknet_leaf_40_i_clk),
    .D(_0500_),
    .Q(\core_1.execute.pc_high_out[1] ));
 sky130_fd_sc_hd__dfxtp_2 _7287_ (.CLK(clknet_leaf_40_i_clk),
    .D(_0501_),
    .Q(\core_1.execute.pc_high_out[2] ));
 sky130_fd_sc_hd__dfxtp_2 _7288_ (.CLK(clknet_leaf_40_i_clk),
    .D(_0502_),
    .Q(\core_1.execute.pc_high_out[3] ));
 sky130_fd_sc_hd__dfxtp_2 _7289_ (.CLK(clknet_leaf_39_i_clk),
    .D(_0503_),
    .Q(\core_1.execute.pc_high_out[4] ));
 sky130_fd_sc_hd__dfxtp_2 _7290_ (.CLK(clknet_leaf_39_i_clk),
    .D(_0504_),
    .Q(\core_1.execute.pc_high_out[5] ));
 sky130_fd_sc_hd__dfxtp_2 _7291_ (.CLK(clknet_leaf_39_i_clk),
    .D(_0505_),
    .Q(\core_1.execute.pc_high_out[6] ));
 sky130_fd_sc_hd__dfxtp_2 _7292_ (.CLK(clknet_leaf_41_i_clk),
    .D(_0506_),
    .Q(\core_1.execute.pc_high_out[7] ));
 sky130_fd_sc_hd__dfxtp_1 _7293_ (.CLK(clknet_leaf_41_i_clk),
    .D(_0507_),
    .Q(\core_1.execute.pc_high_buff_out[0] ));
 sky130_fd_sc_hd__dfxtp_1 _7294_ (.CLK(clknet_leaf_40_i_clk),
    .D(_0508_),
    .Q(\core_1.execute.pc_high_buff_out[1] ));
 sky130_fd_sc_hd__dfxtp_1 _7295_ (.CLK(clknet_leaf_41_i_clk),
    .D(_0509_),
    .Q(\core_1.execute.pc_high_buff_out[2] ));
 sky130_fd_sc_hd__dfxtp_1 _7296_ (.CLK(clknet_leaf_40_i_clk),
    .D(_0510_),
    .Q(\core_1.execute.pc_high_buff_out[3] ));
 sky130_fd_sc_hd__dfxtp_1 _7297_ (.CLK(clknet_leaf_41_i_clk),
    .D(_0511_),
    .Q(\core_1.execute.pc_high_buff_out[4] ));
 sky130_fd_sc_hd__dfxtp_1 _7298_ (.CLK(clknet_leaf_40_i_clk),
    .D(_0512_),
    .Q(\core_1.execute.pc_high_buff_out[5] ));
 sky130_fd_sc_hd__dfxtp_2 _7299_ (.CLK(clknet_leaf_41_i_clk),
    .D(_0513_),
    .Q(\core_1.execute.pc_high_buff_out[6] ));
 sky130_fd_sc_hd__dfxtp_2 _7300_ (.CLK(clknet_leaf_42_i_clk),
    .D(_0514_),
    .Q(\core_1.execute.pc_high_buff_out[7] ));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_0_i_clk (.A(clknet_2_0_0_i_clk),
    .X(clknet_leaf_0_i_clk));
 sky130_fd_sc_hd__decap_3 PHY_0 ();
 sky130_fd_sc_hd__decap_3 PHY_1 ();
 sky130_fd_sc_hd__decap_3 PHY_2 ();
 sky130_fd_sc_hd__decap_3 PHY_3 ();
 sky130_fd_sc_hd__decap_3 PHY_4 ();
 sky130_fd_sc_hd__decap_3 PHY_5 ();
 sky130_fd_sc_hd__decap_3 PHY_6 ();
 sky130_fd_sc_hd__decap_3 PHY_7 ();
 sky130_fd_sc_hd__decap_3 PHY_8 ();
 sky130_fd_sc_hd__decap_3 PHY_9 ();
 sky130_fd_sc_hd__decap_3 PHY_10 ();
 sky130_fd_sc_hd__decap_3 PHY_11 ();
 sky130_fd_sc_hd__decap_3 PHY_12 ();
 sky130_fd_sc_hd__decap_3 PHY_13 ();
 sky130_fd_sc_hd__decap_3 PHY_14 ();
 sky130_fd_sc_hd__decap_3 PHY_15 ();
 sky130_fd_sc_hd__decap_3 PHY_16 ();
 sky130_fd_sc_hd__decap_3 PHY_17 ();
 sky130_fd_sc_hd__decap_3 PHY_18 ();
 sky130_fd_sc_hd__decap_3 PHY_19 ();
 sky130_fd_sc_hd__decap_3 PHY_20 ();
 sky130_fd_sc_hd__decap_3 PHY_21 ();
 sky130_fd_sc_hd__decap_3 PHY_22 ();
 sky130_fd_sc_hd__decap_3 PHY_23 ();
 sky130_fd_sc_hd__decap_3 PHY_24 ();
 sky130_fd_sc_hd__decap_3 PHY_25 ();
 sky130_fd_sc_hd__decap_3 PHY_26 ();
 sky130_fd_sc_hd__decap_3 PHY_27 ();
 sky130_fd_sc_hd__decap_3 PHY_28 ();
 sky130_fd_sc_hd__decap_3 PHY_29 ();
 sky130_fd_sc_hd__decap_3 PHY_30 ();
 sky130_fd_sc_hd__decap_3 PHY_31 ();
 sky130_fd_sc_hd__decap_3 PHY_32 ();
 sky130_fd_sc_hd__decap_3 PHY_33 ();
 sky130_fd_sc_hd__decap_3 PHY_34 ();
 sky130_fd_sc_hd__decap_3 PHY_35 ();
 sky130_fd_sc_hd__decap_3 PHY_36 ();
 sky130_fd_sc_hd__decap_3 PHY_37 ();
 sky130_fd_sc_hd__decap_3 PHY_38 ();
 sky130_fd_sc_hd__decap_3 PHY_39 ();
 sky130_fd_sc_hd__decap_3 PHY_40 ();
 sky130_fd_sc_hd__decap_3 PHY_41 ();
 sky130_fd_sc_hd__decap_3 PHY_42 ();
 sky130_fd_sc_hd__decap_3 PHY_43 ();
 sky130_fd_sc_hd__decap_3 PHY_44 ();
 sky130_fd_sc_hd__decap_3 PHY_45 ();
 sky130_fd_sc_hd__decap_3 PHY_46 ();
 sky130_fd_sc_hd__decap_3 PHY_47 ();
 sky130_fd_sc_hd__decap_3 PHY_48 ();
 sky130_fd_sc_hd__decap_3 PHY_49 ();
 sky130_fd_sc_hd__decap_3 PHY_50 ();
 sky130_fd_sc_hd__decap_3 PHY_51 ();
 sky130_fd_sc_hd__decap_3 PHY_52 ();
 sky130_fd_sc_hd__decap_3 PHY_53 ();
 sky130_fd_sc_hd__decap_3 PHY_54 ();
 sky130_fd_sc_hd__decap_3 PHY_55 ();
 sky130_fd_sc_hd__decap_3 PHY_56 ();
 sky130_fd_sc_hd__decap_3 PHY_57 ();
 sky130_fd_sc_hd__decap_3 PHY_58 ();
 sky130_fd_sc_hd__decap_3 PHY_59 ();
 sky130_fd_sc_hd__decap_3 PHY_60 ();
 sky130_fd_sc_hd__decap_3 PHY_61 ();
 sky130_fd_sc_hd__decap_3 PHY_62 ();
 sky130_fd_sc_hd__decap_3 PHY_63 ();
 sky130_fd_sc_hd__decap_3 PHY_64 ();
 sky130_fd_sc_hd__decap_3 PHY_65 ();
 sky130_fd_sc_hd__decap_3 PHY_66 ();
 sky130_fd_sc_hd__decap_3 PHY_67 ();
 sky130_fd_sc_hd__decap_3 PHY_68 ();
 sky130_fd_sc_hd__decap_3 PHY_69 ();
 sky130_fd_sc_hd__decap_3 PHY_70 ();
 sky130_fd_sc_hd__decap_3 PHY_71 ();
 sky130_fd_sc_hd__decap_3 PHY_72 ();
 sky130_fd_sc_hd__decap_3 PHY_73 ();
 sky130_fd_sc_hd__decap_3 PHY_74 ();
 sky130_fd_sc_hd__decap_3 PHY_75 ();
 sky130_fd_sc_hd__decap_3 PHY_76 ();
 sky130_fd_sc_hd__decap_3 PHY_77 ();
 sky130_fd_sc_hd__decap_3 PHY_78 ();
 sky130_fd_sc_hd__decap_3 PHY_79 ();
 sky130_fd_sc_hd__decap_3 PHY_80 ();
 sky130_fd_sc_hd__decap_3 PHY_81 ();
 sky130_fd_sc_hd__decap_3 PHY_82 ();
 sky130_fd_sc_hd__decap_3 PHY_83 ();
 sky130_fd_sc_hd__decap_3 PHY_84 ();
 sky130_fd_sc_hd__decap_3 PHY_85 ();
 sky130_fd_sc_hd__decap_3 PHY_86 ();
 sky130_fd_sc_hd__decap_3 PHY_87 ();
 sky130_fd_sc_hd__decap_3 PHY_88 ();
 sky130_fd_sc_hd__decap_3 PHY_89 ();
 sky130_fd_sc_hd__decap_3 PHY_90 ();
 sky130_fd_sc_hd__decap_3 PHY_91 ();
 sky130_fd_sc_hd__decap_3 PHY_92 ();
 sky130_fd_sc_hd__decap_3 PHY_93 ();
 sky130_fd_sc_hd__decap_3 PHY_94 ();
 sky130_fd_sc_hd__decap_3 PHY_95 ();
 sky130_fd_sc_hd__decap_3 PHY_96 ();
 sky130_fd_sc_hd__decap_3 PHY_97 ();
 sky130_fd_sc_hd__decap_3 PHY_98 ();
 sky130_fd_sc_hd__decap_3 PHY_99 ();
 sky130_fd_sc_hd__decap_3 PHY_100 ();
 sky130_fd_sc_hd__decap_3 PHY_101 ();
 sky130_fd_sc_hd__decap_3 PHY_102 ();
 sky130_fd_sc_hd__decap_3 PHY_103 ();
 sky130_fd_sc_hd__decap_3 PHY_104 ();
 sky130_fd_sc_hd__decap_3 PHY_105 ();
 sky130_fd_sc_hd__decap_3 PHY_106 ();
 sky130_fd_sc_hd__decap_3 PHY_107 ();
 sky130_fd_sc_hd__decap_3 PHY_108 ();
 sky130_fd_sc_hd__decap_3 PHY_109 ();
 sky130_fd_sc_hd__decap_3 PHY_110 ();
 sky130_fd_sc_hd__decap_3 PHY_111 ();
 sky130_fd_sc_hd__decap_3 PHY_112 ();
 sky130_fd_sc_hd__decap_3 PHY_113 ();
 sky130_fd_sc_hd__decap_3 PHY_114 ();
 sky130_fd_sc_hd__decap_3 PHY_115 ();
 sky130_fd_sc_hd__decap_3 PHY_116 ();
 sky130_fd_sc_hd__decap_3 PHY_117 ();
 sky130_fd_sc_hd__decap_3 PHY_118 ();
 sky130_fd_sc_hd__decap_3 PHY_119 ();
 sky130_fd_sc_hd__decap_3 PHY_120 ();
 sky130_fd_sc_hd__decap_3 PHY_121 ();
 sky130_fd_sc_hd__decap_3 PHY_122 ();
 sky130_fd_sc_hd__decap_3 PHY_123 ();
 sky130_fd_sc_hd__decap_3 PHY_124 ();
 sky130_fd_sc_hd__decap_3 PHY_125 ();
 sky130_fd_sc_hd__decap_3 PHY_126 ();
 sky130_fd_sc_hd__decap_3 PHY_127 ();
 sky130_fd_sc_hd__decap_3 PHY_128 ();
 sky130_fd_sc_hd__decap_3 PHY_129 ();
 sky130_fd_sc_hd__decap_3 PHY_130 ();
 sky130_fd_sc_hd__decap_3 PHY_131 ();
 sky130_fd_sc_hd__decap_3 PHY_132 ();
 sky130_fd_sc_hd__decap_3 PHY_133 ();
 sky130_fd_sc_hd__decap_3 PHY_134 ();
 sky130_fd_sc_hd__decap_3 PHY_135 ();
 sky130_fd_sc_hd__decap_3 PHY_136 ();
 sky130_fd_sc_hd__decap_3 PHY_137 ();
 sky130_fd_sc_hd__decap_3 PHY_138 ();
 sky130_fd_sc_hd__decap_3 PHY_139 ();
 sky130_fd_sc_hd__decap_3 PHY_140 ();
 sky130_fd_sc_hd__decap_3 PHY_141 ();
 sky130_fd_sc_hd__decap_3 PHY_142 ();
 sky130_fd_sc_hd__decap_3 PHY_143 ();
 sky130_fd_sc_hd__decap_3 PHY_144 ();
 sky130_fd_sc_hd__decap_3 PHY_145 ();
 sky130_fd_sc_hd__decap_3 PHY_146 ();
 sky130_fd_sc_hd__decap_3 PHY_147 ();
 sky130_fd_sc_hd__decap_3 PHY_148 ();
 sky130_fd_sc_hd__decap_3 PHY_149 ();
 sky130_fd_sc_hd__decap_3 PHY_150 ();
 sky130_fd_sc_hd__decap_3 PHY_151 ();
 sky130_fd_sc_hd__decap_3 PHY_152 ();
 sky130_fd_sc_hd__decap_3 PHY_153 ();
 sky130_fd_sc_hd__decap_3 PHY_154 ();
 sky130_fd_sc_hd__decap_3 PHY_155 ();
 sky130_fd_sc_hd__decap_3 PHY_156 ();
 sky130_fd_sc_hd__decap_3 PHY_157 ();
 sky130_fd_sc_hd__decap_3 PHY_158 ();
 sky130_fd_sc_hd__decap_3 PHY_159 ();
 sky130_fd_sc_hd__decap_3 PHY_160 ();
 sky130_fd_sc_hd__decap_3 PHY_161 ();
 sky130_fd_sc_hd__decap_3 PHY_162 ();
 sky130_fd_sc_hd__decap_3 PHY_163 ();
 sky130_fd_sc_hd__decap_3 PHY_164 ();
 sky130_fd_sc_hd__decap_3 PHY_165 ();
 sky130_fd_sc_hd__decap_3 PHY_166 ();
 sky130_fd_sc_hd__decap_3 PHY_167 ();
 sky130_fd_sc_hd__decap_3 PHY_168 ();
 sky130_fd_sc_hd__decap_3 PHY_169 ();
 sky130_fd_sc_hd__decap_3 PHY_170 ();
 sky130_fd_sc_hd__decap_3 PHY_171 ();
 sky130_fd_sc_hd__decap_3 PHY_172 ();
 sky130_fd_sc_hd__decap_3 PHY_173 ();
 sky130_fd_sc_hd__decap_3 PHY_174 ();
 sky130_fd_sc_hd__decap_3 PHY_175 ();
 sky130_fd_sc_hd__decap_3 PHY_176 ();
 sky130_fd_sc_hd__decap_3 PHY_177 ();
 sky130_fd_sc_hd__decap_3 PHY_178 ();
 sky130_fd_sc_hd__decap_3 PHY_179 ();
 sky130_fd_sc_hd__decap_3 PHY_180 ();
 sky130_fd_sc_hd__decap_3 PHY_181 ();
 sky130_fd_sc_hd__decap_3 PHY_182 ();
 sky130_fd_sc_hd__decap_3 PHY_183 ();
 sky130_fd_sc_hd__decap_3 PHY_184 ();
 sky130_fd_sc_hd__decap_3 PHY_185 ();
 sky130_fd_sc_hd__decap_3 PHY_186 ();
 sky130_fd_sc_hd__decap_3 PHY_187 ();
 sky130_fd_sc_hd__decap_3 PHY_188 ();
 sky130_fd_sc_hd__decap_3 PHY_189 ();
 sky130_fd_sc_hd__decap_3 PHY_190 ();
 sky130_fd_sc_hd__decap_3 PHY_191 ();
 sky130_fd_sc_hd__decap_3 PHY_192 ();
 sky130_fd_sc_hd__decap_3 PHY_193 ();
 sky130_fd_sc_hd__decap_3 PHY_194 ();
 sky130_fd_sc_hd__decap_3 PHY_195 ();
 sky130_fd_sc_hd__decap_3 PHY_196 ();
 sky130_fd_sc_hd__decap_3 PHY_197 ();
 sky130_fd_sc_hd__decap_3 PHY_198 ();
 sky130_fd_sc_hd__decap_3 PHY_199 ();
 sky130_fd_sc_hd__decap_3 PHY_200 ();
 sky130_fd_sc_hd__decap_3 PHY_201 ();
 sky130_fd_sc_hd__decap_3 PHY_202 ();
 sky130_fd_sc_hd__decap_3 PHY_203 ();
 sky130_fd_sc_hd__decap_3 PHY_204 ();
 sky130_fd_sc_hd__decap_3 PHY_205 ();
 sky130_fd_sc_hd__decap_3 PHY_206 ();
 sky130_fd_sc_hd__decap_3 PHY_207 ();
 sky130_fd_sc_hd__decap_3 PHY_208 ();
 sky130_fd_sc_hd__decap_3 PHY_209 ();
 sky130_fd_sc_hd__decap_3 PHY_210 ();
 sky130_fd_sc_hd__decap_3 PHY_211 ();
 sky130_fd_sc_hd__decap_3 PHY_212 ();
 sky130_fd_sc_hd__decap_3 PHY_213 ();
 sky130_fd_sc_hd__decap_3 PHY_214 ();
 sky130_fd_sc_hd__decap_3 PHY_215 ();
 sky130_fd_sc_hd__decap_3 PHY_216 ();
 sky130_fd_sc_hd__decap_3 PHY_217 ();
 sky130_fd_sc_hd__decap_3 PHY_218 ();
 sky130_fd_sc_hd__decap_3 PHY_219 ();
 sky130_fd_sc_hd__decap_3 PHY_220 ();
 sky130_fd_sc_hd__decap_3 PHY_221 ();
 sky130_fd_sc_hd__decap_3 PHY_222 ();
 sky130_fd_sc_hd__decap_3 PHY_223 ();
 sky130_fd_sc_hd__decap_3 PHY_224 ();
 sky130_fd_sc_hd__decap_3 PHY_225 ();
 sky130_fd_sc_hd__decap_3 PHY_226 ();
 sky130_fd_sc_hd__decap_3 PHY_227 ();
 sky130_fd_sc_hd__decap_3 PHY_228 ();
 sky130_fd_sc_hd__decap_3 PHY_229 ();
 sky130_fd_sc_hd__decap_3 PHY_230 ();
 sky130_fd_sc_hd__decap_3 PHY_231 ();
 sky130_fd_sc_hd__decap_3 PHY_232 ();
 sky130_fd_sc_hd__decap_3 PHY_233 ();
 sky130_fd_sc_hd__decap_3 PHY_234 ();
 sky130_fd_sc_hd__decap_3 PHY_235 ();
 sky130_fd_sc_hd__decap_3 PHY_236 ();
 sky130_fd_sc_hd__decap_3 PHY_237 ();
 sky130_fd_sc_hd__decap_3 PHY_238 ();
 sky130_fd_sc_hd__decap_3 PHY_239 ();
 sky130_fd_sc_hd__decap_3 PHY_240 ();
 sky130_fd_sc_hd__decap_3 PHY_241 ();
 sky130_fd_sc_hd__decap_3 PHY_242 ();
 sky130_fd_sc_hd__decap_3 PHY_243 ();
 sky130_fd_sc_hd__decap_3 PHY_244 ();
 sky130_fd_sc_hd__decap_3 PHY_245 ();
 sky130_fd_sc_hd__decap_3 PHY_246 ();
 sky130_fd_sc_hd__decap_3 PHY_247 ();
 sky130_fd_sc_hd__decap_3 PHY_248 ();
 sky130_fd_sc_hd__decap_3 PHY_249 ();
 sky130_fd_sc_hd__decap_3 PHY_250 ();
 sky130_fd_sc_hd__decap_3 PHY_251 ();
 sky130_fd_sc_hd__decap_3 PHY_252 ();
 sky130_fd_sc_hd__decap_3 PHY_253 ();
 sky130_fd_sc_hd__decap_3 PHY_254 ();
 sky130_fd_sc_hd__decap_3 PHY_255 ();
 sky130_fd_sc_hd__decap_3 PHY_256 ();
 sky130_fd_sc_hd__decap_3 PHY_257 ();
 sky130_fd_sc_hd__decap_3 PHY_258 ();
 sky130_fd_sc_hd__decap_3 PHY_259 ();
 sky130_fd_sc_hd__decap_3 PHY_260 ();
 sky130_fd_sc_hd__decap_3 PHY_261 ();
 sky130_fd_sc_hd__decap_3 PHY_262 ();
 sky130_fd_sc_hd__decap_3 PHY_263 ();
 sky130_fd_sc_hd__decap_3 PHY_264 ();
 sky130_fd_sc_hd__decap_3 PHY_265 ();
 sky130_fd_sc_hd__decap_3 PHY_266 ();
 sky130_fd_sc_hd__decap_3 PHY_267 ();
 sky130_fd_sc_hd__decap_3 PHY_268 ();
 sky130_fd_sc_hd__decap_3 PHY_269 ();
 sky130_fd_sc_hd__decap_3 PHY_270 ();
 sky130_fd_sc_hd__decap_3 PHY_271 ();
 sky130_fd_sc_hd__decap_3 PHY_272 ();
 sky130_fd_sc_hd__decap_3 PHY_273 ();
 sky130_fd_sc_hd__decap_3 PHY_274 ();
 sky130_fd_sc_hd__decap_3 PHY_275 ();
 sky130_fd_sc_hd__decap_3 PHY_276 ();
 sky130_fd_sc_hd__decap_3 PHY_277 ();
 sky130_fd_sc_hd__decap_3 PHY_278 ();
 sky130_fd_sc_hd__decap_3 PHY_279 ();
 sky130_fd_sc_hd__decap_3 PHY_280 ();
 sky130_fd_sc_hd__decap_3 PHY_281 ();
 sky130_fd_sc_hd__decap_3 PHY_282 ();
 sky130_fd_sc_hd__decap_3 PHY_283 ();
 sky130_fd_sc_hd__decap_3 PHY_284 ();
 sky130_fd_sc_hd__decap_3 PHY_285 ();
 sky130_fd_sc_hd__decap_3 PHY_286 ();
 sky130_fd_sc_hd__decap_3 PHY_287 ();
 sky130_fd_sc_hd__decap_3 PHY_288 ();
 sky130_fd_sc_hd__decap_3 PHY_289 ();
 sky130_fd_sc_hd__decap_3 PHY_290 ();
 sky130_fd_sc_hd__decap_3 PHY_291 ();
 sky130_fd_sc_hd__decap_3 PHY_292 ();
 sky130_fd_sc_hd__decap_3 PHY_293 ();
 sky130_fd_sc_hd__decap_3 PHY_294 ();
 sky130_fd_sc_hd__decap_3 PHY_295 ();
 sky130_fd_sc_hd__decap_3 PHY_296 ();
 sky130_fd_sc_hd__decap_3 PHY_297 ();
 sky130_fd_sc_hd__decap_3 PHY_298 ();
 sky130_fd_sc_hd__decap_3 PHY_299 ();
 sky130_fd_sc_hd__decap_3 PHY_300 ();
 sky130_fd_sc_hd__decap_3 PHY_301 ();
 sky130_fd_sc_hd__decap_3 PHY_302 ();
 sky130_fd_sc_hd__decap_3 PHY_303 ();
 sky130_fd_sc_hd__decap_3 PHY_304 ();
 sky130_fd_sc_hd__decap_3 PHY_305 ();
 sky130_fd_sc_hd__decap_3 PHY_306 ();
 sky130_fd_sc_hd__decap_3 PHY_307 ();
 sky130_fd_sc_hd__decap_3 PHY_308 ();
 sky130_fd_sc_hd__decap_3 PHY_309 ();
 sky130_fd_sc_hd__decap_3 PHY_310 ();
 sky130_fd_sc_hd__decap_3 PHY_311 ();
 sky130_fd_sc_hd__decap_3 PHY_312 ();
 sky130_fd_sc_hd__decap_3 PHY_313 ();
 sky130_fd_sc_hd__decap_3 PHY_314 ();
 sky130_fd_sc_hd__decap_3 PHY_315 ();
 sky130_fd_sc_hd__decap_3 PHY_316 ();
 sky130_fd_sc_hd__decap_3 PHY_317 ();
 sky130_fd_sc_hd__decap_3 PHY_318 ();
 sky130_fd_sc_hd__decap_3 PHY_319 ();
 sky130_fd_sc_hd__decap_3 PHY_320 ();
 sky130_fd_sc_hd__decap_3 PHY_321 ();
 sky130_fd_sc_hd__decap_3 PHY_322 ();
 sky130_fd_sc_hd__decap_3 PHY_323 ();
 sky130_fd_sc_hd__decap_3 PHY_324 ();
 sky130_fd_sc_hd__decap_3 PHY_325 ();
 sky130_fd_sc_hd__decap_3 PHY_326 ();
 sky130_fd_sc_hd__decap_3 PHY_327 ();
 sky130_fd_sc_hd__decap_3 PHY_328 ();
 sky130_fd_sc_hd__decap_3 PHY_329 ();
 sky130_fd_sc_hd__decap_3 PHY_330 ();
 sky130_fd_sc_hd__decap_3 PHY_331 ();
 sky130_fd_sc_hd__decap_3 PHY_332 ();
 sky130_fd_sc_hd__decap_3 PHY_333 ();
 sky130_fd_sc_hd__decap_3 PHY_334 ();
 sky130_fd_sc_hd__decap_3 PHY_335 ();
 sky130_fd_sc_hd__decap_3 PHY_336 ();
 sky130_fd_sc_hd__decap_3 PHY_337 ();
 sky130_fd_sc_hd__decap_3 PHY_338 ();
 sky130_fd_sc_hd__decap_3 PHY_339 ();
 sky130_fd_sc_hd__decap_3 PHY_340 ();
 sky130_fd_sc_hd__decap_3 PHY_341 ();
 sky130_fd_sc_hd__decap_3 PHY_342 ();
 sky130_fd_sc_hd__decap_3 PHY_343 ();
 sky130_fd_sc_hd__decap_3 PHY_344 ();
 sky130_fd_sc_hd__decap_3 PHY_345 ();
 sky130_fd_sc_hd__decap_3 PHY_346 ();
 sky130_fd_sc_hd__decap_3 PHY_347 ();
 sky130_fd_sc_hd__decap_3 PHY_348 ();
 sky130_fd_sc_hd__decap_3 PHY_349 ();
 sky130_fd_sc_hd__decap_3 PHY_350 ();
 sky130_fd_sc_hd__decap_3 PHY_351 ();
 sky130_fd_sc_hd__decap_3 PHY_352 ();
 sky130_fd_sc_hd__decap_3 PHY_353 ();
 sky130_fd_sc_hd__decap_3 PHY_354 ();
 sky130_fd_sc_hd__decap_3 PHY_355 ();
 sky130_fd_sc_hd__decap_3 PHY_356 ();
 sky130_fd_sc_hd__decap_3 PHY_357 ();
 sky130_fd_sc_hd__decap_3 PHY_358 ();
 sky130_fd_sc_hd__decap_3 PHY_359 ();
 sky130_fd_sc_hd__decap_3 PHY_360 ();
 sky130_fd_sc_hd__decap_3 PHY_361 ();
 sky130_fd_sc_hd__decap_3 PHY_362 ();
 sky130_fd_sc_hd__decap_3 PHY_363 ();
 sky130_fd_sc_hd__decap_3 PHY_364 ();
 sky130_fd_sc_hd__decap_3 PHY_365 ();
 sky130_fd_sc_hd__decap_3 PHY_366 ();
 sky130_fd_sc_hd__decap_3 PHY_367 ();
 sky130_fd_sc_hd__decap_3 PHY_368 ();
 sky130_fd_sc_hd__decap_3 PHY_369 ();
 sky130_fd_sc_hd__decap_3 PHY_370 ();
 sky130_fd_sc_hd__decap_3 PHY_371 ();
 sky130_fd_sc_hd__decap_3 PHY_372 ();
 sky130_fd_sc_hd__decap_3 PHY_373 ();
 sky130_fd_sc_hd__decap_3 PHY_374 ();
 sky130_fd_sc_hd__decap_3 PHY_375 ();
 sky130_fd_sc_hd__decap_3 PHY_376 ();
 sky130_fd_sc_hd__decap_3 PHY_377 ();
 sky130_fd_sc_hd__decap_3 PHY_378 ();
 sky130_fd_sc_hd__decap_3 PHY_379 ();
 sky130_fd_sc_hd__decap_3 PHY_380 ();
 sky130_fd_sc_hd__decap_3 PHY_381 ();
 sky130_fd_sc_hd__decap_3 PHY_382 ();
 sky130_fd_sc_hd__decap_3 PHY_383 ();
 sky130_fd_sc_hd__decap_3 PHY_384 ();
 sky130_fd_sc_hd__decap_3 PHY_385 ();
 sky130_fd_sc_hd__decap_3 PHY_386 ();
 sky130_fd_sc_hd__decap_3 PHY_387 ();
 sky130_fd_sc_hd__decap_3 PHY_388 ();
 sky130_fd_sc_hd__decap_3 PHY_389 ();
 sky130_fd_sc_hd__decap_3 PHY_390 ();
 sky130_fd_sc_hd__decap_3 PHY_391 ();
 sky130_fd_sc_hd__decap_3 PHY_392 ();
 sky130_fd_sc_hd__decap_3 PHY_393 ();
 sky130_fd_sc_hd__decap_3 PHY_394 ();
 sky130_fd_sc_hd__decap_3 PHY_395 ();
 sky130_fd_sc_hd__decap_3 PHY_396 ();
 sky130_fd_sc_hd__decap_3 PHY_397 ();
 sky130_fd_sc_hd__decap_3 PHY_398 ();
 sky130_fd_sc_hd__decap_3 PHY_399 ();
 sky130_fd_sc_hd__decap_3 PHY_400 ();
 sky130_fd_sc_hd__decap_3 PHY_401 ();
 sky130_fd_sc_hd__decap_3 PHY_402 ();
 sky130_fd_sc_hd__decap_3 PHY_403 ();
 sky130_fd_sc_hd__decap_3 PHY_404 ();
 sky130_fd_sc_hd__decap_3 PHY_405 ();
 sky130_fd_sc_hd__decap_3 PHY_406 ();
 sky130_fd_sc_hd__decap_3 PHY_407 ();
 sky130_fd_sc_hd__decap_3 PHY_408 ();
 sky130_fd_sc_hd__decap_3 PHY_409 ();
 sky130_fd_sc_hd__decap_3 PHY_410 ();
 sky130_fd_sc_hd__decap_3 PHY_411 ();
 sky130_fd_sc_hd__decap_3 PHY_412 ();
 sky130_fd_sc_hd__decap_3 PHY_413 ();
 sky130_fd_sc_hd__decap_3 PHY_414 ();
 sky130_fd_sc_hd__decap_3 PHY_415 ();
 sky130_fd_sc_hd__decap_3 PHY_416 ();
 sky130_fd_sc_hd__decap_3 PHY_417 ();
 sky130_fd_sc_hd__decap_3 PHY_418 ();
 sky130_fd_sc_hd__decap_3 PHY_419 ();
 sky130_fd_sc_hd__decap_3 PHY_420 ();
 sky130_fd_sc_hd__decap_3 PHY_421 ();
 sky130_fd_sc_hd__decap_3 PHY_422 ();
 sky130_fd_sc_hd__decap_3 PHY_423 ();
 sky130_fd_sc_hd__decap_3 PHY_424 ();
 sky130_fd_sc_hd__decap_3 PHY_425 ();
 sky130_fd_sc_hd__decap_3 PHY_426 ();
 sky130_fd_sc_hd__decap_3 PHY_427 ();
 sky130_fd_sc_hd__decap_3 PHY_428 ();
 sky130_fd_sc_hd__decap_3 PHY_429 ();
 sky130_fd_sc_hd__decap_3 PHY_430 ();
 sky130_fd_sc_hd__decap_3 PHY_431 ();
 sky130_fd_sc_hd__decap_3 PHY_432 ();
 sky130_fd_sc_hd__decap_3 PHY_433 ();
 sky130_fd_sc_hd__decap_3 PHY_434 ();
 sky130_fd_sc_hd__decap_3 PHY_435 ();
 sky130_fd_sc_hd__decap_3 PHY_436 ();
 sky130_fd_sc_hd__decap_3 PHY_437 ();
 sky130_fd_sc_hd__decap_3 PHY_438 ();
 sky130_fd_sc_hd__decap_3 PHY_439 ();
 sky130_fd_sc_hd__decap_3 PHY_440 ();
 sky130_fd_sc_hd__decap_3 PHY_441 ();
 sky130_fd_sc_hd__decap_3 PHY_442 ();
 sky130_fd_sc_hd__decap_3 PHY_443 ();
 sky130_fd_sc_hd__decap_3 PHY_444 ();
 sky130_fd_sc_hd__decap_3 PHY_445 ();
 sky130_fd_sc_hd__decap_3 PHY_446 ();
 sky130_fd_sc_hd__decap_3 PHY_447 ();
 sky130_fd_sc_hd__decap_3 PHY_448 ();
 sky130_fd_sc_hd__decap_3 PHY_449 ();
 sky130_fd_sc_hd__decap_3 PHY_450 ();
 sky130_fd_sc_hd__decap_3 PHY_451 ();
 sky130_fd_sc_hd__decap_3 PHY_452 ();
 sky130_fd_sc_hd__decap_3 PHY_453 ();
 sky130_fd_sc_hd__decap_3 PHY_454 ();
 sky130_fd_sc_hd__decap_3 PHY_455 ();
 sky130_fd_sc_hd__decap_3 PHY_456 ();
 sky130_fd_sc_hd__decap_3 PHY_457 ();
 sky130_fd_sc_hd__decap_3 PHY_458 ();
 sky130_fd_sc_hd__decap_3 PHY_459 ();
 sky130_fd_sc_hd__decap_3 PHY_460 ();
 sky130_fd_sc_hd__decap_3 PHY_461 ();
 sky130_fd_sc_hd__decap_3 PHY_462 ();
 sky130_fd_sc_hd__decap_3 PHY_463 ();
 sky130_fd_sc_hd__decap_3 PHY_464 ();
 sky130_fd_sc_hd__decap_3 PHY_465 ();
 sky130_fd_sc_hd__decap_3 PHY_466 ();
 sky130_fd_sc_hd__decap_3 PHY_467 ();
 sky130_fd_sc_hd__decap_3 PHY_468 ();
 sky130_fd_sc_hd__decap_3 PHY_469 ();
 sky130_fd_sc_hd__decap_3 PHY_470 ();
 sky130_fd_sc_hd__decap_3 PHY_471 ();
 sky130_fd_sc_hd__decap_3 PHY_472 ();
 sky130_fd_sc_hd__decap_3 PHY_473 ();
 sky130_fd_sc_hd__decap_3 PHY_474 ();
 sky130_fd_sc_hd__decap_3 PHY_475 ();
 sky130_fd_sc_hd__decap_3 PHY_476 ();
 sky130_fd_sc_hd__decap_3 PHY_477 ();
 sky130_fd_sc_hd__decap_3 PHY_478 ();
 sky130_fd_sc_hd__decap_3 PHY_479 ();
 sky130_fd_sc_hd__decap_3 PHY_480 ();
 sky130_fd_sc_hd__decap_3 PHY_481 ();
 sky130_fd_sc_hd__decap_3 PHY_482 ();
 sky130_fd_sc_hd__decap_3 PHY_483 ();
 sky130_fd_sc_hd__decap_3 PHY_484 ();
 sky130_fd_sc_hd__decap_3 PHY_485 ();
 sky130_fd_sc_hd__decap_3 PHY_486 ();
 sky130_fd_sc_hd__decap_3 PHY_487 ();
 sky130_fd_sc_hd__decap_3 PHY_488 ();
 sky130_fd_sc_hd__decap_3 PHY_489 ();
 sky130_fd_sc_hd__decap_3 PHY_490 ();
 sky130_fd_sc_hd__decap_3 PHY_491 ();
 sky130_fd_sc_hd__decap_3 PHY_492 ();
 sky130_fd_sc_hd__decap_3 PHY_493 ();
 sky130_fd_sc_hd__decap_3 PHY_494 ();
 sky130_fd_sc_hd__decap_3 PHY_495 ();
 sky130_fd_sc_hd__decap_3 PHY_496 ();
 sky130_fd_sc_hd__decap_3 PHY_497 ();
 sky130_fd_sc_hd__decap_3 PHY_498 ();
 sky130_fd_sc_hd__decap_3 PHY_499 ();
 sky130_fd_sc_hd__decap_3 PHY_500 ();
 sky130_fd_sc_hd__decap_3 PHY_501 ();
 sky130_fd_sc_hd__decap_3 PHY_502 ();
 sky130_fd_sc_hd__decap_3 PHY_503 ();
 sky130_fd_sc_hd__decap_3 PHY_504 ();
 sky130_fd_sc_hd__decap_3 PHY_505 ();
 sky130_fd_sc_hd__decap_3 PHY_506 ();
 sky130_fd_sc_hd__decap_3 PHY_507 ();
 sky130_fd_sc_hd__decap_3 PHY_508 ();
 sky130_fd_sc_hd__decap_3 PHY_509 ();
 sky130_fd_sc_hd__decap_3 PHY_510 ();
 sky130_fd_sc_hd__decap_3 PHY_511 ();
 sky130_fd_sc_hd__decap_3 PHY_512 ();
 sky130_fd_sc_hd__decap_3 PHY_513 ();
 sky130_fd_sc_hd__decap_3 PHY_514 ();
 sky130_fd_sc_hd__decap_3 PHY_515 ();
 sky130_fd_sc_hd__decap_3 PHY_516 ();
 sky130_fd_sc_hd__decap_3 PHY_517 ();
 sky130_fd_sc_hd__decap_3 PHY_518 ();
 sky130_fd_sc_hd__decap_3 PHY_519 ();
 sky130_fd_sc_hd__decap_3 PHY_520 ();
 sky130_fd_sc_hd__decap_3 PHY_521 ();
 sky130_fd_sc_hd__decap_3 PHY_522 ();
 sky130_fd_sc_hd__decap_3 PHY_523 ();
 sky130_fd_sc_hd__decap_3 PHY_524 ();
 sky130_fd_sc_hd__decap_3 PHY_525 ();
 sky130_fd_sc_hd__decap_3 PHY_526 ();
 sky130_fd_sc_hd__decap_3 PHY_527 ();
 sky130_fd_sc_hd__decap_3 PHY_528 ();
 sky130_fd_sc_hd__decap_3 PHY_529 ();
 sky130_fd_sc_hd__decap_3 PHY_530 ();
 sky130_fd_sc_hd__decap_3 PHY_531 ();
 sky130_fd_sc_hd__decap_3 PHY_532 ();
 sky130_fd_sc_hd__decap_3 PHY_533 ();
 sky130_fd_sc_hd__decap_3 PHY_534 ();
 sky130_fd_sc_hd__decap_3 PHY_535 ();
 sky130_fd_sc_hd__decap_3 PHY_536 ();
 sky130_fd_sc_hd__decap_3 PHY_537 ();
 sky130_fd_sc_hd__decap_3 PHY_538 ();
 sky130_fd_sc_hd__decap_3 PHY_539 ();
 sky130_fd_sc_hd__decap_3 PHY_540 ();
 sky130_fd_sc_hd__decap_3 PHY_541 ();
 sky130_fd_sc_hd__decap_3 PHY_542 ();
 sky130_fd_sc_hd__decap_3 PHY_543 ();
 sky130_fd_sc_hd__decap_3 PHY_544 ();
 sky130_fd_sc_hd__decap_3 PHY_545 ();
 sky130_fd_sc_hd__decap_3 PHY_546 ();
 sky130_fd_sc_hd__decap_3 PHY_547 ();
 sky130_fd_sc_hd__decap_3 PHY_548 ();
 sky130_fd_sc_hd__decap_3 PHY_549 ();
 sky130_fd_sc_hd__decap_3 PHY_550 ();
 sky130_fd_sc_hd__decap_3 PHY_551 ();
 sky130_fd_sc_hd__decap_3 PHY_552 ();
 sky130_fd_sc_hd__decap_3 PHY_553 ();
 sky130_fd_sc_hd__decap_3 PHY_554 ();
 sky130_fd_sc_hd__decap_3 PHY_555 ();
 sky130_fd_sc_hd__decap_3 PHY_556 ();
 sky130_fd_sc_hd__decap_3 PHY_557 ();
 sky130_fd_sc_hd__decap_3 PHY_558 ();
 sky130_fd_sc_hd__decap_3 PHY_559 ();
 sky130_fd_sc_hd__decap_3 PHY_560 ();
 sky130_fd_sc_hd__decap_3 PHY_561 ();
 sky130_fd_sc_hd__decap_3 PHY_562 ();
 sky130_fd_sc_hd__decap_3 PHY_563 ();
 sky130_fd_sc_hd__decap_3 PHY_564 ();
 sky130_fd_sc_hd__decap_3 PHY_565 ();
 sky130_fd_sc_hd__decap_3 PHY_566 ();
 sky130_fd_sc_hd__decap_3 PHY_567 ();
 sky130_fd_sc_hd__decap_3 PHY_568 ();
 sky130_fd_sc_hd__decap_3 PHY_569 ();
 sky130_fd_sc_hd__decap_3 PHY_570 ();
 sky130_fd_sc_hd__decap_3 PHY_571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4891 ();
 sky130_fd_sc_hd__clkbuf_1 input1 (.A(i_core_int_sreg[0]),
    .X(net1));
 sky130_fd_sc_hd__clkbuf_1 input2 (.A(i_core_int_sreg[10]),
    .X(net2));
 sky130_fd_sc_hd__clkbuf_1 input3 (.A(i_core_int_sreg[11]),
    .X(net3));
 sky130_fd_sc_hd__clkbuf_1 input4 (.A(i_core_int_sreg[12]),
    .X(net4));
 sky130_fd_sc_hd__clkbuf_1 input5 (.A(i_core_int_sreg[13]),
    .X(net5));
 sky130_fd_sc_hd__clkbuf_1 input6 (.A(i_core_int_sreg[14]),
    .X(net6));
 sky130_fd_sc_hd__dlymetal6s2s_1 input7 (.A(i_core_int_sreg[15]),
    .X(net7));
 sky130_fd_sc_hd__clkbuf_1 input8 (.A(i_core_int_sreg[1]),
    .X(net8));
 sky130_fd_sc_hd__clkbuf_1 input9 (.A(i_core_int_sreg[2]),
    .X(net9));
 sky130_fd_sc_hd__clkbuf_1 input10 (.A(i_core_int_sreg[3]),
    .X(net10));
 sky130_fd_sc_hd__clkbuf_1 input11 (.A(i_core_int_sreg[4]),
    .X(net11));
 sky130_fd_sc_hd__dlymetal6s2s_1 input12 (.A(i_core_int_sreg[5]),
    .X(net12));
 sky130_fd_sc_hd__clkbuf_1 input13 (.A(i_core_int_sreg[6]),
    .X(net13));
 sky130_fd_sc_hd__clkbuf_1 input14 (.A(i_core_int_sreg[7]),
    .X(net14));
 sky130_fd_sc_hd__clkbuf_1 input15 (.A(i_core_int_sreg[8]),
    .X(net15));
 sky130_fd_sc_hd__clkbuf_1 input16 (.A(i_core_int_sreg[9]),
    .X(net16));
 sky130_fd_sc_hd__clkbuf_1 input17 (.A(i_disable),
    .X(net17));
 sky130_fd_sc_hd__clkbuf_1 input18 (.A(i_irq),
    .X(net18));
 sky130_fd_sc_hd__clkbuf_1 input19 (.A(i_mc_core_int),
    .X(net19));
 sky130_fd_sc_hd__clkbuf_4 input20 (.A(i_mem_ack),
    .X(net20));
 sky130_fd_sc_hd__buf_2 input21 (.A(i_mem_data[0]),
    .X(net21));
 sky130_fd_sc_hd__clkbuf_1 input22 (.A(i_mem_data[10]),
    .X(net22));
 sky130_fd_sc_hd__clkbuf_2 input23 (.A(i_mem_data[11]),
    .X(net23));
 sky130_fd_sc_hd__dlymetal6s2s_1 input24 (.A(i_mem_data[12]),
    .X(net24));
 sky130_fd_sc_hd__clkbuf_2 input25 (.A(i_mem_data[13]),
    .X(net25));
 sky130_fd_sc_hd__clkbuf_2 input26 (.A(i_mem_data[14]),
    .X(net26));
 sky130_fd_sc_hd__clkbuf_2 input27 (.A(i_mem_data[15]),
    .X(net27));
 sky130_fd_sc_hd__buf_2 input28 (.A(i_mem_data[1]),
    .X(net28));
 sky130_fd_sc_hd__buf_2 input29 (.A(i_mem_data[2]),
    .X(net29));
 sky130_fd_sc_hd__clkbuf_2 input30 (.A(i_mem_data[3]),
    .X(net30));
 sky130_fd_sc_hd__clkbuf_2 input31 (.A(i_mem_data[4]),
    .X(net31));
 sky130_fd_sc_hd__dlymetal6s2s_1 input32 (.A(i_mem_data[5]),
    .X(net32));
 sky130_fd_sc_hd__clkbuf_1 input33 (.A(i_mem_data[6]),
    .X(net33));
 sky130_fd_sc_hd__clkbuf_1 input34 (.A(i_mem_data[7]),
    .X(net34));
 sky130_fd_sc_hd__clkbuf_1 input35 (.A(i_mem_data[8]),
    .X(net35));
 sky130_fd_sc_hd__clkbuf_1 input36 (.A(i_mem_data[9]),
    .X(net36));
 sky130_fd_sc_hd__buf_6 input37 (.A(i_mem_exception),
    .X(net37));
 sky130_fd_sc_hd__clkbuf_1 input38 (.A(i_req_data[0]),
    .X(net38));
 sky130_fd_sc_hd__clkbuf_1 input39 (.A(i_req_data[10]),
    .X(net39));
 sky130_fd_sc_hd__clkbuf_1 input40 (.A(i_req_data[11]),
    .X(net40));
 sky130_fd_sc_hd__clkbuf_1 input41 (.A(i_req_data[12]),
    .X(net41));
 sky130_fd_sc_hd__clkbuf_1 input42 (.A(i_req_data[13]),
    .X(net42));
 sky130_fd_sc_hd__clkbuf_1 input43 (.A(i_req_data[14]),
    .X(net43));
 sky130_fd_sc_hd__clkbuf_1 input44 (.A(i_req_data[15]),
    .X(net44));
 sky130_fd_sc_hd__clkbuf_1 input45 (.A(i_req_data[16]),
    .X(net45));
 sky130_fd_sc_hd__clkbuf_1 input46 (.A(i_req_data[17]),
    .X(net46));
 sky130_fd_sc_hd__dlymetal6s2s_1 input47 (.A(i_req_data[18]),
    .X(net47));
 sky130_fd_sc_hd__dlymetal6s2s_1 input48 (.A(i_req_data[19]),
    .X(net48));
 sky130_fd_sc_hd__clkbuf_1 input49 (.A(i_req_data[1]),
    .X(net49));
 sky130_fd_sc_hd__clkbuf_1 input50 (.A(i_req_data[20]),
    .X(net50));
 sky130_fd_sc_hd__clkbuf_1 input51 (.A(i_req_data[21]),
    .X(net51));
 sky130_fd_sc_hd__clkbuf_1 input52 (.A(i_req_data[22]),
    .X(net52));
 sky130_fd_sc_hd__clkbuf_1 input53 (.A(i_req_data[23]),
    .X(net53));
 sky130_fd_sc_hd__clkbuf_1 input54 (.A(i_req_data[24]),
    .X(net54));
 sky130_fd_sc_hd__clkbuf_1 input55 (.A(i_req_data[25]),
    .X(net55));
 sky130_fd_sc_hd__clkbuf_1 input56 (.A(i_req_data[26]),
    .X(net56));
 sky130_fd_sc_hd__clkbuf_1 input57 (.A(i_req_data[27]),
    .X(net57));
 sky130_fd_sc_hd__clkbuf_1 input58 (.A(i_req_data[28]),
    .X(net58));
 sky130_fd_sc_hd__clkbuf_1 input59 (.A(i_req_data[29]),
    .X(net59));
 sky130_fd_sc_hd__clkbuf_1 input60 (.A(i_req_data[2]),
    .X(net60));
 sky130_fd_sc_hd__clkbuf_1 input61 (.A(i_req_data[30]),
    .X(net61));
 sky130_fd_sc_hd__dlymetal6s2s_1 input62 (.A(i_req_data[31]),
    .X(net62));
 sky130_fd_sc_hd__clkbuf_1 input63 (.A(i_req_data[3]),
    .X(net63));
 sky130_fd_sc_hd__clkbuf_1 input64 (.A(i_req_data[4]),
    .X(net64));
 sky130_fd_sc_hd__clkbuf_1 input65 (.A(i_req_data[5]),
    .X(net65));
 sky130_fd_sc_hd__clkbuf_1 input66 (.A(i_req_data[6]),
    .X(net66));
 sky130_fd_sc_hd__clkbuf_1 input67 (.A(i_req_data[7]),
    .X(net67));
 sky130_fd_sc_hd__clkbuf_1 input68 (.A(i_req_data[8]),
    .X(net68));
 sky130_fd_sc_hd__dlymetal6s2s_1 input69 (.A(i_req_data[9]),
    .X(net69));
 sky130_fd_sc_hd__buf_6 input70 (.A(i_req_data_valid),
    .X(net70));
 sky130_fd_sc_hd__buf_12 input71 (.A(i_rst),
    .X(net71));
 sky130_fd_sc_hd__buf_2 output72 (.A(net211),
    .X(dbg_pc[0]));
 sky130_fd_sc_hd__buf_2 output73 (.A(net73),
    .X(dbg_pc[10]));
 sky130_fd_sc_hd__buf_2 output74 (.A(net74),
    .X(dbg_pc[11]));
 sky130_fd_sc_hd__buf_2 output75 (.A(net75),
    .X(dbg_pc[12]));
 sky130_fd_sc_hd__buf_2 output76 (.A(net76),
    .X(dbg_pc[13]));
 sky130_fd_sc_hd__buf_2 output77 (.A(net77),
    .X(dbg_pc[14]));
 sky130_fd_sc_hd__buf_2 output78 (.A(net78),
    .X(dbg_pc[15]));
 sky130_fd_sc_hd__buf_2 output79 (.A(net79),
    .X(dbg_pc[1]));
 sky130_fd_sc_hd__buf_2 output80 (.A(net80),
    .X(dbg_pc[2]));
 sky130_fd_sc_hd__buf_2 output81 (.A(net81),
    .X(dbg_pc[3]));
 sky130_fd_sc_hd__buf_2 output82 (.A(net82),
    .X(dbg_pc[4]));
 sky130_fd_sc_hd__buf_2 output83 (.A(net83),
    .X(dbg_pc[5]));
 sky130_fd_sc_hd__buf_2 output84 (.A(net84),
    .X(dbg_pc[6]));
 sky130_fd_sc_hd__buf_2 output85 (.A(net85),
    .X(dbg_pc[7]));
 sky130_fd_sc_hd__buf_2 output86 (.A(net86),
    .X(dbg_pc[8]));
 sky130_fd_sc_hd__buf_2 output87 (.A(net87),
    .X(dbg_pc[9]));
 sky130_fd_sc_hd__buf_2 output88 (.A(net88),
    .X(dbg_r0[0]));
 sky130_fd_sc_hd__buf_2 output89 (.A(net89),
    .X(dbg_r0[10]));
 sky130_fd_sc_hd__buf_2 output90 (.A(net90),
    .X(dbg_r0[11]));
 sky130_fd_sc_hd__buf_2 output91 (.A(net91),
    .X(dbg_r0[12]));
 sky130_fd_sc_hd__buf_2 output92 (.A(net92),
    .X(dbg_r0[13]));
 sky130_fd_sc_hd__buf_2 output93 (.A(net93),
    .X(dbg_r0[14]));
 sky130_fd_sc_hd__buf_2 output94 (.A(net94),
    .X(dbg_r0[15]));
 sky130_fd_sc_hd__buf_2 output95 (.A(net95),
    .X(dbg_r0[1]));
 sky130_fd_sc_hd__buf_2 output96 (.A(net96),
    .X(dbg_r0[2]));
 sky130_fd_sc_hd__buf_2 output97 (.A(net97),
    .X(dbg_r0[3]));
 sky130_fd_sc_hd__buf_2 output98 (.A(net98),
    .X(dbg_r0[4]));
 sky130_fd_sc_hd__buf_2 output99 (.A(net99),
    .X(dbg_r0[5]));
 sky130_fd_sc_hd__buf_2 output100 (.A(net100),
    .X(dbg_r0[6]));
 sky130_fd_sc_hd__buf_2 output101 (.A(net101),
    .X(dbg_r0[7]));
 sky130_fd_sc_hd__buf_2 output102 (.A(net102),
    .X(dbg_r0[8]));
 sky130_fd_sc_hd__buf_2 output103 (.A(net103),
    .X(dbg_r0[9]));
 sky130_fd_sc_hd__buf_2 output104 (.A(net104),
    .X(o_c_data_page));
 sky130_fd_sc_hd__buf_2 output105 (.A(net105),
    .X(o_c_instr_long));
 sky130_fd_sc_hd__buf_2 output106 (.A(net106),
    .X(o_c_instr_page));
 sky130_fd_sc_hd__buf_2 output107 (.A(net107),
    .X(o_icache_flush));
 sky130_fd_sc_hd__buf_2 output108 (.A(net108),
    .X(o_instr_long_addr[0]));
 sky130_fd_sc_hd__buf_2 output109 (.A(net109),
    .X(o_instr_long_addr[1]));
 sky130_fd_sc_hd__buf_2 output110 (.A(net110),
    .X(o_instr_long_addr[2]));
 sky130_fd_sc_hd__buf_2 output111 (.A(net111),
    .X(o_instr_long_addr[3]));
 sky130_fd_sc_hd__buf_2 output112 (.A(net112),
    .X(o_instr_long_addr[4]));
 sky130_fd_sc_hd__buf_2 output113 (.A(net113),
    .X(o_instr_long_addr[5]));
 sky130_fd_sc_hd__buf_2 output114 (.A(net114),
    .X(o_instr_long_addr[6]));
 sky130_fd_sc_hd__buf_2 output115 (.A(net115),
    .X(o_instr_long_addr[7]));
 sky130_fd_sc_hd__buf_2 output116 (.A(net116),
    .X(o_mem_addr[0]));
 sky130_fd_sc_hd__buf_2 output117 (.A(net117),
    .X(o_mem_addr[10]));
 sky130_fd_sc_hd__buf_2 output118 (.A(net118),
    .X(o_mem_addr[11]));
 sky130_fd_sc_hd__buf_2 output119 (.A(net119),
    .X(o_mem_addr[12]));
 sky130_fd_sc_hd__buf_2 output120 (.A(net120),
    .X(o_mem_addr[13]));
 sky130_fd_sc_hd__buf_2 output121 (.A(net121),
    .X(o_mem_addr[14]));
 sky130_fd_sc_hd__buf_2 output122 (.A(net122),
    .X(o_mem_addr[15]));
 sky130_fd_sc_hd__buf_2 output123 (.A(net123),
    .X(o_mem_addr[1]));
 sky130_fd_sc_hd__buf_2 output124 (.A(net124),
    .X(o_mem_addr[2]));
 sky130_fd_sc_hd__buf_2 output125 (.A(net125),
    .X(o_mem_addr[3]));
 sky130_fd_sc_hd__buf_2 output126 (.A(net126),
    .X(o_mem_addr[4]));
 sky130_fd_sc_hd__buf_2 output127 (.A(net127),
    .X(o_mem_addr[5]));
 sky130_fd_sc_hd__buf_2 output128 (.A(net128),
    .X(o_mem_addr[6]));
 sky130_fd_sc_hd__buf_2 output129 (.A(net129),
    .X(o_mem_addr[7]));
 sky130_fd_sc_hd__buf_2 output130 (.A(net130),
    .X(o_mem_addr[8]));
 sky130_fd_sc_hd__buf_2 output131 (.A(net131),
    .X(o_mem_addr[9]));
 sky130_fd_sc_hd__buf_2 output132 (.A(net132),
    .X(o_mem_addr_high[0]));
 sky130_fd_sc_hd__buf_2 output133 (.A(net133),
    .X(o_mem_addr_high[1]));
 sky130_fd_sc_hd__buf_2 output134 (.A(net134),
    .X(o_mem_addr_high[2]));
 sky130_fd_sc_hd__buf_2 output135 (.A(net135),
    .X(o_mem_addr_high[3]));
 sky130_fd_sc_hd__buf_2 output136 (.A(net136),
    .X(o_mem_addr_high[4]));
 sky130_fd_sc_hd__buf_2 output137 (.A(net137),
    .X(o_mem_addr_high[5]));
 sky130_fd_sc_hd__buf_2 output138 (.A(net138),
    .X(o_mem_addr_high[6]));
 sky130_fd_sc_hd__buf_2 output139 (.A(net139),
    .X(o_mem_data[0]));
 sky130_fd_sc_hd__buf_2 output140 (.A(net140),
    .X(o_mem_data[10]));
 sky130_fd_sc_hd__buf_2 output141 (.A(net141),
    .X(o_mem_data[11]));
 sky130_fd_sc_hd__buf_2 output142 (.A(net142),
    .X(o_mem_data[12]));
 sky130_fd_sc_hd__buf_2 output143 (.A(net143),
    .X(o_mem_data[13]));
 sky130_fd_sc_hd__buf_2 output144 (.A(net144),
    .X(o_mem_data[14]));
 sky130_fd_sc_hd__buf_2 output145 (.A(net145),
    .X(o_mem_data[15]));
 sky130_fd_sc_hd__buf_2 output146 (.A(net146),
    .X(o_mem_data[1]));
 sky130_fd_sc_hd__buf_2 output147 (.A(net147),
    .X(o_mem_data[2]));
 sky130_fd_sc_hd__buf_2 output148 (.A(net148),
    .X(o_mem_data[3]));
 sky130_fd_sc_hd__buf_2 output149 (.A(net149),
    .X(o_mem_data[4]));
 sky130_fd_sc_hd__buf_2 output150 (.A(net150),
    .X(o_mem_data[5]));
 sky130_fd_sc_hd__buf_2 output151 (.A(net151),
    .X(o_mem_data[6]));
 sky130_fd_sc_hd__buf_2 output152 (.A(net152),
    .X(o_mem_data[7]));
 sky130_fd_sc_hd__buf_2 output153 (.A(net153),
    .X(o_mem_data[8]));
 sky130_fd_sc_hd__buf_2 output154 (.A(net154),
    .X(o_mem_data[9]));
 sky130_fd_sc_hd__buf_2 output155 (.A(net155),
    .X(o_mem_long));
 sky130_fd_sc_hd__buf_2 output156 (.A(net156),
    .X(o_mem_req));
 sky130_fd_sc_hd__buf_2 output157 (.A(net157),
    .X(o_mem_sel[0]));
 sky130_fd_sc_hd__buf_2 output158 (.A(net158),
    .X(o_mem_sel[1]));
 sky130_fd_sc_hd__buf_2 output159 (.A(net159),
    .X(o_mem_we));
 sky130_fd_sc_hd__buf_2 output160 (.A(net160),
    .X(o_req_active));
 sky130_fd_sc_hd__buf_2 output161 (.A(net161),
    .X(o_req_addr[0]));
 sky130_fd_sc_hd__buf_2 output162 (.A(net162),
    .X(o_req_addr[10]));
 sky130_fd_sc_hd__buf_2 output163 (.A(net163),
    .X(o_req_addr[11]));
 sky130_fd_sc_hd__buf_2 output164 (.A(net164),
    .X(o_req_addr[12]));
 sky130_fd_sc_hd__buf_2 output165 (.A(net165),
    .X(o_req_addr[13]));
 sky130_fd_sc_hd__buf_2 output166 (.A(net166),
    .X(o_req_addr[14]));
 sky130_fd_sc_hd__buf_2 output167 (.A(net167),
    .X(o_req_addr[15]));
 sky130_fd_sc_hd__buf_2 output168 (.A(net168),
    .X(o_req_addr[1]));
 sky130_fd_sc_hd__buf_2 output169 (.A(net169),
    .X(o_req_addr[2]));
 sky130_fd_sc_hd__buf_2 output170 (.A(net170),
    .X(o_req_addr[3]));
 sky130_fd_sc_hd__buf_2 output171 (.A(net171),
    .X(o_req_addr[4]));
 sky130_fd_sc_hd__buf_2 output172 (.A(net172),
    .X(o_req_addr[5]));
 sky130_fd_sc_hd__buf_2 output173 (.A(net173),
    .X(o_req_addr[6]));
 sky130_fd_sc_hd__buf_2 output174 (.A(net174),
    .X(o_req_addr[7]));
 sky130_fd_sc_hd__buf_2 output175 (.A(net175),
    .X(o_req_addr[8]));
 sky130_fd_sc_hd__buf_2 output176 (.A(net176),
    .X(o_req_addr[9]));
 sky130_fd_sc_hd__buf_2 output177 (.A(net177),
    .X(o_req_ppl_submit));
 sky130_fd_sc_hd__buf_2 output178 (.A(net178),
    .X(sr_bus_addr[0]));
 sky130_fd_sc_hd__buf_2 output179 (.A(net179),
    .X(sr_bus_addr[10]));
 sky130_fd_sc_hd__buf_2 output180 (.A(net180),
    .X(sr_bus_addr[11]));
 sky130_fd_sc_hd__buf_2 output181 (.A(net181),
    .X(sr_bus_addr[12]));
 sky130_fd_sc_hd__buf_2 output182 (.A(net182),
    .X(sr_bus_addr[13]));
 sky130_fd_sc_hd__buf_2 output183 (.A(net183),
    .X(sr_bus_addr[14]));
 sky130_fd_sc_hd__buf_2 output184 (.A(net184),
    .X(sr_bus_addr[15]));
 sky130_fd_sc_hd__buf_2 output185 (.A(net185),
    .X(sr_bus_addr[1]));
 sky130_fd_sc_hd__buf_2 output186 (.A(net186),
    .X(sr_bus_addr[2]));
 sky130_fd_sc_hd__buf_2 output187 (.A(net187),
    .X(sr_bus_addr[3]));
 sky130_fd_sc_hd__buf_2 output188 (.A(net188),
    .X(sr_bus_addr[4]));
 sky130_fd_sc_hd__buf_2 output189 (.A(net189),
    .X(sr_bus_addr[5]));
 sky130_fd_sc_hd__buf_2 output190 (.A(net190),
    .X(sr_bus_addr[6]));
 sky130_fd_sc_hd__buf_2 output191 (.A(net191),
    .X(sr_bus_addr[7]));
 sky130_fd_sc_hd__buf_2 output192 (.A(net192),
    .X(sr_bus_addr[8]));
 sky130_fd_sc_hd__buf_2 output193 (.A(net193),
    .X(sr_bus_addr[9]));
 sky130_fd_sc_hd__buf_2 output194 (.A(net194),
    .X(sr_bus_data_o[0]));
 sky130_fd_sc_hd__buf_2 output195 (.A(net195),
    .X(sr_bus_data_o[10]));
 sky130_fd_sc_hd__buf_2 output196 (.A(net196),
    .X(sr_bus_data_o[11]));
 sky130_fd_sc_hd__buf_2 output197 (.A(net197),
    .X(sr_bus_data_o[12]));
 sky130_fd_sc_hd__buf_2 output198 (.A(net198),
    .X(sr_bus_data_o[13]));
 sky130_fd_sc_hd__buf_2 output199 (.A(net199),
    .X(sr_bus_data_o[14]));
 sky130_fd_sc_hd__buf_2 output200 (.A(net200),
    .X(sr_bus_data_o[15]));
 sky130_fd_sc_hd__buf_2 output201 (.A(net201),
    .X(sr_bus_data_o[1]));
 sky130_fd_sc_hd__buf_2 output202 (.A(net202),
    .X(sr_bus_data_o[2]));
 sky130_fd_sc_hd__buf_2 output203 (.A(net203),
    .X(sr_bus_data_o[3]));
 sky130_fd_sc_hd__buf_2 output204 (.A(net204),
    .X(sr_bus_data_o[4]));
 sky130_fd_sc_hd__buf_2 output205 (.A(net205),
    .X(sr_bus_data_o[5]));
 sky130_fd_sc_hd__buf_2 output206 (.A(net206),
    .X(sr_bus_data_o[6]));
 sky130_fd_sc_hd__buf_2 output207 (.A(net207),
    .X(sr_bus_data_o[7]));
 sky130_fd_sc_hd__buf_2 output208 (.A(net208),
    .X(sr_bus_data_o[8]));
 sky130_fd_sc_hd__buf_2 output209 (.A(net209),
    .X(sr_bus_data_o[9]));
 sky130_fd_sc_hd__buf_2 output210 (.A(net210),
    .X(sr_bus_we));
 sky130_fd_sc_hd__buf_6 fanout211 (.A(net72),
    .X(net211));
 sky130_fd_sc_hd__conb_1 core1_212 (.LO(net212));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_1_i_clk (.A(clknet_2_0_0_i_clk),
    .X(clknet_leaf_1_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_2_i_clk (.A(clknet_2_0_0_i_clk),
    .X(clknet_leaf_2_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_3_i_clk (.A(clknet_2_0_0_i_clk),
    .X(clknet_leaf_3_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_4_i_clk (.A(clknet_2_0_0_i_clk),
    .X(clknet_leaf_4_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_5_i_clk (.A(clknet_2_2_0_i_clk),
    .X(clknet_leaf_5_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_6_i_clk (.A(clknet_2_2_0_i_clk),
    .X(clknet_leaf_6_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_7_i_clk (.A(clknet_2_2_0_i_clk),
    .X(clknet_leaf_7_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_8_i_clk (.A(clknet_2_2_0_i_clk),
    .X(clknet_leaf_8_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_9_i_clk (.A(clknet_2_2_0_i_clk),
    .X(clknet_leaf_9_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_10_i_clk (.A(clknet_2_2_0_i_clk),
    .X(clknet_leaf_10_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_11_i_clk (.A(clknet_2_2_0_i_clk),
    .X(clknet_leaf_11_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_12_i_clk (.A(clknet_2_2_0_i_clk),
    .X(clknet_leaf_12_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_13_i_clk (.A(clknet_2_2_0_i_clk),
    .X(clknet_leaf_13_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_14_i_clk (.A(clknet_2_2_0_i_clk),
    .X(clknet_leaf_14_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_15_i_clk (.A(clknet_2_2_0_i_clk),
    .X(clknet_leaf_15_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_16_i_clk (.A(clknet_2_3_0_i_clk),
    .X(clknet_leaf_16_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_17_i_clk (.A(clknet_2_3_0_i_clk),
    .X(clknet_leaf_17_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_18_i_clk (.A(clknet_2_3_0_i_clk),
    .X(clknet_leaf_18_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_19_i_clk (.A(clknet_2_3_0_i_clk),
    .X(clknet_leaf_19_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_20_i_clk (.A(clknet_2_3_0_i_clk),
    .X(clknet_leaf_20_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_21_i_clk (.A(clknet_2_3_0_i_clk),
    .X(clknet_leaf_21_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_22_i_clk (.A(clknet_2_3_0_i_clk),
    .X(clknet_leaf_22_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_23_i_clk (.A(clknet_opt_2_1_i_clk),
    .X(clknet_leaf_23_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_24_i_clk (.A(clknet_2_3_0_i_clk),
    .X(clknet_leaf_24_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_25_i_clk (.A(clknet_2_3_0_i_clk),
    .X(clknet_leaf_25_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_26_i_clk (.A(clknet_2_3_0_i_clk),
    .X(clknet_leaf_26_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_27_i_clk (.A(clknet_2_3_0_i_clk),
    .X(clknet_leaf_27_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_28_i_clk (.A(clknet_2_3_0_i_clk),
    .X(clknet_leaf_28_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_29_i_clk (.A(clknet_2_3_0_i_clk),
    .X(clknet_leaf_29_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_30_i_clk (.A(clknet_2_3_0_i_clk),
    .X(clknet_leaf_30_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_31_i_clk (.A(clknet_2_1_0_i_clk),
    .X(clknet_leaf_31_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_32_i_clk (.A(clknet_2_1_0_i_clk),
    .X(clknet_leaf_32_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_33_i_clk (.A(clknet_2_1_0_i_clk),
    .X(clknet_leaf_33_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_34_i_clk (.A(clknet_2_1_0_i_clk),
    .X(clknet_leaf_34_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_35_i_clk (.A(clknet_2_1_0_i_clk),
    .X(clknet_leaf_35_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_36_i_clk (.A(clknet_2_1_0_i_clk),
    .X(clknet_leaf_36_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_37_i_clk (.A(clknet_2_1_0_i_clk),
    .X(clknet_leaf_37_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_38_i_clk (.A(clknet_2_1_0_i_clk),
    .X(clknet_leaf_38_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_39_i_clk (.A(clknet_2_1_0_i_clk),
    .X(clknet_leaf_39_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_40_i_clk (.A(clknet_2_1_0_i_clk),
    .X(clknet_leaf_40_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_41_i_clk (.A(clknet_2_1_0_i_clk),
    .X(clknet_leaf_41_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_42_i_clk (.A(clknet_2_1_0_i_clk),
    .X(clknet_leaf_42_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_43_i_clk (.A(clknet_2_1_0_i_clk),
    .X(clknet_leaf_43_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_44_i_clk (.A(clknet_2_0_0_i_clk),
    .X(clknet_leaf_44_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_45_i_clk (.A(clknet_2_1_0_i_clk),
    .X(clknet_leaf_45_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_46_i_clk (.A(clknet_2_1_0_i_clk),
    .X(clknet_leaf_46_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_47_i_clk (.A(clknet_2_0_0_i_clk),
    .X(clknet_leaf_47_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_48_i_clk (.A(clknet_opt_1_1_i_clk),
    .X(clknet_leaf_48_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_49_i_clk (.A(clknet_2_0_0_i_clk),
    .X(clknet_leaf_49_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_50_i_clk (.A(clknet_2_0_0_i_clk),
    .X(clknet_leaf_50_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_i_clk (.A(i_clk),
    .X(clknet_0_i_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_1_0_0_i_clk (.A(clknet_0_i_clk),
    .X(clknet_1_0_0_i_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_1_0_1_i_clk (.A(clknet_1_0_0_i_clk),
    .X(clknet_1_0_1_i_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_1_1_0_i_clk (.A(clknet_0_i_clk),
    .X(clknet_1_1_0_i_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_1_1_1_i_clk (.A(clknet_1_1_0_i_clk),
    .X(clknet_1_1_1_i_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_2_0_0_i_clk (.A(clknet_1_0_1_i_clk),
    .X(clknet_2_0_0_i_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_2_1_0_i_clk (.A(clknet_1_0_1_i_clk),
    .X(clknet_2_1_0_i_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_2_2_0_i_clk (.A(clknet_1_1_1_i_clk),
    .X(clknet_2_2_0_i_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_2_3_0_i_clk (.A(clknet_1_1_1_i_clk),
    .X(clknet_2_3_0_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_opt_1_0_i_clk (.A(clknet_2_0_0_i_clk),
    .X(clknet_opt_1_0_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_opt_1_1_i_clk (.A(clknet_opt_1_0_i_clk),
    .X(clknet_opt_1_1_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_opt_2_0_i_clk (.A(clknet_2_3_0_i_clk),
    .X(clknet_opt_2_0_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_opt_2_1_i_clk (.A(clknet_opt_2_0_i_clk),
    .X(clknet_opt_2_1_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6784__D (.DIODE(_0015_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3893__B1 (.DIODE(_0015_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3887__B1 (.DIODE(_0015_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3882__B1 (.DIODE(_0015_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3874__B1 (.DIODE(_0015_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3858__B1 (.DIODE(_0015_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3855__B1 (.DIODE(_0015_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3844__B1 (.DIODE(_0015_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3825__B1 (.DIODE(_0015_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3818__B1 (.DIODE(_0015_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6792__D (.DIODE(_0023_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6793__D (.DIODE(_0024_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6794__D (.DIODE(_0025_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6884__D (.DIODE(_0115_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7013__D (.DIODE(_0228_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5666__C1 (.DIODE(_0228_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5159__B1_N (.DIODE(_0228_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3520__B (.DIODE(_0519_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3512__B (.DIODE(_0519_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3505__A2 (.DIODE(_0519_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3482__B1 (.DIODE(_0519_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3474__B (.DIODE(_0519_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3466__B (.DIODE(_0519_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3458__B1 (.DIODE(_0519_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3450__B (.DIODE(_0519_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3418__B1 (.DIODE(_0519_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3365__A (.DIODE(_0519_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4418__A2 (.DIODE(_0520_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4414__A2 (.DIODE(_0520_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4401__A2 (.DIODE(_0520_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4396__A2 (.DIODE(_0520_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3496__B1 (.DIODE(_0520_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3443__A2 (.DIODE(_0520_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3434__A2 (.DIODE(_0520_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3425__B1 (.DIODE(_0520_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3402__A2 (.DIODE(_0520_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3390__A2 (.DIODE(_0520_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3516__A2 (.DIODE(_0521_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3488__A2 (.DIODE(_0521_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3481__A2 (.DIODE(_0521_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3473__A2 (.DIODE(_0521_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3457__A2 (.DIODE(_0521_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3417__A2 (.DIODE(_0521_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3367__A (.DIODE(_0521_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3511__A2 (.DIODE(_0522_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3499__A2 (.DIODE(_0522_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3495__A2 (.DIODE(_0522_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3465__A2 (.DIODE(_0522_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3449__A2 (.DIODE(_0522_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3442__A2 (.DIODE(_0522_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3433__A2 (.DIODE(_0522_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3424__A2 (.DIODE(_0522_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3394__A2 (.DIODE(_0522_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3376__A2 (.DIODE(_0522_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3518__D (.DIODE(_0523_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3517__B (.DIODE(_0523_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3472__C (.DIODE(_0523_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3460__A (.DIODE(_0523_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3414__B (.DIODE(_0523_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3413__A_N (.DIODE(_0523_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3392__A (.DIODE(_0523_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3387__A (.DIODE(_0523_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3374__A (.DIODE(_0523_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3371__A_N (.DIODE(_0523_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3516__B1 (.DIODE(_0526_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3508__A2 (.DIODE(_0526_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3492__A2 (.DIODE(_0526_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3469__A2 (.DIODE(_0526_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3462__A2 (.DIODE(_0526_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3394__B1 (.DIODE(_0526_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3376__B1 (.DIODE(_0526_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3441__B (.DIODE(_0527_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3440__C (.DIODE(_0527_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3436__B (.DIODE(_0527_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3429__B_N (.DIODE(_0527_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3423__C (.DIODE(_0527_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3422__B (.DIODE(_0527_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3398__B (.DIODE(_0527_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3397__B_N (.DIODE(_0527_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3388__B_N (.DIODE(_0527_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3375__A_N (.DIODE(_0527_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3502__D (.DIODE(_0528_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3498__C (.DIODE(_0528_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3494__A_N (.DIODE(_0528_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3448__C (.DIODE(_0528_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3432__D (.DIODE(_0528_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3431__C (.DIODE(_0528_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3427__B (.DIODE(_0528_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3388__C (.DIODE(_0528_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3386__A_N (.DIODE(_0528_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3375__B (.DIODE(_0528_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4046__A1 (.DIODE(_0532_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3557__S1 (.DIODE(_0532_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3555__S1 (.DIODE(_0532_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3464__B (.DIODE(_0532_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3463__A_N (.DIODE(_0532_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3438__A_N (.DIODE(_0532_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3437__B_N (.DIODE(_0532_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3399__C (.DIODE(_0532_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3393__A_N (.DIODE(_0532_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3379__A (.DIODE(_0532_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4044__A1 (.DIODE(_0533_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3557__S0 (.DIODE(_0533_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3555__S0 (.DIODE(_0533_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3464__A_N (.DIODE(_0533_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3463__B_N (.DIODE(_0533_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3438__B (.DIODE(_0533_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3399__D (.DIODE(_0533_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3398__A_N (.DIODE(_0533_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3393__B (.DIODE(_0533_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3379__B (.DIODE(_0533_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3504__A1 (.DIODE(_0534_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3400__A1 (.DIODE(_0534_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3389__A1 (.DIODE(_0534_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3510__B (.DIODE(_0536_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3509__C (.DIODE(_0536_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3501__D (.DIODE(_0536_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3494__C (.DIODE(_0536_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3493__B (.DIODE(_0536_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3480__B (.DIODE(_0536_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3479__A_N (.DIODE(_0536_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3447__B (.DIODE(_0536_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3386__C (.DIODE(_0536_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3384__B (.DIODE(_0536_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3518__A_N (.DIODE(_0537_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3517__C (.DIODE(_0537_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3510__C (.DIODE(_0537_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3509__B (.DIODE(_0537_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3494__B (.DIODE(_0537_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3493__C (.DIODE(_0537_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3480__C (.DIODE(_0537_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3479__B (.DIODE(_0537_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3447__C (.DIODE(_0537_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3384__C (.DIODE(_0537_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3518__B (.DIODE(_0538_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3517__D (.DIODE(_0538_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3510__D (.DIODE(_0538_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3509__A_N (.DIODE(_0538_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3501__B (.DIODE(_0538_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3493__D (.DIODE(_0538_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3480__D (.DIODE(_0538_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3479__C (.DIODE(_0538_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3447__D (.DIODE(_0538_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3384__D (.DIODE(_0538_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3503__B (.DIODE(_0540_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3502__C (.DIODE(_0540_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3501__A_N (.DIODE(_0540_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3498__B (.DIODE(_0540_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3448__B (.DIODE(_0540_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3432__C (.DIODE(_0540_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3431__B (.DIODE(_0540_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3428__B (.DIODE(_0540_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3427__A_N (.DIODE(_0540_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3386__B (.DIODE(_0540_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3498__A_N (.DIODE(_0542_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3463__D (.DIODE(_0542_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3440__B (.DIODE(_0542_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3436__C (.DIODE(_0542_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3429__A_N (.DIODE(_0542_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3423__B (.DIODE(_0542_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3422__A_N (.DIODE(_0542_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3398__C (.DIODE(_0542_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3397__A_N (.DIODE(_0542_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3388__A_N (.DIODE(_0542_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6632__A (.DIODE(_0545_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3391__A (.DIODE(_0545_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4049__A1 (.DIODE(_0546_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3559__A1 (.DIODE(_0546_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3556__A (.DIODE(_0546_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3464__C (.DIODE(_0546_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3441__A_N (.DIODE(_0546_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3438__D (.DIODE(_0546_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3437__A_N (.DIODE(_0546_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3399__B (.DIODE(_0546_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3395__B_N (.DIODE(_0546_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3393__D (.DIODE(_0546_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3503__A_N (.DIODE(_0550_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3441__C (.DIODE(_0550_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3440__D (.DIODE(_0550_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3437__C (.DIODE(_0550_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3436__A_N (.DIODE(_0550_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3429__C (.DIODE(_0550_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3428__A_N (.DIODE(_0550_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3423__D (.DIODE(_0550_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3422__C (.DIODE(_0550_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3397__C (.DIODE(_0550_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6628__A (.DIODE(_0556_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6495__A1 (.DIODE(_0556_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3403__A (.DIODE(_0556_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3485__A2 (.DIODE(_0557_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3453__A2 (.DIODE(_0557_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3405__A (.DIODE(_0557_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3515__A2 (.DIODE(_0558_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3508__B1 (.DIODE(_0558_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3499__B1 (.DIODE(_0558_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3492__B1 (.DIODE(_0558_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3478__A2 (.DIODE(_0558_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3469__B1 (.DIODE(_0558_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3462__B1 (.DIODE(_0558_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3446__A2 (.DIODE(_0558_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3420__A2 (.DIODE(_0558_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3407__A2 (.DIODE(_0558_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3515__B1 (.DIODE(_0559_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3485__B1 (.DIODE(_0559_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3478__B1 (.DIODE(_0559_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3453__B1 (.DIODE(_0559_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3446__B1 (.DIODE(_0559_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3420__B1 (.DIODE(_0559_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3407__B1 (.DIODE(_0559_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3507__A2 (.DIODE(_0562_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3491__A2 (.DIODE(_0562_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3484__A2 (.DIODE(_0562_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3477__A2 (.DIODE(_0562_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3470__A2 (.DIODE(_0562_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3461__A2 (.DIODE(_0562_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3454__A2 (.DIODE(_0562_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3445__A2 (.DIODE(_0562_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3421__A2 (.DIODE(_0562_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3412__A2 (.DIODE(_0562_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3519__A2 (.DIODE(_0564_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3507__B1 (.DIODE(_0564_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3491__B1 (.DIODE(_0564_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3477__B1 (.DIODE(_0564_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3454__B1 (.DIODE(_0564_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3445__B1 (.DIODE(_0564_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3439__A2 (.DIODE(_0564_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3430__A2 (.DIODE(_0564_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3421__B1 (.DIODE(_0564_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3412__B1 (.DIODE(_0564_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3519__D1 (.DIODE(_0569_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3511__D1 (.DIODE(_0569_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3495__D1 (.DIODE(_0569_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3481__D1 (.DIODE(_0569_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3465__D1 (.DIODE(_0569_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3449__D1 (.DIODE(_0569_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3442__D1 (.DIODE(_0569_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3433__D1 (.DIODE(_0569_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3424__D1 (.DIODE(_0569_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3417__D1 (.DIODE(_0569_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6624__A (.DIODE(_0571_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4406__A1 (.DIODE(_0571_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3419__A (.DIODE(_0571_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6619__A (.DIODE(_0577_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6483__A1 (.DIODE(_0577_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5665__B (.DIODE(_0577_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4409__A2 (.DIODE(_0577_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3426__A (.DIODE(_0577_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6615__A (.DIODE(_0585_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5637__A2 (.DIODE(_0585_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3435__A (.DIODE(_0585_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6611__A (.DIODE(_0593_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3444__A (.DIODE(_0593_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6607__A (.DIODE(_0600_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6465__A1 (.DIODE(_0600_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4423__A2 (.DIODE(_0600_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3452__A (.DIODE(_0600_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6603__A (.DIODE(_0606_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3459__A (.DIODE(_0606_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3470__B1 (.DIODE(_0607_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3461__B1 (.DIODE(_0607_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6781__A1 (.DIODE(_0614_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6599__A (.DIODE(_0614_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4793__A2 (.DIODE(_0614_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4429__A2 (.DIODE(_0614_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3468__A (.DIODE(_0614_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3475__A3 (.DIODE(_0619_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6778__A1 (.DIODE(_0621_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6595__A (.DIODE(_0621_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6446__A (.DIODE(_0621_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3476__A (.DIODE(_0621_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6775__A1 (.DIODE(_0627_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6591__A (.DIODE(_0627_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6439__A (.DIODE(_0627_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4792__A2 (.DIODE(_0627_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4437__A2 (.DIODE(_0627_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3483__A (.DIODE(_0627_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6772__A1 (.DIODE(_0633_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6733__A (.DIODE(_0633_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6587__A (.DIODE(_0633_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5401__A1 (.DIODE(_0633_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4444__A1 (.DIODE(_0633_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3490__A (.DIODE(_0633_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4785__A2 (.DIODE(_0639_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3497__A (.DIODE(_0639_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6766__A1 (.DIODE(_0647_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6577__A (.DIODE(_0647_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6423__B1 (.DIODE(_0647_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4463__A1 (.DIODE(_0647_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3506__A (.DIODE(_0647_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3514__A (.DIODE(_0654_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6760__A1 (.DIODE(_0661_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3522__A (.DIODE(_0661_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5931__A (.DIODE(_0662_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5157__A (.DIODE(_0662_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5137__A (.DIODE(_0662_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4973__A (.DIODE(_0662_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4385__A (.DIODE(_0662_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4282__B (.DIODE(_0662_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3991__A (.DIODE(_0662_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3896__A (.DIODE(_0662_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3644__A (.DIODE(_0662_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3683__A1 (.DIODE(_0664_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3676__A1 (.DIODE(_0664_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3659__A1 (.DIODE(_0664_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3628__A1 (.DIODE(_0664_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3615__A1 (.DIODE(_0664_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3612__S (.DIODE(_0664_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3611__S (.DIODE(_0664_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3604__S (.DIODE(_0664_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3603__S (.DIODE(_0664_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3526__A (.DIODE(_0664_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3703__S (.DIODE(_0665_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3702__S (.DIODE(_0665_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3701__S (.DIODE(_0665_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3650__A1 (.DIODE(_0665_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3640__S (.DIODE(_0665_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3607__S (.DIODE(_0665_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3606__S (.DIODE(_0665_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3602__S (.DIODE(_0665_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3601__S (.DIODE(_0665_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3527__A (.DIODE(_0665_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4392__S (.DIODE(_0666_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4342__S (.DIODE(_0666_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4339__S (.DIODE(_0666_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4336__S (.DIODE(_0666_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4333__S (.DIODE(_0666_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4330__S (.DIODE(_0666_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4273__B1 (.DIODE(_0666_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3947__A1 (.DIODE(_0666_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3704__S (.DIODE(_0666_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3642__A1 (.DIODE(_0666_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6646__A (.DIODE(_0670_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6636__A (.DIODE(_0670_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6563__B1 (.DIODE(_0670_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6561__B1 (.DIODE(_0670_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6415__B (.DIODE(_0670_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4779__B1 (.DIODE(_0670_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4144__B (.DIODE(_0670_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4141__A (.DIODE(_0670_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3985__C1 (.DIODE(_0670_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3551__A (.DIODE(_0670_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6755__A1 (.DIODE(_0671_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6704__A (.DIODE(_0671_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6701__A1 (.DIODE(_0671_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6699__A (.DIODE(_0671_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6652__B2 (.DIODE(_0671_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5283__B2 (.DIODE(_0671_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3546__B (.DIODE(_0671_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3538__B (.DIODE(_0671_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3534__B (.DIODE(_0671_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3533__B (.DIODE(_0671_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6766__A0 (.DIODE(_0672_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4963__B (.DIODE(_0672_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3791__A (.DIODE(_0672_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3541__B1 (.DIODE(_0672_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3537__A2 (.DIODE(_0672_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6781__A0 (.DIODE(_0673_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4968__B (.DIODE(_0673_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3796__A (.DIODE(_0673_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3537__B1 (.DIODE(_0673_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3536__A2_N (.DIODE(_0673_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6778__A0 (.DIODE(_0677_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4967__B (.DIODE(_0677_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3795__A (.DIODE(_0677_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3541__A2 (.DIODE(_0677_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3540__A2_N (.DIODE(_0677_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6775__A0 (.DIODE(_0681_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4966__B (.DIODE(_0681_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3794__A (.DIODE(_0681_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3543__B (.DIODE(_0681_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3988__C1 (.DIODE(_0689_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3551__B (.DIODE(_0689_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4959__D (.DIODE(_0692_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4957__D (.DIODE(_0692_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4922__A (.DIODE(_0692_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3599__A (.DIODE(_0692_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3598__C (.DIODE(_0692_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4742__B (.DIODE(_0699_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4726__B_N (.DIODE(_0699_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4717__A_N (.DIODE(_0699_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4716__B (.DIODE(_0699_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4715__B (.DIODE(_0699_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4704__B (.DIODE(_0699_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4648__A (.DIODE(_0699_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4647__C_N (.DIODE(_0699_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4613__A (.DIODE(_0699_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3561__A (.DIODE(_0699_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4692__A2 (.DIODE(_0701_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4685__B (.DIODE(_0701_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4679__B (.DIODE(_0701_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4669__B (.DIODE(_0701_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4634__A2 (.DIODE(_0701_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4615__A2 (.DIODE(_0701_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4609__A (.DIODE(_0701_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3585__C1 (.DIODE(_0701_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3580__A1 (.DIODE(_0701_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3577__A (.DIODE(_0701_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4749__C (.DIODE(_0702_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4742__C (.DIODE(_0702_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4716__A_N (.DIODE(_0702_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4706__C (.DIODE(_0702_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4705__B (.DIODE(_0702_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4704__A_N (.DIODE(_0702_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4647__A (.DIODE(_0702_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4613__B (.DIODE(_0702_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3582__A (.DIODE(_0702_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3565__A (.DIODE(_0702_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4756__A (.DIODE(_0703_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4725__B1 (.DIODE(_0703_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4718__B1 (.DIODE(_0703_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4707__B1 (.DIODE(_0703_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4647__B (.DIODE(_0703_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4628__A2 (.DIODE(_0703_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4618__C (.DIODE(_0703_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3582__B_N (.DIODE(_0703_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3568__A (.DIODE(_0703_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3565__B (.DIODE(_0703_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4749__B (.DIODE(_0706_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4733__B (.DIODE(_0706_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4706__B (.DIODE(_0706_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4705__A_N (.DIODE(_0706_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4644__B (.DIODE(_0706_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4618__A (.DIODE(_0706_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4617__A (.DIODE(_0706_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4036__A1 (.DIODE(_0706_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3588__C1 (.DIODE(_0706_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3576__A (.DIODE(_0706_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4751__B2 (.DIODE(_0707_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4744__A (.DIODE(_0707_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4738__B2 (.DIODE(_0707_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4693__A2 (.DIODE(_0707_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4680__A2 (.DIODE(_0707_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4653__B (.DIODE(_0707_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4650__A1 (.DIODE(_0707_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4635__A2 (.DIODE(_0707_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4616__A2 (.DIODE(_0707_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3569__A (.DIODE(_0707_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4819__B2 (.DIODE(_0708_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4683__A2 (.DIODE(_0708_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4671__B (.DIODE(_0708_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4032__A1 (.DIODE(_0708_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3586__A (.DIODE(_0708_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3583__A (.DIODE(_0708_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3581__B (.DIODE(_0708_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3578__S0 (.DIODE(_0708_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3575__B2 (.DIODE(_0708_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3572__A_N (.DIODE(_0708_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4733__C (.DIODE(_0710_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4644__C (.DIODE(_0710_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4618__B (.DIODE(_0710_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4034__A1 (.DIODE(_0710_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3586__C_N (.DIODE(_0710_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3583__C_N (.DIODE(_0710_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3581__A (.DIODE(_0710_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3578__S1 (.DIODE(_0710_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3574__A (.DIODE(_0710_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3572__C (.DIODE(_0710_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4727__B2 (.DIODE(_0712_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4692__B1 (.DIODE(_0712_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4686__B2 (.DIODE(_0712_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4680__B2 (.DIODE(_0712_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4672__B2 (.DIODE(_0712_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4656__B2 (.DIODE(_0712_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4634__B1 (.DIODE(_0712_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4628__B2 (.DIODE(_0712_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4615__B1 (.DIODE(_0712_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3575__A2 (.DIODE(_0712_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4609__B (.DIODE(_0721_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3587__B1 (.DIODE(_0721_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3584__B1 (.DIODE(_0721_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4959__B (.DIODE(_0729_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4957__B (.DIODE(_0729_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4920__A (.DIODE(_0729_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3995__B (.DIODE(_0729_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3598__A (.DIODE(_0729_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6360__B (.DIODE(_0731_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4917__S (.DIODE(_0731_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4390__B (.DIODE(_0731_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3597__B (.DIODE(_0731_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5752__B1_N (.DIODE(_0732_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5721__B1_N (.DIODE(_0732_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5582__B1_N (.DIODE(_0732_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5548__B1_N (.DIODE(_0732_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5365__B1_N (.DIODE(_0732_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5336__B1_N (.DIODE(_0732_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5292__B1_N (.DIODE(_0732_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4487__A (.DIODE(_0732_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3594__B (.DIODE(_0732_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6273__B1 (.DIODE(_0734_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6199__A (.DIODE(_0734_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6184__A (.DIODE(_0734_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6181__A (.DIODE(_0734_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3596__B (.DIODE(_0734_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4910__A (.DIODE(_0735_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4904__A (.DIODE(_0735_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4202__A1 (.DIODE(_0735_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4200__B (.DIODE(_0735_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3597__C (.DIODE(_0735_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4959__C (.DIODE(_0736_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4957__C (.DIODE(_0736_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4921__A (.DIODE(_0736_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3995__C (.DIODE(_0736_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3598__B (.DIODE(_0736_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6756__A (.DIODE(_0737_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6635__C (.DIODE(_0737_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4776__A (.DIODE(_0737_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4774__A (.DIODE(_0737_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3984__A (.DIODE(_0737_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3981__B1 (.DIODE(_0737_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3951__A (.DIODE(_0737_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3599__B (.DIODE(_0737_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4274__C (.DIODE(_0739_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4204__B (.DIODE(_0739_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3947__B1 (.DIODE(_0739_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3642__B1 (.DIODE(_0739_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4319__A0 (.DIODE(_0740_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3706__B (.DIODE(_0740_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3641__A (.DIODE(_0740_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4317__A0 (.DIODE(_0741_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3706__C (.DIODE(_0741_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3641__B (.DIODE(_0741_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4307__A0 (.DIODE(_0742_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3616__D_N (.DIODE(_0742_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3605__A (.DIODE(_0742_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4309__A0 (.DIODE(_0743_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3707__D_N (.DIODE(_0743_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3616__A (.DIODE(_0743_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3605__B_N (.DIODE(_0743_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4311__A0 (.DIODE(_0745_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3638__B1 (.DIODE(_0745_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3608__A (.DIODE(_0745_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4313__A0 (.DIODE(_0746_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3638__C1 (.DIODE(_0746_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3608__B (.DIODE(_0746_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4362__A0 (.DIODE(_0749_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3755__A1 (.DIODE(_0749_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3651__A (.DIODE(_0749_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3637__A (.DIODE(_0749_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4366__A0 (.DIODE(_0750_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3746__A1 (.DIODE(_0750_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3668__B1 (.DIODE(_0750_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3655__B1 (.DIODE(_0750_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3637__B (.DIODE(_0750_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4347__A0 (.DIODE(_0751_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3784__A1 (.DIODE(_0751_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3692__B (.DIODE(_0751_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3679__B (.DIODE(_0751_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3678__A2 (.DIODE(_0751_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3616__B (.DIODE(_0751_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4351__A0 (.DIODE(_0754_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3776__A1 (.DIODE(_0754_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3616__C (.DIODE(_0754_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4360__A0 (.DIODE(_0756_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3760__A1 (.DIODE(_0756_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3686__B1 (.DIODE(_0756_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3672__B (.DIODE(_0756_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3622__A (.DIODE(_0756_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4354__A0 (.DIODE(_0759_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3772__A1 (.DIODE(_0759_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3690__B1 (.DIODE(_0759_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3685__B1 (.DIODE(_0759_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3622__C (.DIODE(_0759_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4374__A0 (.DIODE(_0760_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3732__A1 (.DIODE(_0760_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3662__B2 (.DIODE(_0760_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3658__B1 (.DIODE(_0760_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3622__D (.DIODE(_0760_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4370__A0 (.DIODE(_0765_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3739__A1 (.DIODE(_0765_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3629__C (.DIODE(_0765_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4376__A0 (.DIODE(_0767_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3713__A1 (.DIODE(_0767_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3629__D (.DIODE(_0767_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4358__A0 (.DIODE(_0769_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3764__A1 (.DIODE(_0769_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3686__A2 (.DIODE(_0769_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3682__A2 (.DIODE(_0769_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3635__A (.DIODE(_0769_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4368__A0 (.DIODE(_0770_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3743__A1 (.DIODE(_0770_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3668__A2 (.DIODE(_0770_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3667__B2 (.DIODE(_0770_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3635__B (.DIODE(_0770_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4364__A0 (.DIODE(_0772_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3751__A1 (.DIODE(_0772_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3635__C (.DIODE(_0772_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4372__A0 (.DIODE(_0773_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3735__A1 (.DIODE(_0773_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3697__A2 (.DIODE(_0773_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3664__A2 (.DIODE(_0773_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3658__A2 (.DIODE(_0773_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3635__D (.DIODE(_0773_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4315__A0 (.DIODE(_0779_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3707__A (.DIODE(_0779_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3641__D_N (.DIODE(_0779_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4303__A1 (.DIODE(_0784_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4302__A1 (.DIODE(_0784_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4301__A1 (.DIODE(_0784_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4300__A1 (.DIODE(_0784_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4293__S (.DIODE(_0784_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4290__S (.DIODE(_0784_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4283__S (.DIODE(_0784_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4276__S (.DIODE(_0784_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3646__A (.DIODE(_0784_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4902__A (.DIODE(_0785_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4274__A (.DIODE(_0785_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4201__A (.DIODE(_0785_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4134__A (.DIODE(_0785_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3994__A (.DIODE(_0785_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3946__A (.DIODE(_0785_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3801__A (.DIODE(_0785_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3798__A (.DIODE(_0785_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3711__B (.DIODE(_0785_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3648__B (.DIODE(_0785_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4287__A (.DIODE(_0819_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3690__A1 (.DIODE(_0819_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3682__B2 (.DIODE(_0819_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4285__A (.DIODE(_0822_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3690__B2 (.DIODE(_0822_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3685__B2 (.DIODE(_0822_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3708__A1 (.DIODE(_0838_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4323__A0 (.DIODE(_0839_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3705__A1 (.DIODE(_0839_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4321__A0 (.DIODE(_0840_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3705__A2 (.DIODE(_0840_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4325__A0 (.DIODE(_0842_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3705__A4 (.DIODE(_0842_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3906__A1 (.DIODE(_0846_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3754__A1 (.DIODE(_0846_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3750__A1 (.DIODE(_0846_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3745__B1_N (.DIODE(_0846_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3734__B1_N (.DIODE(_0846_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3709__A (.DIODE(_0846_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4117__B (.DIODE(_0912_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4064__C (.DIODE(_0912_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4062__B (.DIODE(_0912_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4060__B (.DIODE(_0912_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4055__B (.DIODE(_0912_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4001__A2 (.DIODE(_0912_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3898__A2 (.DIODE(_0912_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3895__A (.DIODE(_0912_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3799__B (.DIODE(_0912_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4125__B1 (.DIODE(_0913_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4074__B1 (.DIODE(_0913_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4073__B1 (.DIODE(_0913_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4072__B1 (.DIODE(_0913_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4047__A (.DIODE(_0913_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3890__A (.DIODE(_0913_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3847__A (.DIODE(_0913_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3800__A (.DIODE(_0913_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4127__B1 (.DIODE(_0914_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4076__B1 (.DIODE(_0914_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3887__A2 (.DIODE(_0914_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3882__A2 (.DIODE(_0914_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3874__A2 (.DIODE(_0914_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3858__A2 (.DIODE(_0914_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3855__A2 (.DIODE(_0914_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3844__A2 (.DIODE(_0914_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3825__A2 (.DIODE(_0914_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3818__A2 (.DIODE(_0914_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3999__B (.DIODE(_0915_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3998__A (.DIODE(_0915_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3802__B (.DIODE(_0915_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4915__S (.DIODE(_0916_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4108__S (.DIODE(_0916_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4106__S (.DIODE(_0916_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4085__A (.DIODE(_0916_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3845__A (.DIODE(_0916_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3803__A (.DIODE(_0916_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4128__A (.DIODE(_0921_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4037__A (.DIODE(_0921_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4020__B1 (.DIODE(_0921_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4018__A (.DIODE(_0921_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3998__C (.DIODE(_0921_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3903__A (.DIODE(_0921_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3901__A (.DIODE(_0921_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3854__A2 (.DIODE(_0921_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3824__B1 (.DIODE(_0921_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3810__A (.DIODE(_0921_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3894__A (.DIODE(_0925_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3891__A (.DIODE(_0925_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3885__A (.DIODE(_0925_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3884__A (.DIODE(_0925_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3872__A (.DIODE(_0925_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3871__A_N (.DIODE(_0925_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3867__A (.DIODE(_0925_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3857__A_N (.DIODE(_0925_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3840__A (.DIODE(_0925_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3816__A (.DIODE(_0925_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5738__B2 (.DIODE(_0931_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5654__A1 (.DIODE(_0931_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5556__B2 (.DIODE(_0931_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5521__A1 (.DIODE(_0931_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5503__A1 (.DIODE(_0931_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5463__B2 (.DIODE(_0931_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5430__B2 (.DIODE(_0931_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5382__B2 (.DIODE(_0931_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5311__A1 (.DIODE(_0931_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3825__A1 (.DIODE(_0931_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4050__D (.DIODE(_0932_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4028__B2 (.DIODE(_0932_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3862__A (.DIODE(_0932_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3860__A (.DIODE(_0932_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3850__A1 (.DIODE(_0932_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3834__B (.DIODE(_0932_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3821__B (.DIODE(_0932_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5736__B1 (.DIODE(_0937_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5652__A1 (.DIODE(_0937_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5554__A1 (.DIODE(_0937_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5519__A1 (.DIODE(_0937_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5502__A1 (.DIODE(_0937_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5462__A1 (.DIODE(_0937_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5429__A1 (.DIODE(_0937_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5339__A1 (.DIODE(_0937_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5316__A1 (.DIODE(_0937_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3844__A1 (.DIODE(_0937_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4074__A3 (.DIODE(_0940_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4073__A3 (.DIODE(_0940_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4072__A3 (.DIODE(_0940_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4071__A3 (.DIODE(_0940_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3838__A (.DIODE(_0940_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4132__B1 (.DIODE(_0955_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4131__B1 (.DIODE(_0955_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4129__B1 (.DIODE(_0955_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4125__A1 (.DIODE(_0955_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4123__B1 (.DIODE(_0955_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4121__B1 (.DIODE(_0955_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4114__B1 (.DIODE(_0955_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4113__B1 (.DIODE(_0955_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3889__A2 (.DIODE(_0955_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3850__A2 (.DIODE(_0955_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4040__B (.DIODE(_0956_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4026__A (.DIODE(_0956_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3889__A3 (.DIODE(_0956_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3850__A3 (.DIODE(_0956_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4132__A2 (.DIODE(_0957_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4131__A2 (.DIODE(_0957_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4129__A2 (.DIODE(_0957_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4123__A2 (.DIODE(_0957_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4121__A2 (.DIODE(_0957_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4120__A2 (.DIODE(_0957_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4114__A2 (.DIODE(_0957_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4071__B1 (.DIODE(_0957_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3889__B1 (.DIODE(_0957_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3850__B1 (.DIODE(_0957_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5750__A1 (.DIODE(_0958_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5719__A1 (.DIODE(_0958_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5600__A1 (.DIODE(_0958_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5506__A1 (.DIODE(_0958_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5468__A1 (.DIODE(_0958_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5433__A1 (.DIODE(_0958_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5385__A1 (.DIODE(_0958_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5219__A (.DIODE(_0958_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4784__A (.DIODE(_0958_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3849__A (.DIODE(_0958_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6180__A (.DIODE(_0959_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6162__B (.DIODE(_0959_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5692__A1 (.DIODE(_0959_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5661__A1 (.DIODE(_0959_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5627__A1 (.DIODE(_0959_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5626__A (.DIODE(_0959_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5528__A1 (.DIODE(_0959_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5359__A1 (.DIODE(_0959_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4892__A1 (.DIODE(_0959_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3850__B2 (.DIODE(_0959_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5737__A1 (.DIODE(_0960_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5652__B2 (.DIODE(_0960_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5554__C1 (.DIODE(_0960_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5520__A1 (.DIODE(_0960_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5502__C1 (.DIODE(_0960_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5463__A1 (.DIODE(_0960_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5430__A1 (.DIODE(_0960_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5339__C1 (.DIODE(_0960_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5316__B2 (.DIODE(_0960_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3855__A1 (.DIODE(_0960_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5693__A2 (.DIODE(_0964_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5662__A2 (.DIODE(_0964_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5628__A2 (.DIODE(_0964_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5529__A2 (.DIODE(_0964_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5508__A2 (.DIODE(_0964_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5470__A2 (.DIODE(_0964_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5435__A2 (.DIODE(_0964_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5360__A2 (.DIODE(_0964_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4893__A2 (.DIODE(_0964_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3858__A1 (.DIODE(_0964_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4040__C (.DIODE(_0965_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4029__A (.DIODE(_0965_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3858__B2 (.DIODE(_0965_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5746__B1 (.DIODE(_0966_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5689__A1 (.DIODE(_0966_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5611__B1 (.DIODE(_0966_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5598__C (.DIODE(_0966_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5458__B1 (.DIODE(_0966_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5420__B1 (.DIODE(_0966_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5342__B2 (.DIODE(_0966_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5313__A1_N (.DIODE(_0966_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5092__C1 (.DIODE(_0966_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3874__A1 (.DIODE(_0966_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4132__B2 (.DIODE(_0979_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4130__A2 (.DIODE(_0979_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4112__A (.DIODE(_0979_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4028__B1 (.DIODE(_0979_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4025__A2 (.DIODE(_0979_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4008__C (.DIODE(_0979_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3873__D (.DIODE(_0979_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6532__A1 (.DIODE(_0981_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6531__A (.DIODE(_0981_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5690__A1 (.DIODE(_0981_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5624__A (.DIODE(_0981_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5599__A1 (.DIODE(_0981_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5566__A1 (.DIODE(_0981_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5342__A1 (.DIODE(_0981_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5134__A1 (.DIODE(_0981_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4888__A1 (.DIODE(_0981_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3882__A1 (.DIODE(_0981_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5303__A1 (.DIODE(_0988_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5302__A1 (.DIODE(_0988_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5301__A1 (.DIODE(_0988_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5111__A1 (.DIODE(_0988_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4853__A1 (.DIODE(_0988_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4851__A (.DIODE(_0988_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4845__A1 (.DIODE(_0988_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4836__A1 (.DIODE(_0988_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4831__B (.DIODE(_0988_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3887__A1 (.DIODE(_0988_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5692__C1 (.DIODE(_0992_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5661__C1 (.DIODE(_0992_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5627__C1 (.DIODE(_0992_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5569__C1 (.DIODE(_0992_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5528__C1 (.DIODE(_0992_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5359__C1 (.DIODE(_0992_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5321__C1 (.DIODE(_0992_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5218__A2 (.DIODE(_0992_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4892__C1 (.DIODE(_0992_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3889__B2 (.DIODE(_0992_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4046__A2 (.DIODE(_0993_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4044__A2 (.DIODE(_0993_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4036__A2 (.DIODE(_0993_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4034__A2 (.DIODE(_0993_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4032__A2 (.DIODE(_0993_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4024__A2 (.DIODE(_0993_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4023__A2 (.DIODE(_0993_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4014__A2 (.DIODE(_0993_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3905__A2 (.DIODE(_0993_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3893__A2 (.DIODE(_0993_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4017__C_N (.DIODE(_0996_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3895__B (.DIODE(_0996_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6711__A (.DIODE(_0998_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6672__A (.DIODE(_0998_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6621__A (.DIODE(_0998_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6580__A (.DIODE(_0998_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4971__B (.DIODE(_0998_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4969__B (.DIODE(_0998_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4168__A (.DIODE(_0998_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4066__A (.DIODE(_0998_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4000__A (.DIODE(_0998_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3897__A (.DIODE(_0998_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6783__A (.DIODE(_0999_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6695__B1 (.DIODE(_0999_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4940__C1 (.DIODE(_0999_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4937__C1 (.DIODE(_0999_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4932__C1 (.DIODE(_0999_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4928__C1 (.DIODE(_0999_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4926__C1 (.DIODE(_0999_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4924__C1 (.DIODE(_0999_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4901__B1 (.DIODE(_0999_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3898__C1 (.DIODE(_0999_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5653__B2 (.DIODE(_1000_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5556__A1 (.DIODE(_1000_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5517__A (.DIODE(_1000_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5504__A1 (.DIODE(_1000_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5465__A1 (.DIODE(_1000_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5431__A1 (.DIODE(_1000_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5382__A1 (.DIODE(_1000_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5339__B2 (.DIODE(_1000_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5317__A1 (.DIODE(_1000_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3905__A1 (.DIODE(_1000_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4049__B1 (.DIODE(_1001_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4046__B1 (.DIODE(_1001_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4044__B1 (.DIODE(_1001_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4036__B1 (.DIODE(_1001_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4034__B1 (.DIODE(_1001_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4032__B1 (.DIODE(_1001_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4024__B1 (.DIODE(_1001_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4023__B1 (.DIODE(_1001_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4014__B1 (.DIODE(_1001_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3905__B1 (.DIODE(_1001_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5855__S (.DIODE(_1007_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5850__S (.DIODE(_1007_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5845__S (.DIODE(_1007_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5840__S (.DIODE(_1007_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5835__S (.DIODE(_1007_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5830__S (.DIODE(_1007_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3909__A (.DIODE(_1007_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5824__S (.DIODE(_1008_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5817__S (.DIODE(_1008_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3941__S (.DIODE(_1008_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3939__S (.DIODE(_1008_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3937__S (.DIODE(_1008_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3935__S (.DIODE(_1008_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3933__S (.DIODE(_1008_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3931__S (.DIODE(_1008_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3929__S (.DIODE(_1008_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3910__A (.DIODE(_1008_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3940__A (.DIODE(_1023_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3942__A (.DIODE(_1024_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3944__A (.DIODE(_1025_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4376__S (.DIODE(_1027_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4374__S (.DIODE(_1027_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4353__A (.DIODE(_1027_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4327__A (.DIODE(_1027_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4306__A (.DIODE(_1027_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3948__A (.DIODE(_1027_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3950__A (.DIODE(_1028_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6709__A (.DIODE(_1029_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6702__A (.DIODE(_1029_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6511__B1 (.DIODE(_1029_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6159__A2 (.DIODE(_1029_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5137__B (.DIODE(_1029_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4973__B (.DIODE(_1029_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4930__A (.DIODE(_1029_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4900__A (.DIODE(_1029_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4771__A2 (.DIODE(_1029_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3952__A (.DIODE(_1029_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4948__A2 (.DIODE(_1030_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4946__A2 (.DIODE(_1030_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4944__A2 (.DIODE(_1030_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4940__A2 (.DIODE(_1030_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4937__A2 (.DIODE(_1030_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4932__A2 (.DIODE(_1030_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4928__A2 (.DIODE(_1030_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4926__A2 (.DIODE(_1030_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4924__A2 (.DIODE(_1030_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3990__A1 (.DIODE(_1030_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5209__B (.DIODE(_1050_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5206__B (.DIODE(_1050_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4463__A0 (.DIODE(_1050_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3974__B (.DIODE(_1050_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5209__C (.DIODE(_1051_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5206__C (.DIODE(_1051_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5202__C (.DIODE(_1051_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5197__C (.DIODE(_1051_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3984__B (.DIODE(_1051_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3974__C (.DIODE(_1051_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5198__B (.DIODE(_1053_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5194__C (.DIODE(_1053_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4135__C (.DIODE(_1053_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3984__C (.DIODE(_1053_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3977__C (.DIODE(_1053_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5198__C (.DIODE(_1054_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5194__D (.DIODE(_1054_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4135__D (.DIODE(_1054_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3977__D (.DIODE(_1054_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6505__A2 (.DIODE(_1057_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6411__A (.DIODE(_1057_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5702__B (.DIODE(_1057_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5672__B (.DIODE(_1057_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5642__B (.DIODE(_1057_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5579__B (.DIODE(_1057_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4780__A (.DIODE(_1057_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4140__A (.DIODE(_1057_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4126__A (.DIODE(_1057_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3980__B1 (.DIODE(_1057_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6704__B (.DIODE(_1059_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6699__B (.DIODE(_1059_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6652__A2 (.DIODE(_1059_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6649__A2 (.DIODE(_1059_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6646__B (.DIODE(_1059_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3986__B (.DIODE(_1059_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3985__A2 (.DIODE(_1059_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3984__D (.DIODE(_1061_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3985__B1 (.DIODE(_1062_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3992__B (.DIODE(_1066_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3989__B1 (.DIODE(_1066_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3990__A2 (.DIODE(_1067_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6698__A3 (.DIODE(_1068_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4934__B1 (.DIODE(_1068_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4166__A (.DIODE(_1068_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4163__A (.DIODE(_1068_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4160__A (.DIODE(_1068_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4157__A (.DIODE(_1068_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4154__A (.DIODE(_1068_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4151__A (.DIODE(_1068_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4148__A (.DIODE(_1068_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3992__A (.DIODE(_1068_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6655__B (.DIODE(_1071_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6563__A1 (.DIODE(_1071_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6561__A1 (.DIODE(_1071_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5157__B (.DIODE(_1071_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4971__C (.DIODE(_1071_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4969__C (.DIODE(_1071_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4935__A2 (.DIODE(_1071_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4133__B (.DIODE(_1071_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3996__C (.DIODE(_1071_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4127__A2_N (.DIODE(_1073_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4001__B1 (.DIODE(_1073_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4076__A2_N (.DIODE(_1074_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4001__C1 (.DIODE(_1074_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6780__C1 (.DIODE(_1075_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6777__C1 (.DIODE(_1075_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6774__C1 (.DIODE(_1075_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6771__C1 (.DIODE(_1075_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6697__A2 (.DIODE(_1075_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6696__A2 (.DIODE(_1075_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6692__A3 (.DIODE(_1075_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4120__B2 (.DIODE(_1075_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4118__C1 (.DIODE(_1075_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4001__D1 (.DIODE(_1075_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4797__A1 (.DIODE(_1076_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4796__A1 (.DIODE(_1076_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4437__A1 (.DIODE(_1076_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4436__A (.DIODE(_1076_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4428__A (.DIODE(_1076_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4423__A1 (.DIODE(_1076_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4422__A (.DIODE(_1076_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4409__A1 (.DIODE(_1076_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4408__A (.DIODE(_1076_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4003__A (.DIODE(_1076_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4995__A1 (.DIODE(_1077_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4978__A1 (.DIODE(_1077_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4793__A1 (.DIODE(_1077_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4792__A1 (.DIODE(_1077_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4785__A1 (.DIODE(_1077_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4448__A1 (.DIODE(_1077_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4429__A1 (.DIODE(_1077_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4415__A1 (.DIODE(_1077_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4397__A1 (.DIODE(_1077_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4014__A1 (.DIODE(_1077_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4030__A (.DIODE(_1095_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4023__B2 (.DIODE(_1095_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4118__A1 (.DIODE(_1096_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4038__B (.DIODE(_1096_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4035__A2 (.DIODE(_1096_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4033__A2 (.DIODE(_1096_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4031__A2 (.DIODE(_1096_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4035__B1 (.DIODE(_1101_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4033__B1 (.DIODE(_1101_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4031__B1 (.DIODE(_1101_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4119__A1 (.DIODE(_1107_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4048__A2 (.DIODE(_1107_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4045__A2 (.DIODE(_1107_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4043__A2 (.DIODE(_1107_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4119__A2 (.DIODE(_1110_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4118__A2 (.DIODE(_1110_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4048__B1 (.DIODE(_1110_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4045__B1 (.DIODE(_1110_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4043__B1 (.DIODE(_1110_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4113__A2 (.DIODE(_1113_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4070__A2 (.DIODE(_1113_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4069__A2 (.DIODE(_1113_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4068__A2 (.DIODE(_1113_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4067__A2 (.DIODE(_1113_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4065__A2 (.DIODE(_1113_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4063__A2 (.DIODE(_1113_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4061__A2 (.DIODE(_1113_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4059__A2 (.DIODE(_1113_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4049__A2 (.DIODE(_1113_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4064__D (.DIODE(_1118_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4062__C (.DIODE(_1118_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4054__B (.DIODE(_1118_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6536__B1 (.DIODE(_1121_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4292__B (.DIODE(_1121_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4289__B (.DIODE(_1121_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4287__B (.DIODE(_1121_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4285__B (.DIODE(_1121_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4280__A (.DIODE(_1121_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4278__B (.DIODE(_1121_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4275__B (.DIODE(_1121_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4075__A (.DIODE(_1121_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4057__A (.DIODE(_1121_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6753__C1 (.DIODE(_1122_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6648__B1 (.DIODE(_1122_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6558__A (.DIODE(_1122_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4968__A (.DIODE(_1122_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4967__A (.DIODE(_1122_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4383__A (.DIODE(_1122_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4378__A (.DIODE(_1122_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4274__B (.DIODE(_1122_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4134__B (.DIODE(_1122_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4058__A (.DIODE(_1122_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6360__A (.DIODE(_1128_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5813__A (.DIODE(_1128_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4966__A (.DIODE(_1128_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4965__A (.DIODE(_1128_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4964__A (.DIODE(_1128_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4963__A (.DIODE(_1128_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4962__A (.DIODE(_1128_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4961__A (.DIODE(_1128_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4127__A1_N (.DIODE(_1128_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4076__A1_N (.DIODE(_1128_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4104__S (.DIODE(_1133_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4102__S (.DIODE(_1133_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4100__S (.DIODE(_1133_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4098__S (.DIODE(_1133_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4096__S (.DIODE(_1133_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4094__S (.DIODE(_1133_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4092__S (.DIODE(_1133_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4090__S (.DIODE(_1133_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4088__S (.DIODE(_1133_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4086__S (.DIODE(_1133_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5755__S (.DIODE(_1146_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5725__S (.DIODE(_1146_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5695__S (.DIODE(_1146_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5604__S (.DIODE(_1146_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5572__S (.DIODE(_1146_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5538__S (.DIODE(_1146_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5510__S (.DIODE(_1146_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5472__S (.DIODE(_1146_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5437__S (.DIODE(_1146_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4111__A (.DIODE(_1146_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5807__A0 (.DIODE(_1147_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5666__A1 (.DIODE(_1147_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5665__A (.DIODE(_1147_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5637__A1 (.DIODE(_1147_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5636__C1 (.DIODE(_1147_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5362__S (.DIODE(_1147_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5324__S (.DIODE(_1147_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5278__S (.DIODE(_1147_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5257__S (.DIODE(_1147_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4113__A1 (.DIODE(_1147_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4113__B2 (.DIODE(_1148_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6754__A (.DIODE(_1153_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6707__A (.DIODE(_1153_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6655__A (.DIODE(_1153_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6635__B (.DIODE(_1153_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6559__A (.DIODE(_1153_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6411__B (.DIODE(_1153_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6410__B (.DIODE(_1153_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4896__B (.DIODE(_1153_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4780__B (.DIODE(_1153_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4123__A1 (.DIODE(_1153_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6479__A2 (.DIODE(_1155_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6459__A2 (.DIODE(_1155_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6447__A2 (.DIODE(_1155_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6440__A2 (.DIODE(_1155_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6435__A2 (.DIODE(_1155_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6430__A2 (.DIODE(_1155_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6423__A2 (.DIODE(_1155_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6161__A1 (.DIODE(_1155_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6159__A1 (.DIODE(_1155_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4127__B2 (.DIODE(_1155_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5444__A2 (.DIODE(_1161_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5407__A2 (.DIODE(_1161_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5393__A2 (.DIODE(_1161_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5328__A2 (.DIODE(_1161_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5287__B1 (.DIODE(_1161_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5270__A2 (.DIODE(_1161_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4138__A (.DIODE(_1161_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5730__A2 (.DIODE(_1162_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5700__A2 (.DIODE(_1162_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5670__A2 (.DIODE(_1162_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5640__A2 (.DIODE(_1162_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5631__A2 (.DIODE(_1162_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5577__A2 (.DIODE(_1162_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5543__A2 (.DIODE(_1162_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5532__A2 (.DIODE(_1162_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5480__A2 (.DIODE(_1162_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4139__B (.DIODE(_1162_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4187__A2 (.DIODE(_1164_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4184__A2 (.DIODE(_1164_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4181__A2 (.DIODE(_1164_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4178__A2 (.DIODE(_1164_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4175__A2 (.DIODE(_1164_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4143__A (.DIODE(_1164_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4141__B (.DIODE(_1164_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4187__B1 (.DIODE(_1165_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4184__B1 (.DIODE(_1165_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4181__B1 (.DIODE(_1165_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4178__B1 (.DIODE(_1165_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4175__B1 (.DIODE(_1165_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4142__A (.DIODE(_1165_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4172__B1 (.DIODE(_1166_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4169__B1 (.DIODE(_1166_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4165__B1 (.DIODE(_1166_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4162__B1 (.DIODE(_1166_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4159__B1 (.DIODE(_1166_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4156__B1 (.DIODE(_1166_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4153__B1 (.DIODE(_1166_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4150__B1 (.DIODE(_1166_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4147__B1 (.DIODE(_1166_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4146__A2 (.DIODE(_1166_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4172__A2 (.DIODE(_1167_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4169__A2 (.DIODE(_1167_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4165__A2 (.DIODE(_1167_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4162__A2 (.DIODE(_1167_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4159__A2 (.DIODE(_1167_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4156__A2 (.DIODE(_1167_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4153__A2 (.DIODE(_1167_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4150__A2 (.DIODE(_1167_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4147__A2 (.DIODE(_1167_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4145__A2 (.DIODE(_1167_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6529__A (.DIODE(_1184_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6525__A (.DIODE(_1184_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4918__A (.DIODE(_1184_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4188__A (.DIODE(_1184_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4185__A (.DIODE(_1184_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4182__A (.DIODE(_1184_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4179__A (.DIODE(_1184_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4176__A (.DIODE(_1184_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4173__A (.DIODE(_1184_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4170__A (.DIODE(_1184_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6315__A1 (.DIODE(_1199_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6301__B1 (.DIODE(_1199_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6290__B1 (.DIODE(_1199_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6267__A1 (.DIODE(_1199_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6244__A (.DIODE(_1199_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6239__A1 (.DIODE(_1199_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6238__B (.DIODE(_1199_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6214__A1 (.DIODE(_1199_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4702__A (.DIODE(_1199_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4191__A (.DIODE(_1199_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6387__A (.DIODE(_1200_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6384__A1 (.DIODE(_1200_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6353__A1 (.DIODE(_1200_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6178__A1 (.DIODE(_1200_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6173__A1 (.DIODE(_1200_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6171__B1 (.DIODE(_1200_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4914__A1 (.DIODE(_1200_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4912__A (.DIODE(_1200_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4495__A (.DIODE(_1200_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4198__A (.DIODE(_1200_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6404__A (.DIODE(_1202_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6401__A1 (.DIODE(_1202_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6382__A (.DIODE(_1202_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6379__A1 (.DIODE(_1202_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6278__A1 (.DIODE(_1202_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6267__A2 (.DIODE(_1202_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6255__S (.DIODE(_1202_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6173__C1 (.DIODE(_1202_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4764__S (.DIODE(_1202_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4197__A (.DIODE(_1202_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6376__B (.DIODE(_1205_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6176__A1 (.DIODE(_1205_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6174__A1 (.DIODE(_1205_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4197__B (.DIODE(_1205_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4594__A (.DIODE(_1207_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4569__A (.DIODE(_1207_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4556__A (.DIODE(_1207_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4528__A (.DIODE(_1207_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4504__A (.DIODE(_1207_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4493__A1 (.DIODE(_1207_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4199__A (.DIODE(_1207_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4602__A1 (.DIODE(_1208_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4588__A1 (.DIODE(_1208_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4581__A1 (.DIODE(_1208_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4580__A (.DIODE(_1208_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4563__A1 (.DIODE(_1208_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4551__A1 (.DIODE(_1208_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4536__A1 (.DIODE(_1208_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4523__A1 (.DIODE(_1208_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4489__A1 (.DIODE(_1208_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4202__A2 (.DIODE(_1208_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4910__B (.DIODE(_1210_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4202__B1_N (.DIODE(_1210_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4304__S (.DIODE(_1213_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4271__S (.DIODE(_1213_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4269__S (.DIODE(_1213_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4248__A (.DIODE(_1213_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4227__A (.DIODE(_1213_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4206__A (.DIODE(_1213_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4225__S (.DIODE(_1214_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4223__S (.DIODE(_1214_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4221__S (.DIODE(_1214_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4219__S (.DIODE(_1214_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4217__S (.DIODE(_1214_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4215__S (.DIODE(_1214_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4213__S (.DIODE(_1214_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4211__S (.DIODE(_1214_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4209__S (.DIODE(_1214_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4207__S (.DIODE(_1214_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4246__S (.DIODE(_1225_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4244__S (.DIODE(_1225_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4242__S (.DIODE(_1225_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4240__S (.DIODE(_1225_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4238__S (.DIODE(_1225_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4236__S (.DIODE(_1225_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4234__S (.DIODE(_1225_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4232__S (.DIODE(_1225_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4230__S (.DIODE(_1225_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4228__S (.DIODE(_1225_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4381__B (.DIODE(_1262_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4303__B1 (.DIODE(_1262_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4302__B1 (.DIODE(_1262_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4301__B1 (.DIODE(_1262_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4300__B1 (.DIODE(_1262_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4299__B1 (.DIODE(_1262_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4298__B1 (.DIODE(_1262_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4297__B1 (.DIODE(_1262_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4296__B1 (.DIODE(_1262_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4325__S (.DIODE(_1264_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4323__S (.DIODE(_1264_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4321__S (.DIODE(_1264_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4319__S (.DIODE(_1264_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4317__S (.DIODE(_1264_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4315__S (.DIODE(_1264_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4313__S (.DIODE(_1264_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4311__S (.DIODE(_1264_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4309__S (.DIODE(_1264_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4307__S (.DIODE(_1264_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4351__S (.DIODE(_1275_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4349__S (.DIODE(_1275_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4347__S (.DIODE(_1275_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4345__S (.DIODE(_1275_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4343__S (.DIODE(_1275_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4340__S (.DIODE(_1275_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4337__S (.DIODE(_1275_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4334__S (.DIODE(_1275_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4331__S (.DIODE(_1275_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4328__S (.DIODE(_1275_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6653__A (.DIODE(_1307_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6650__A (.DIODE(_1307_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6644__A (.DIODE(_1307_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6641__A (.DIODE(_1307_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6638__A (.DIODE(_1307_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5909__A (.DIODE(_1307_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5877__A (.DIODE(_1307_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5828__A (.DIODE(_1307_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4943__A (.DIODE(_1307_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4390__A (.DIODE(_1307_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5861__B (.DIODE(_1309_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5856__S (.DIODE(_1309_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5851__S (.DIODE(_1309_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5846__S (.DIODE(_1309_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5841__S (.DIODE(_1309_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5836__S (.DIODE(_1309_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5831__S (.DIODE(_1309_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5825__S (.DIODE(_1309_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5818__S (.DIODE(_1309_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4388__A (.DIODE(_1309_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5892__B2 (.DIODE(_1310_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5888__B2 (.DIODE(_1310_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5884__B2 (.DIODE(_1310_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5880__B2 (.DIODE(_1310_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5875__B2 (.DIODE(_1310_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5872__B2 (.DIODE(_1310_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5868__B2 (.DIODE(_1310_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5864__B2 (.DIODE(_1310_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5807__A1 (.DIODE(_1310_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4389__A1 (.DIODE(_1310_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4393__A1 (.DIODE(_1313_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4458__C1 (.DIODE(_1315_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4455__C1 (.DIODE(_1315_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4440__S (.DIODE(_1315_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4426__S (.DIODE(_1315_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4400__A (.DIODE(_1315_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4396__C1 (.DIODE(_1315_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4978__B1 (.DIODE(_1316_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4796__B1 (.DIODE(_1316_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4397__B1 (.DIODE(_1316_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6166__B (.DIODE(_1317_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5151__A (.DIODE(_1317_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5091__A (.DIODE(_1317_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4980__A (.DIODE(_1317_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4485__B (.DIODE(_1317_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4398__B (.DIODE(_1317_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4795__S (.DIODE(_1320_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4463__S (.DIODE(_1320_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4451__S (.DIODE(_1320_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4447__A (.DIODE(_1320_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4444__S (.DIODE(_1320_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4431__S (.DIODE(_1320_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4418__C1 (.DIODE(_1320_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4414__C1 (.DIODE(_1320_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4406__S (.DIODE(_1320_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4401__C1 (.DIODE(_1320_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4796__D1 (.DIODE(_1321_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4402__B (.DIODE(_1321_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6169__A1 (.DIODE(_1323_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5713__A2 (.DIODE(_1323_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4985__A (.DIODE(_1323_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4984__A (.DIODE(_1323_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4481__B (.DIODE(_1323_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4404__A (.DIODE(_1323_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5067__A1 (.DIODE(_1326_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4990__A (.DIODE(_1326_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4988__A (.DIODE(_1326_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4987__A (.DIODE(_1326_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4482__B (.DIODE(_1326_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4407__B (.DIODE(_1326_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6168__B (.DIODE(_1329_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5652__A2 (.DIODE(_1329_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5060__A (.DIODE(_1329_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5059__A (.DIODE(_1329_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4798__B (.DIODE(_1329_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4410__A (.DIODE(_1329_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4995__B1 (.DIODE(_1334_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4797__B1 (.DIODE(_1334_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4415__B1 (.DIODE(_1334_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5063__A1 (.DIODE(_1335_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4478__B (.DIODE(_1335_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4416__B (.DIODE(_1335_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4797__D1 (.DIODE(_1338_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4419__B (.DIODE(_1338_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6176__B1 (.DIODE(_1340_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5591__A2 (.DIODE(_1340_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5052__A (.DIODE(_1340_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5051__A (.DIODE(_1340_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4474__B (.DIODE(_1340_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4421__A (.DIODE(_1340_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5001__A (.DIODE(_1341_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5000__A1 (.DIODE(_1341_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4477__A2 (.DIODE(_1341_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6177__B2 (.DIODE(_1343_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5554__A2 (.DIODE(_1343_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5055__A (.DIODE(_1343_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5054__A1 (.DIODE(_1343_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5005__A (.DIODE(_1343_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5004__A (.DIODE(_1343_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4794__A (.DIODE(_1343_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4560__B (.DIODE(_1343_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4475__B_N (.DIODE(_1343_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4424__A_N (.DIODE(_1343_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6177__A2 (.DIODE(_1347_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5519__A2 (.DIODE(_1347_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5517__B (.DIODE(_1347_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5044__A (.DIODE(_1347_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5043__A (.DIODE(_1347_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5008__A (.DIODE(_1347_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5007__A1 (.DIODE(_1347_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4794__B (.DIODE(_1347_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4473__A2 (.DIODE(_1347_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4471__B (.DIODE(_1347_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6171__A2 (.DIODE(_1349_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5047__A (.DIODE(_1349_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5046__A1 (.DIODE(_1349_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4547__B (.DIODE(_1349_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4469__B (.DIODE(_1349_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4430__B (.DIODE(_1349_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6172__A1 (.DIODE(_1351_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5462__A2 (.DIODE(_1351_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5018__A (.DIODE(_1351_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5017__A (.DIODE(_1351_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5015__B1 (.DIODE(_1351_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4794__D (.DIODE(_1351_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4432__A (.DIODE(_1351_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5080__A (.DIODE(_1352_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5013__A1 (.DIODE(_1352_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4434__B (.DIODE(_1352_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4433__B (.DIODE(_1352_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5023__A (.DIODE(_1357_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5021__A1 (.DIODE(_1357_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4853__B1 (.DIODE(_1357_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4840__B (.DIODE(_1357_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4467__B (.DIODE(_1357_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4438__B (.DIODE(_1357_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6170__A2 (.DIODE(_1361_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5381__A2 (.DIODE(_1361_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5244__A (.DIODE(_1361_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5034__A (.DIODE(_1361_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4852__A (.DIODE(_1361_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4832__A (.DIODE(_1361_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4442__B (.DIODE(_1361_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4532__B1 (.DIODE(_1362_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4468__B1 (.DIODE(_1362_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4446__A (.DIODE(_1362_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5380__A1 (.DIODE(_1364_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5082__A (.DIODE(_1364_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5025__A (.DIODE(_1364_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5024__A1 (.DIODE(_1364_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4839__B1 (.DIODE(_1364_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4445__B (.DIODE(_1364_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5031__A (.DIODE(_1368_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5030__A (.DIODE(_1368_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4839__A1 (.DIODE(_1368_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4449__A (.DIODE(_1368_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5460__A (.DIODE(_1369_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5374__A1 (.DIODE(_1369_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5356__A (.DIODE(_1369_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5296__A (.DIODE(_1369_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5248__A1 (.DIODE(_1369_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5245__A (.DIODE(_1369_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4856__A (.DIODE(_1369_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4518__B (.DIODE(_1369_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4462__B (.DIODE(_1369_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4450__B (.DIODE(_1369_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5426__A (.DIODE(_1372_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5355__A1 (.DIODE(_1372_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5354__A (.DIODE(_1372_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5246__A1 (.DIODE(_1372_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5225__A (.DIODE(_1372_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5029__A (.DIODE(_1372_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5027__A (.DIODE(_1372_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4860__A (.DIODE(_1372_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4830__B (.DIODE(_1372_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4453__B (.DIODE(_1372_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4825__A (.DIODE(_1374_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4801__A (.DIODE(_1374_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4786__A (.DIODE(_1374_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4460__B (.DIODE(_1374_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4456__A1 (.DIODE(_1374_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4825__B (.DIODE(_1375_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4801__B (.DIODE(_1375_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4786__B (.DIODE(_1375_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4460__C (.DIODE(_1375_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4456__A2 (.DIODE(_1375_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4874__A1 (.DIODE(_1377_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4873__A (.DIODE(_1377_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4866__A1 (.DIODE(_1377_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4825__C (.DIODE(_1377_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4788__A (.DIODE(_1377_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4497__A (.DIODE(_1377_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4459__A1 (.DIODE(_1377_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4874__A2 (.DIODE(_1378_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4873__B (.DIODE(_1378_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4866__A2 (.DIODE(_1378_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4825__D (.DIODE(_1378_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4788__B (.DIODE(_1378_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4497__B (.DIODE(_1378_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4459__A2 (.DIODE(_1378_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5075__A (.DIODE(_1383_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4839__A2 (.DIODE(_1383_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4464__A (.DIODE(_1383_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5738__A1 (.DIODE(_1384_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5499__A (.DIODE(_1384_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5295__S (.DIODE(_1384_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5243__C1 (.DIODE(_1384_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5112__A (.DIODE(_1384_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5074__A (.DIODE(_1384_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4854__A (.DIODE(_1384_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4818__B (.DIODE(_1384_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4813__S (.DIODE(_1384_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4465__B (.DIODE(_1384_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4532__A3 (.DIODE(_1386_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4526__B (.DIODE(_1386_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4468__A3 (.DIODE(_1386_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4540__A2 (.DIODE(_1388_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4539__C (.DIODE(_1388_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4470__A3 (.DIODE(_1388_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6365__A (.DIODE(_1406_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6361__A (.DIODE(_1406_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4602__C1 (.DIODE(_1406_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4595__C1 (.DIODE(_1406_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4588__C1 (.DIODE(_1406_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4543__S (.DIODE(_1406_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4515__S (.DIODE(_1406_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4505__A (.DIODE(_1406_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4493__A2 (.DIODE(_1406_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4489__A2 (.DIODE(_1406_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5675__B1_N (.DIODE(_1407_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5645__B1_N (.DIODE(_1407_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5609__B1_N (.DIODE(_1407_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5513__B1_N (.DIODE(_1407_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5485__B1_N (.DIODE(_1407_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5448__B1_N (.DIODE(_1407_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5414__B1_N (.DIODE(_1407_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4783__B1_N (.DIODE(_1407_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4605__B (.DIODE(_1407_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4488__B (.DIODE(_1407_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4768__A2 (.DIODE(_1409_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4604__A2 (.DIODE(_1409_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4597__A2 (.DIODE(_1409_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4590__A2 (.DIODE(_1409_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4583__A2 (.DIODE(_1409_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4578__A2 (.DIODE(_1409_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4490__A (.DIODE(_1409_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4572__A2 (.DIODE(_1410_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4566__A2 (.DIODE(_1410_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4559__A2 (.DIODE(_1410_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4553__A2 (.DIODE(_1410_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4545__A2 (.DIODE(_1410_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4538__A2 (.DIODE(_1410_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4531__A2 (.DIODE(_1410_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4525__A2 (.DIODE(_1410_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4517__A2 (.DIODE(_1410_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4510__A2 (.DIODE(_1410_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4582__A2 (.DIODE(_1412_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4577__A2 (.DIODE(_1412_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4571__A2 (.DIODE(_1412_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4564__A2 (.DIODE(_1412_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4558__A2 (.DIODE(_1412_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4552__A2 (.DIODE(_1412_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4537__A2 (.DIODE(_1412_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4530__A2 (.DIODE(_1412_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4524__A2 (.DIODE(_1412_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4507__A2 (.DIODE(_1412_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4767__C1 (.DIODE(_1413_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4603__B1 (.DIODE(_1413_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4596__B1 (.DIODE(_1413_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4589__B1 (.DIODE(_1413_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4544__A (.DIODE(_1413_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4516__A (.DIODE(_1413_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4494__A (.DIODE(_1413_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4582__B1 (.DIODE(_1414_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4577__B1 (.DIODE(_1414_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4571__B1 (.DIODE(_1414_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4564__B1 (.DIODE(_1414_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4558__B1 (.DIODE(_1414_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4552__B1 (.DIODE(_1414_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4537__B1 (.DIODE(_1414_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4530__B1 (.DIODE(_1414_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4524__B1 (.DIODE(_1414_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4507__B1 (.DIODE(_1414_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4601__A (.DIODE(_1415_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4587__A (.DIODE(_1415_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4562__A (.DIODE(_1415_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4550__A (.DIODE(_1415_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4542__S (.DIODE(_1415_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4535__A (.DIODE(_1415_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4522__A (.DIODE(_1415_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4514__S (.DIODE(_1415_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4496__A (.DIODE(_1415_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6362__A1 (.DIODE(_1416_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4913__A (.DIODE(_1416_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4767__A1 (.DIODE(_1416_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4595__A1 (.DIODE(_1416_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4576__A1 (.DIODE(_1416_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4575__A (.DIODE(_1416_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4570__A1 (.DIODE(_1416_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4557__A1 (.DIODE(_1416_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4529__A1 (.DIODE(_1416_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4506__A1 (.DIODE(_1416_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5101__A (.DIODE(_1417_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4865__A1 (.DIODE(_1417_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4824__B (.DIODE(_1417_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4498__A (.DIODE(_1417_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5415__S (.DIODE(_1418_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5124__S (.DIODE(_1418_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5120__S (.DIODE(_1418_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5117__S (.DIODE(_1418_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5105__S (.DIODE(_1418_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5098__A1 (.DIODE(_1418_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5097__A (.DIODE(_1418_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4805__A (.DIODE(_1418_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4803__A (.DIODE(_1418_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4499__A (.DIODE(_1418_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6184__B (.DIODE(_1419_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5685__S (.DIODE(_1419_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5613__S (.DIODE(_1419_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5560__S (.DIODE(_1419_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5493__A1 (.DIODE(_1419_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5452__A (.DIODE(_1419_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5350__S (.DIODE(_1419_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5304__S (.DIODE(_1419_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4849__S (.DIODE(_1419_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4500__B (.DIODE(_1419_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4581__C1 (.DIODE(_1425_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4576__C1 (.DIODE(_1425_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4570__C1 (.DIODE(_1425_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4563__C1 (.DIODE(_1425_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4557__C1 (.DIODE(_1425_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4551__C1 (.DIODE(_1425_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4536__C1 (.DIODE(_1425_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4529__C1 (.DIODE(_1425_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4523__C1 (.DIODE(_1425_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4506__C1 (.DIODE(_1425_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6402__A (.DIODE(_1428_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6397__A (.DIODE(_1428_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6394__A (.DIODE(_1428_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6391__A (.DIODE(_1428_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6385__A (.DIODE(_1428_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6380__A (.DIODE(_1428_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6163__A2 (.DIODE(_1428_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4768__C1 (.DIODE(_1428_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4565__A (.DIODE(_1428_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4509__A (.DIODE(_1428_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6405__B1 (.DIODE(_1429_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6383__B1 (.DIODE(_1429_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4559__C1 (.DIODE(_1429_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4553__C1 (.DIODE(_1429_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4545__C1 (.DIODE(_1429_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4538__C1 (.DIODE(_1429_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4531__C1 (.DIODE(_1429_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4525__C1 (.DIODE(_1429_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4517__C1 (.DIODE(_1429_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4510__C1 (.DIODE(_1429_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6374__A (.DIODE(_1477_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6371__A (.DIODE(_1477_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6368__A (.DIODE(_1477_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4604__C1 (.DIODE(_1477_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4597__C1 (.DIODE(_1477_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4590__C1 (.DIODE(_1477_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4583__C1 (.DIODE(_1477_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4578__C1 (.DIODE(_1477_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4572__C1 (.DIODE(_1477_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4566__C1 (.DIODE(_1477_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4759__B1 (.DIODE(_1512_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4752__A1 (.DIODE(_1512_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4741__B1 (.DIODE(_1512_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4737__B1 (.DIODE(_1512_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4729__B (.DIODE(_1512_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4713__B (.DIODE(_1512_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4711__B (.DIODE(_1512_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4608__A (.DIODE(_1512_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4791__A2 (.DIODE(_1513_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4696__A2 (.DIODE(_1513_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4688__A2 (.DIODE(_1513_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4681__B1 (.DIODE(_1513_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4674__A2 (.DIODE(_1513_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4658__A2 (.DIODE(_1513_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4651__A2 (.DIODE(_1513_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4637__A2 (.DIODE(_1513_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4630__A2 (.DIODE(_1513_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4624__A2 (.DIODE(_1513_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4691__A2 (.DIODE(_1514_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4687__A2 (.DIODE(_1514_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4678__A2 (.DIODE(_1514_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4668__A2 (.DIODE(_1514_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4654__A2 (.DIODE(_1514_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4633__A2 (.DIODE(_1514_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4626__A2 (.DIODE(_1514_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4612__A2 (.DIODE(_1514_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4758__B1 (.DIODE(_1515_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4739__B1 (.DIODE(_1515_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4735__B1 (.DIODE(_1515_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4728__B1 (.DIODE(_1515_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4719__B1 (.DIODE(_1515_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4708__B1 (.DIODE(_1515_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4611__A (.DIODE(_1515_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4748__A2 (.DIODE(_1516_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4694__A2 (.DIODE(_1516_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4687__B1 (.DIODE(_1516_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4678__B1 (.DIODE(_1516_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4672__A2 (.DIODE(_1516_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4654__B1 (.DIODE(_1516_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4646__B1 (.DIODE(_1516_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4635__B1 (.DIODE(_1516_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4626__B1 (.DIODE(_1516_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4612__B1 (.DIODE(_1516_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4757__A2 (.DIODE(_1518_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4740__A2 (.DIODE(_1518_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4727__A2 (.DIODE(_1518_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4719__A2 (.DIODE(_1518_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4708__A2 (.DIODE(_1518_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4614__A (.DIODE(_1518_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4747__A2 (.DIODE(_1519_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4735__A2 (.DIODE(_1519_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4693__A3 (.DIODE(_1519_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4680__A3 (.DIODE(_1519_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4670__A (.DIODE(_1519_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4653__C (.DIODE(_1519_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4649__A2 (.DIODE(_1519_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4635__A3 (.DIODE(_1519_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4628__A3 (.DIODE(_1519_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4616__A3 (.DIODE(_1519_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4693__B1 (.DIODE(_1522_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4686__A2 (.DIODE(_1522_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4676__B1 (.DIODE(_1522_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4668__B1 (.DIODE(_1522_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4657__B1 (.DIODE(_1522_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4632__A2 (.DIODE(_1522_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4625__B (.DIODE(_1522_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4622__A2 (.DIODE(_1522_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4695__A2 (.DIODE(_1523_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4684__A2 (.DIODE(_1523_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4676__A2 (.DIODE(_1523_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4673__A2 (.DIODE(_1523_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4657__A2 (.DIODE(_1523_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4636__A2 (.DIODE(_1523_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4629__A2 (.DIODE(_1523_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4621__A2 (.DIODE(_1523_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4758__A2 (.DIODE(_1524_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4739__A2 (.DIODE(_1524_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4736__A2 (.DIODE(_1524_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4728__A2 (.DIODE(_1524_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4714__A2 (.DIODE(_1524_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4709__A2 (.DIODE(_1524_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4620__A (.DIODE(_1524_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4747__B1 (.DIODE(_1525_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4691__B1 (.DIODE(_1525_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4683__B1 (.DIODE(_1525_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4677__A2 (.DIODE(_1525_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4673__B1 (.DIODE(_1525_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4656__A2 (.DIODE(_1525_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4646__A2 (.DIODE(_1525_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4632__B1 (.DIODE(_1525_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4629__B1 (.DIODE(_1525_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4621__B1 (.DIODE(_1525_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6533__S (.DIODE(_1529_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6357__B1 (.DIODE(_1529_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6352__A3 (.DIODE(_1529_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5749__A1 (.DIODE(_1529_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5736__A2 (.DIODE(_1529_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5498__A (.DIODE(_1529_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5224__A1 (.DIODE(_1529_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4979__B (.DIODE(_1529_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4842__B (.DIODE(_1529_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4769__A2 (.DIODE(_1529_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6303__A0 (.DIODE(_1535_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6285__B1 (.DIODE(_1535_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6277__A3 (.DIODE(_1535_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5554__B1 (.DIODE(_1535_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5220__A1_N (.DIODE(_1535_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5115__A2 (.DIODE(_1535_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5005__B (.DIODE(_1535_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5004__B (.DIODE(_1535_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4631__A (.DIODE(_1535_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5055__B (.DIODE(_1536_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5054__A2 (.DIODE(_1536_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4811__B2 (.DIODE(_1536_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4640__A2 (.DIODE(_1536_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5051__B (.DIODE(_1542_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4638__A (.DIODE(_1542_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6304__A0 (.DIODE(_1543_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6298__A1 (.DIODE(_1543_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5591__B1 (.DIODE(_1543_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5222__A1_N (.DIODE(_1543_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5116__A2 (.DIODE(_1543_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5052__B (.DIODE(_1543_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5001__B (.DIODE(_1543_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5000__A2 (.DIODE(_1543_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4811__A1_N (.DIODE(_1543_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4639__B (.DIODE(_1543_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4755__A2 (.DIODE(_1547_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4750__A2 (.DIODE(_1547_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4743__A2 (.DIODE(_1547_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4734__A2 (.DIODE(_1547_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4645__A2 (.DIODE(_1547_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4755__B1 (.DIODE(_1548_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4750__B1 (.DIODE(_1548_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4743__B1 (.DIODE(_1548_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4734__B1 (.DIODE(_1548_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4645__B1 (.DIODE(_1548_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4757__B1 (.DIODE(_1552_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4748__B1 (.DIODE(_1552_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4740__B1 (.DIODE(_1552_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4736__B1 (.DIODE(_1552_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4714__B1 (.DIODE(_1552_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4709__B1 (.DIODE(_1552_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4649__B1 (.DIODE(_1552_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4820__A2 (.DIODE(_1553_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4819__A2 (.DIODE(_1553_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4757__C1 (.DIODE(_1553_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4751__A2 (.DIODE(_1553_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4745__A2 (.DIODE(_1553_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4738__A2 (.DIODE(_1553_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4719__C1 (.DIODE(_1553_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4708__C1 (.DIODE(_1553_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4649__C1 (.DIODE(_1553_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5085__B (.DIODE(_1556_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5047__B (.DIODE(_1556_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5011__B (.DIODE(_1556_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5010__B (.DIODE(_1556_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4652__A (.DIODE(_1556_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6277__A1 (.DIODE(_1557_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6262__B1 (.DIODE(_1557_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6254__A2 (.DIODE(_1557_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5518__B (.DIODE(_1557_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5502__B1 (.DIODE(_1557_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5239__A1_N (.DIODE(_1557_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5100__B (.DIODE(_1557_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5046__A2 (.DIODE(_1557_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4816__B2 (.DIODE(_1557_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4662__A0 (.DIODE(_1557_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5044__B (.DIODE(_1563_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4659__A (.DIODE(_1563_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6303__A1 (.DIODE(_1564_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6277__A2 (.DIODE(_1564_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6274__B1 (.DIODE(_1564_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5519__B1 (.DIODE(_1564_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5517__C (.DIODE(_1564_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5099__A2 (.DIODE(_1564_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5043__B (.DIODE(_1564_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5003__A (.DIODE(_1564_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4816__A1 (.DIODE(_1564_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4662__A1 (.DIODE(_1564_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6226__A1 (.DIODE(_1569_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6225__A (.DIODE(_1569_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6205__A1_N (.DIODE(_1569_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6203__C (.DIODE(_1569_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6196__A1 (.DIODE(_1569_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4703__A (.DIODE(_1569_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4666__A (.DIODE(_1569_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6301__A1 (.DIODE(_1570_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6290__A1 (.DIODE(_1570_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6289__A (.DIODE(_1570_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6224__A1 (.DIODE(_1570_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6214__A2 (.DIODE(_1570_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6204__A2 (.DIODE(_1570_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6189__A (.DIODE(_1570_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4908__A (.DIODE(_1570_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4702__B (.DIODE(_1570_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4666__B (.DIODE(_1570_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5185__A2 (.DIODE(_1575_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5179__A2 (.DIODE(_1575_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5174__A2 (.DIODE(_1575_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5167__A2 (.DIODE(_1575_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5163__A2 (.DIODE(_1575_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5154__A2 (.DIODE(_1575_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5142__B (.DIODE(_1575_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4977__A2 (.DIODE(_1575_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4683__A3 (.DIODE(_1575_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4671__C (.DIODE(_1575_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5059__B (.DIODE(_1579_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4675__A (.DIODE(_1579_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6328__A0 (.DIODE(_1580_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6323__B1 (.DIODE(_1580_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5653__A1 (.DIODE(_1580_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5223__B2 (.DIODE(_1580_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5119__A2 (.DIODE(_1580_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5060__B (.DIODE(_1580_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4993__B (.DIODE(_1580_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4992__A2 (.DIODE(_1580_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4810__A1 (.DIODE(_1580_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4682__A0 (.DIODE(_1580_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6304__A1 (.DIODE(_1586_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5618__B1 (.DIODE(_1586_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5221__B (.DIODE(_1586_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5118__A2 (.DIODE(_1586_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5063__A2 (.DIODE(_1586_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5062__A (.DIODE(_1586_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4998__B (.DIODE(_1586_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4996__B (.DIODE(_1586_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4810__B2 (.DIODE(_1586_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4682__A1 (.DIODE(_1586_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5123__A2 (.DIODE(_1593_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4689__A (.DIODE(_1593_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6351__A2 (.DIODE(_1594_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6346__A1 (.DIODE(_1594_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5715__A1 (.DIODE(_1594_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5224__B2 (.DIODE(_1594_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5069__B (.DIODE(_1594_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4985__B (.DIODE(_1594_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4984__B (.DIODE(_1594_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4982__A2 (.DIODE(_1594_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4806__A1_N (.DIODE(_1594_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4701__B1 (.DIODE(_1594_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6396__A2 (.DIODE(_1595_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6373__A2 (.DIODE(_1595_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4906__B (.DIODE(_1595_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4701__B2 (.DIODE(_1595_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4990__B (.DIODE(_1601_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4988__B (.DIODE(_1601_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4983__A (.DIODE(_1601_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4806__B2 (.DIODE(_1601_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4700__A (.DIODE(_1601_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6364__B (.DIODE(_1603_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6329__A (.DIODE(_1603_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6305__S (.DIODE(_1603_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6278__A2 (.DIODE(_1603_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6277__S1 (.DIODE(_1603_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6265__S (.DIODE(_1603_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6234__A (.DIODE(_1603_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6196__A3 (.DIODE(_1603_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4905__B (.DIODE(_1603_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4699__B (.DIODE(_1603_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6366__A (.DIODE(_1608_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6352__A1 (.DIODE(_1608_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6327__A (.DIODE(_1608_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6278__B1 (.DIODE(_1608_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6257__A1 (.DIODE(_1608_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6256__A (.DIODE(_1608_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6197__A1 (.DIODE(_1608_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6190__A1 (.DIODE(_1608_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6179__A1 (.DIODE(_1608_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4765__A (.DIODE(_1608_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4823__A (.DIODE(_1615_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4712__A1 (.DIODE(_1615_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6194__A2 (.DIODE(_1618_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4847__A (.DIODE(_1618_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4827__A (.DIODE(_1618_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4721__A1 (.DIODE(_1618_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6194__A3 (.DIODE(_1625_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4847__B (.DIODE(_1625_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4827__B (.DIODE(_1625_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4721__A2 (.DIODE(_1625_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6193__A2 (.DIODE(_1632_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4837__A2 (.DIODE(_1632_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4730__A2 (.DIODE(_1632_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6193__A3 (.DIODE(_1633_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4837__A3 (.DIODE(_1633_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4730__A3 (.DIODE(_1633_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6222__B (.DIODE(_1635_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6212__A1 (.DIODE(_1635_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6188__C (.DIODE(_1635_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4874__B1 (.DIODE(_1635_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4873__C (.DIODE(_1635_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4732__B1 (.DIODE(_1635_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6289__B (.DIODE(_1637_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6204__A3 (.DIODE(_1637_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6203__B_N (.DIODE(_1637_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4764__A0 (.DIODE(_1637_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5163__B1 (.DIODE(_1639_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4819__B1 (.DIODE(_1639_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4738__B1 (.DIODE(_1639_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4819__C1 (.DIODE(_1642_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4738__C1 (.DIODE(_1642_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6221__A2 (.DIODE(_1643_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6212__A2 (.DIODE(_1643_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5344__A1 (.DIODE(_1643_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5106__B (.DIODE(_1643_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5035__B (.DIODE(_1643_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5031__B (.DIODE(_1643_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5030__B (.DIODE(_1643_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4746__A0 (.DIODE(_1643_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4820__B1 (.DIODE(_1646_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4745__B1 (.DIODE(_1646_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5167__B1 (.DIODE(_1648_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4744__B (.DIODE(_1648_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6221__A3 (.DIODE(_1650_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5380__A2 (.DIODE(_1650_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5238__B2 (.DIODE(_1650_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5082__B (.DIODE(_1650_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5034__B (.DIODE(_1650_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4746__A1 (.DIODE(_1650_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4752__A2 (.DIODE(_1653_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5018__B (.DIODE(_1657_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4753__A (.DIODE(_1657_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6277__A0 (.DIODE(_1658_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6254__A0 (.DIODE(_1658_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6249__A1 (.DIODE(_1658_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5462__B1 (.DIODE(_1658_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5094__B (.DIODE(_1658_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5017__B (.DIODE(_1658_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5014__A (.DIODE(_1658_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5013__A2 (.DIODE(_1658_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4814__A1 (.DIODE(_1658_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4761__A0 (.DIODE(_1658_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5083__B (.DIODE(_1664_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5081__B (.DIODE(_1664_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5023__B (.DIODE(_1664_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4760__A (.DIODE(_1664_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6254__A3 (.DIODE(_1665_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6243__B2 (.DIODE(_1665_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6235__A3 (.DIODE(_1665_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5429__B1 (.DIODE(_1665_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5238__A1_N (.DIODE(_1665_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5096__A2 (.DIODE(_1665_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5021__A2 (.DIODE(_1665_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5020__A (.DIODE(_1665_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4814__B2 (.DIODE(_1665_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4761__A1 (.DIODE(_1665_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6244__B (.DIODE(_1669_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4765__B (.DIODE(_1669_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6342__B (.DIODE(_1671_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6341__B (.DIODE(_1671_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4767__B1 (.DIODE(_1671_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6504__A (.DIODE(_1679_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6471__B1 (.DIODE(_1679_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6464__A (.DIODE(_1679_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6458__B1 (.DIODE(_1679_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6454__B1 (.DIODE(_1679_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6436__B1 (.DIODE(_1679_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6435__C1 (.DIODE(_1679_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6428__B1 (.DIODE(_1679_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6421__A (.DIODE(_1679_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4779__A2 (.DIODE(_1679_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6701__A3 (.DIODE(_1681_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6497__B (.DIODE(_1681_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6491__A (.DIODE(_1681_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6442__A1 (.DIODE(_1681_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6420__A (.DIODE(_1681_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6418__A3 (.DIODE(_1681_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6413__B (.DIODE(_1681_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4778__C (.DIODE(_1681_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5752__A2 (.DIODE(_1685_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5721__A2 (.DIODE(_1685_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5582__A2 (.DIODE(_1685_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5548__A2 (.DIODE(_1685_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5387__A2 (.DIODE(_1685_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5365__A2 (.DIODE(_1685_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5292__A2 (.DIODE(_1685_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4782__A (.DIODE(_1685_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5675__A2 (.DIODE(_1686_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5645__A2 (.DIODE(_1686_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5609__A2 (.DIODE(_1686_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5513__A2 (.DIODE(_1686_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5485__A2 (.DIODE(_1686_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5448__A2 (.DIODE(_1686_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5414__A2 (.DIODE(_1686_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5336__A2 (.DIODE(_1686_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5252__A1 (.DIODE(_1686_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4783__A2 (.DIODE(_1686_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6174__A2 (.DIODE(_1689_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5617__A (.DIODE(_1689_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5500__B2 (.DIODE(_1689_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5425__B1 (.DIODE(_1689_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5339__A2 (.DIODE(_1689_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5300__A1 (.DIODE(_1689_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5035__A (.DIODE(_1689_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4834__A1 (.DIODE(_1689_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4830__A (.DIODE(_1689_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4818__A (.DIODE(_1689_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5370__S (.DIODE(_1691_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5353__S (.DIODE(_1691_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5346__A1 (.DIODE(_1691_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5345__S (.DIODE(_1691_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5294__S (.DIODE(_1691_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5293__S (.DIODE(_1691_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5243__A1 (.DIODE(_1691_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4822__A (.DIODE(_1691_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4812__S (.DIODE(_1691_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4790__A (.DIODE(_1691_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5492__A (.DIODE(_1692_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5416__S (.DIODE(_1692_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5221__A (.DIODE(_1692_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5126__A1 (.DIODE(_1692_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5110__A1 (.DIODE(_1692_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5109__A (.DIODE(_1692_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5102__A1 (.DIODE(_1692_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4835__A2 (.DIODE(_1692_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4809__A (.DIODE(_1692_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4789__A (.DIODE(_1692_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6175__A2 (.DIODE(_1693_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5741__A1 (.DIODE(_1693_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5740__A (.DIODE(_1693_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5586__A1 (.DIODE(_1693_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5453__A1 (.DIODE(_1693_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5367__S (.DIODE(_1693_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5242__A1 (.DIODE(_1693_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5235__A2 (.DIODE(_1693_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4821__S (.DIODE(_1693_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4790__B (.DIODE(_1693_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5584__A1_N (.DIODE(_1694_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5306__A1 (.DIODE(_1694_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4807__A1_N (.DIODE(_1694_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5125__A (.DIODE(_1695_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5091__B (.DIODE(_1695_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5070__A2 (.DIODE(_1695_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4980__B (.DIODE(_1695_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4800__A (.DIODE(_1695_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6170__B2 (.DIODE(_1696_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5429__A2 (.DIODE(_1696_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5093__A (.DIODE(_1696_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5083__A (.DIODE(_1696_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5081__A (.DIODE(_1696_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5022__A1 (.DIODE(_1696_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4804__A (.DIODE(_1696_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4799__A (.DIODE(_1696_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6169__B2 (.DIODE(_1699_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5680__A2 (.DIODE(_1699_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4798__A (.DIODE(_1699_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4841__B (.DIODE(_1702_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4804__C (.DIODE(_1702_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4799__C (.DIODE(_1702_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5242__B1 (.DIODE(_1703_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5222__B2 (.DIODE(_1703_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4829__A (.DIODE(_1703_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4809__B (.DIODE(_1703_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4803__B (.DIODE(_1703_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4800__B (.DIODE(_1703_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5242__D1 (.DIODE(_1705_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5240__S (.DIODE(_1705_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4886__A2 (.DIODE(_1705_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4870__A (.DIODE(_1705_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4824__A (.DIODE(_1705_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4802__A (.DIODE(_1705_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6175__B2 (.DIODE(_1706_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5372__S (.DIODE(_1706_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5347__A1 (.DIODE(_1706_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5298__A (.DIODE(_1706_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5297__S (.DIODE(_1706_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5226__S0 (.DIODE(_1706_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4869__A (.DIODE(_1706_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4868__A (.DIODE(_1706_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4817__S (.DIODE(_1706_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4807__B1 (.DIODE(_1706_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6235__A1 (.DIODE(_1723_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6218__B1 (.DIODE(_1723_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5241__A1_N (.DIODE(_1723_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4821__A0 (.DIODE(_1723_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6254__A1 (.DIODE(_1724_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6235__A2 (.DIODE(_1724_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6231__A1 (.DIODE(_1724_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5381__B1 (.DIODE(_1724_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5108__A2 (.DIODE(_1724_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5025__B (.DIODE(_1724_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5024__A2 (.DIODE(_1724_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4821__A1 (.DIODE(_1724_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6221__A1 (.DIODE(_1727_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6212__A3 (.DIODE(_1727_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5315__A (.DIODE(_1727_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5241__B2 (.DIODE(_1727_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5103__A (.DIODE(_1727_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5075__B (.DIODE(_1727_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5074__B (.DIODE(_1727_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5029__B (.DIODE(_1727_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5027__B (.DIODE(_1727_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4828__A1 (.DIODE(_1727_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5498__C (.DIODE(_1730_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5369__A2 (.DIODE(_1730_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5355__A3 (.DIODE(_1730_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4859__B (.DIODE(_1730_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4854__B (.DIODE(_1730_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4851__B (.DIODE(_1730_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4839__A3 (.DIODE(_1730_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4828__B1 (.DIODE(_1730_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6221__A0 (.DIODE(_1731_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6212__A0 (.DIODE(_1731_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5242__A2 (.DIODE(_1731_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4885__A (.DIODE(_1731_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4878__B (.DIODE(_1731_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4871__B (.DIODE(_1731_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4828__B2 (.DIODE(_1731_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5617__B (.DIODE(_1736_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5500__C1 (.DIODE(_1736_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5356__B (.DIODE(_1736_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5300__B1 (.DIODE(_1736_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5248__A2 (.DIODE(_1736_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4833__C1 (.DIODE(_1736_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5741__C1 (.DIODE(_1740_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5586__C1 (.DIODE(_1740_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5584__B2 (.DIODE(_1740_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5368__S (.DIODE(_1740_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5127__A1 (.DIODE(_1740_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5126__B1 (.DIODE(_1740_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4850__A (.DIODE(_1740_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6192__B2 (.DIODE(_1741_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6190__A3 (.DIODE(_1741_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5301__A2 (.DIODE(_1741_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5235__B1 (.DIODE(_1741_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4864__A (.DIODE(_1741_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4863__A (.DIODE(_1741_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4845__A2 (.DIODE(_1741_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5106__A (.DIODE(_1742_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4859__A (.DIODE(_1742_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4842__A (.DIODE(_1742_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4840__A (.DIODE(_1742_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4839__C1 (.DIODE(_1742_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5119__B1 (.DIODE(_1747_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5118__B1 (.DIODE(_1747_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5116__B1 (.DIODE(_1747_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5115__B1 (.DIODE(_1747_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5108__B1 (.DIODE(_1747_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5104__B1 (.DIODE(_1747_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5099__B1 (.DIODE(_1747_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5096__B1 (.DIODE(_1747_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4848__B1 (.DIODE(_1747_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4844__A (.DIODE(_1747_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5123__A1 (.DIODE(_1750_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5122__A1 (.DIODE(_1750_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5119__A1 (.DIODE(_1750_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5118__A1 (.DIODE(_1750_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5116__A1 (.DIODE(_1750_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5115__A1 (.DIODE(_1750_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5104__A1 (.DIODE(_1750_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5099__A1 (.DIODE(_1750_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4855__A (.DIODE(_1750_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4848__A1 (.DIODE(_1750_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6201__B2 (.DIODE(_1751_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5302__A2 (.DIODE(_1751_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4870__B (.DIODE(_1751_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4866__C1 (.DIODE(_1751_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4865__C1 (.DIODE(_1751_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4848__A2 (.DIODE(_1751_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5744__A1 (.DIODE(_1757_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5658__C1 (.DIODE(_1757_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5621__A1 (.DIODE(_1757_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5595__A1 (.DIODE(_1757_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5565__B1_N (.DIODE(_1757_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5516__A (.DIODE(_1757_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5227__A (.DIODE(_1757_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4858__A (.DIODE(_1757_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5716__B2 (.DIODE(_1762_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5688__C1 (.DIODE(_1762_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5466__A1 (.DIODE(_1762_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5432__A1 (.DIODE(_1762_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5384__A1 (.DIODE(_1762_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5318__A1 (.DIODE(_1762_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4889__A2 (.DIODE(_1762_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5230__B1 (.DIODE(_1766_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5229__A (.DIODE(_1766_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4875__A1 (.DIODE(_1766_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4864__B (.DIODE(_1766_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4863__B (.DIODE(_1766_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5718__A1 (.DIODE(_1785_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5650__A (.DIODE(_1785_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5550__B1 (.DIODE(_1785_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5526__A1 (.DIODE(_1785_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5487__B1 (.DIODE(_1785_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5376__A (.DIODE(_1785_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5338__A (.DIODE(_1785_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5308__A1_N (.DIODE(_1785_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5230__A1 (.DIODE(_1785_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4883__C (.DIODE(_1785_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5749__A2 (.DIODE(_1787_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5715__A2 (.DIODE(_1787_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5680__B2 (.DIODE(_1787_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5653__A2 (.DIODE(_1787_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5618__B2 (.DIODE(_1787_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5591__B2 (.DIODE(_1787_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5554__B2 (.DIODE(_1787_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5519__B2 (.DIODE(_1787_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4884__B (.DIODE(_1787_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4890__B (.DIODE(_1793_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5760__A1 (.DIODE(_1797_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5277__A1 (.DIODE(_1797_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4899__A2 (.DIODE(_1797_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5483__A1 (.DIODE(_1798_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5446__S (.DIODE(_1798_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5410__A1 (.DIODE(_1798_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5396__S (.DIODE(_1798_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5334__S (.DIODE(_1798_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5290__A2 (.DIODE(_1798_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5272__B1 (.DIODE(_1798_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5191__B (.DIODE(_1798_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4895__A (.DIODE(_1798_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6410__A (.DIODE(_1799_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5732__S (.DIODE(_1799_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5703__A1 (.DIODE(_1799_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5673__A1 (.DIODE(_1799_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5643__A1 (.DIODE(_1799_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5633__S (.DIODE(_1799_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5580__A1 (.DIODE(_1799_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5546__A1 (.DIODE(_1799_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5534__S (.DIODE(_1799_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4896__A (.DIODE(_1799_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6505__B2 (.DIODE(_1801_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6487__A2 (.DIODE(_1801_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6479__B2 (.DIODE(_1801_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6472__A2 (.DIODE(_1801_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6459__B2 (.DIODE(_1801_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6451__A2 (.DIODE(_1801_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6435__B2 (.DIODE(_1801_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6430__B2 (.DIODE(_1801_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6423__B2 (.DIODE(_1801_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4899__B1 (.DIODE(_1801_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4903__A (.DIODE(_1805_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6396__A1 (.DIODE(_1810_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6393__A1 (.DIODE(_1810_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6390__A1 (.DIODE(_1810_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6376__A (.DIODE(_1810_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6373__A1 (.DIODE(_1810_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6370__A1 (.DIODE(_1810_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6367__A1 (.DIODE(_1810_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6178__B1 (.DIODE(_1810_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4911__A1 (.DIODE(_1810_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4909__A (.DIODE(_1810_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4955__B (.DIODE(_1818_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4953__B (.DIODE(_1818_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4951__B (.DIODE(_1818_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4949__B (.DIODE(_1818_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4947__B (.DIODE(_1818_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4945__B (.DIODE(_1818_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4936__B (.DIODE(_1818_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4927__B (.DIODE(_1818_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4925__B (.DIODE(_1818_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4923__B (.DIODE(_1818_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4955__C (.DIODE(_1819_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4953__C (.DIODE(_1819_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4951__C (.DIODE(_1819_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4949__C (.DIODE(_1819_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4947__C (.DIODE(_1819_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4945__C (.DIODE(_1819_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4936__C (.DIODE(_1819_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4927__C (.DIODE(_1819_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4925__C (.DIODE(_1819_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4923__C (.DIODE(_1819_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4955__D (.DIODE(_1820_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4953__D (.DIODE(_1820_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4951__D (.DIODE(_1820_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4949__D (.DIODE(_1820_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4947__D (.DIODE(_1820_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4945__D (.DIODE(_1820_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4936__D (.DIODE(_1820_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4927__D (.DIODE(_1820_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4925__D (.DIODE(_1820_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4923__D (.DIODE(_1820_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4926__B1 (.DIODE(_1822_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4960__A2 (.DIODE(_1825_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4958__A2 (.DIODE(_1825_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4956__A2 (.DIODE(_1825_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4954__A2 (.DIODE(_1825_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4952__A2 (.DIODE(_1825_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4950__A2 (.DIODE(_1825_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4942__B (.DIODE(_1825_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4939__B (.DIODE(_1825_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4934__A2 (.DIODE(_1825_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4931__B (.DIODE(_1825_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5823__C1 (.DIODE(_1834_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4960__C1 (.DIODE(_1834_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4958__C1 (.DIODE(_1834_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4956__C1 (.DIODE(_1834_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4954__C1 (.DIODE(_1834_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4952__C1 (.DIODE(_1834_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4950__C1 (.DIODE(_1834_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4948__C1 (.DIODE(_1834_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4946__C1 (.DIODE(_1834_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4944__C1 (.DIODE(_1834_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5809__S (.DIODE(_1845_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5807__S (.DIODE(_1845_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5805__S (.DIODE(_1845_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5803__S (.DIODE(_1845_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5801__S (.DIODE(_1845_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4974__A (.DIODE(_1845_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5812__A2 (.DIODE(_1846_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5799__S (.DIODE(_1846_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5797__S (.DIODE(_1846_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5795__S (.DIODE(_1846_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5793__S (.DIODE(_1846_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5791__S (.DIODE(_1846_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5667__A2 (.DIODE(_1846_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5637__B1 (.DIODE(_1846_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5189__B (.DIODE(_1846_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4975__S (.DIODE(_1846_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5737__B2 (.DIODE(_1849_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5141__A1 (.DIODE(_1849_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5135__A (.DIODE(_1849_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5070__A1 (.DIODE(_1849_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4979__A (.DIODE(_1849_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6532__A2 (.DIODE(_1852_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6531__B (.DIODE(_1852_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5746__A1 (.DIODE(_1852_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5745__B1 (.DIODE(_1852_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5738__B1 (.DIODE(_1852_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5069__C (.DIODE(_1852_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4982__B1 (.DIODE(_1852_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6338__B1 (.DIODE(_1854_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6328__A1 (.DIODE(_1854_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5680__B1 (.DIODE(_1854_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5223__A1 (.DIODE(_1854_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5122__A2 (.DIODE(_1854_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5067__A2 (.DIODE(_1854_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4987__B (.DIODE(_1854_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6176__A2 (.DIODE(_1866_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5618__A2 (.DIODE(_1866_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5064__A1 (.DIODE(_1866_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4998__A (.DIODE(_1866_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4996__A (.DIODE(_1866_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5521__A2 (.DIODE(_1916_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5514__B (.DIODE(_1916_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5087__B1 (.DIODE(_1916_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5047__C (.DIODE(_1916_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5046__B1 (.DIODE(_1916_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5654__A2 (.DIODE(_1932_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5649__A (.DIODE(_1932_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5089__C1 (.DIODE(_1932_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5063__B1 (.DIODE(_1932_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5062__B (.DIODE(_1932_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6235__A0 (.DIODE(_1974_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6208__A1 (.DIODE(_1974_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5303__A2 (.DIODE(_1974_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5104__A2 (.DIODE(_1974_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5709__S (.DIODE(_1982_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5494__S (.DIODE(_1982_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5417__S (.DIODE(_1982_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5305__A (.DIODE(_1982_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5121__S (.DIODE(_1982_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5113__S0 (.DIODE(_1982_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5134__C1 (.DIODE(_2004_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5811__C (.DIODE(_2009_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5638__A2 (.DIODE(_2009_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5190__A1 (.DIODE(_2009_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5183__S (.DIODE(_2009_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5177__S (.DIODE(_2009_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5172__S (.DIODE(_2009_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5165__S (.DIODE(_2009_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5160__A2 (.DIODE(_2009_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5148__S (.DIODE(_2009_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5139__S (.DIODE(_2009_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5169__C (.DIODE(_2024_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5162__A3 (.DIODE(_2024_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5161__B (.DIODE(_2024_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5159__A2 (.DIODE(_2024_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5156__B (.DIODE(_2024_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5169__D_N (.DIODE(_2030_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5168__B (.DIODE(_2030_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5164__B (.DIODE(_2030_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5180__B (.DIODE(_2039_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5176__A (.DIODE(_2039_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5188__B1 (.DIODE(_2048_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5187__C (.DIODE(_2048_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5445__B2 (.DIODE(_2054_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5408__B2 (.DIODE(_2054_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5395__B2 (.DIODE(_2054_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5333__B2 (.DIODE(_2054_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5289__B1 (.DIODE(_2054_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5274__A (.DIODE(_2054_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5271__B1 (.DIODE(_2054_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5193__B (.DIODE(_2054_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5477__A (.DIODE(_2057_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5442__A2 (.DIODE(_2057_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5406__A2 (.DIODE(_2057_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5390__A2 (.DIODE(_2057_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5330__B1 (.DIODE(_2057_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5283__A2 (.DIODE(_2057_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5267__A2 (.DIODE(_2057_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5201__A2 (.DIODE(_2057_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5480__B1 (.DIODE(_2065_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5442__B1 (.DIODE(_2065_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5407__B1 (.DIODE(_2065_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5390__B1 (.DIODE(_2065_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5329__B1 (.DIODE(_2065_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5265__A2 (.DIODE(_2065_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5208__A2 (.DIODE(_2065_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5441__A (.DIODE(_2071_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5405__B1 (.DIODE(_2071_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5391__B1 (.DIODE(_2071_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5328__B1 (.DIODE(_2071_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5284__B1 (.DIODE(_2071_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5265__B1 (.DIODE(_2071_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5213__A2 (.DIODE(_2071_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5751__A1 (.DIODE(_2081_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5720__A1 (.DIODE(_2081_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5601__A1 (.DIODE(_2081_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5507__A1 (.DIODE(_2081_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5469__A1 (.DIODE(_2081_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5434__A1 (.DIODE(_2081_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5386__A1 (.DIODE(_2081_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5251__A1 (.DIODE(_2081_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6174__B1 (.DIODE(_2087_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5459__A (.DIODE(_2087_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5425__A1 (.DIODE(_2087_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5371__A (.DIODE(_2087_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5369__A1 (.DIODE(_2087_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5348__A1 (.DIODE(_2087_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5346__B1 (.DIODE(_2087_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5316__A2 (.DIODE(_2087_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5299__S (.DIODE(_2087_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5226__S1 (.DIODE(_2087_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5502__B2 (.DIODE(_2094_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5462__B2 (.DIODE(_2094_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5429__B2 (.DIODE(_2094_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5381__B2 (.DIODE(_2094_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5235__B2 (.DIODE(_2094_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5593__A1 (.DIODE(_2095_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5380__B1 (.DIODE(_2095_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5234__A (.DIODE(_2095_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5594__A1 (.DIODE(_2107_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5557__B (.DIODE(_2107_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5522__B2 (.DIODE(_2107_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5348__C1 (.DIODE(_2107_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5246__C1 (.DIODE(_2107_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6541__B (.DIODE(_2110_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6515__B (.DIODE(_2110_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5251__A2 (.DIODE(_2110_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5252__B2 (.DIODE(_2113_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6412__B1 (.DIODE(_2114_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5758__A1 (.DIODE(_2114_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5256__A1 (.DIODE(_2114_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5399__B1_N (.DIODE(_2115_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5254__A (.DIODE(_2115_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5754__S (.DIODE(_2116_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5724__S (.DIODE(_2116_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5694__S (.DIODE(_2116_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5603__S (.DIODE(_2116_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5571__S (.DIODE(_2116_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5536__B1 (.DIODE(_2116_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5509__S (.DIODE(_2116_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5400__A1 (.DIODE(_2116_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5275__B1_N (.DIODE(_2116_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5255__A (.DIODE(_2116_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5664__S (.DIODE(_2117_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5636__A1 (.DIODE(_2117_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5635__B1_N (.DIODE(_2117_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5537__A1 (.DIODE(_2117_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5471__S (.DIODE(_2117_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5436__S (.DIODE(_2117_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5361__S (.DIODE(_2117_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5323__S (.DIODE(_2117_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5277__A2 (.DIODE(_2117_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5256__S (.DIODE(_2117_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5573__S (.DIODE(_2120_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5539__S (.DIODE(_2120_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5511__S (.DIODE(_2120_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5473__S (.DIODE(_2120_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5438__S (.DIODE(_2120_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5403__S (.DIODE(_2120_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5363__S (.DIODE(_2120_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5325__S (.DIODE(_2120_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5279__S (.DIODE(_2120_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5259__S (.DIODE(_2120_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5440__A (.DIODE(_2122_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5408__A2 (.DIODE(_2122_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5395__A2 (.DIODE(_2122_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5333__A2 (.DIODE(_2122_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5281__A2 (.DIODE(_2122_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5262__B (.DIODE(_2122_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6707__B (.DIODE(_2129_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5478__A2 (.DIODE(_2129_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5444__B1 (.DIODE(_2129_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5405__A2 (.DIODE(_2129_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5393__B1 (.DIODE(_2129_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5331__B1 (.DIODE(_2129_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5284__A2 (.DIODE(_2129_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5270__B1 (.DIODE(_2129_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5272__A2 (.DIODE(_2132_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5731__B2 (.DIODE(_2135_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5701__B2 (.DIODE(_2135_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5671__B2 (.DIODE(_2135_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5641__B2 (.DIODE(_2135_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5632__B2 (.DIODE(_2135_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5578__B2 (.DIODE(_2135_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5544__B2 (.DIODE(_2135_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5533__B2 (.DIODE(_2135_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5481__B2 (.DIODE(_2135_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5276__A1 (.DIODE(_2135_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5476__A (.DIODE(_2146_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5443__A2 (.DIODE(_2146_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5406__B1 (.DIODE(_2146_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5391__A2 (.DIODE(_2146_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5329__A2 (.DIODE(_2146_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5288__B1 (.DIODE(_2146_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5742__A1 (.DIODE(_2165_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5686__S (.DIODE(_2165_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5656__S0 (.DIODE(_2165_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5614__S (.DIODE(_2165_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5587__A1 (.DIODE(_2165_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5562__A1 (.DIODE(_2165_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5561__A (.DIODE(_2165_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5454__S (.DIODE(_2165_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5351__S (.DIODE(_2165_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5306__B2 (.DIODE(_2165_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5748__A1 (.DIODE(_2172_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5708__B1 (.DIODE(_2172_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5646__B1 (.DIODE(_2172_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5524__B1 (.DIODE(_2172_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5491__A (.DIODE(_2172_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5451__B (.DIODE(_2172_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5423__B1 (.DIODE(_2172_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5379__A (.DIODE(_2172_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5344__B2 (.DIODE(_2172_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5313__B2 (.DIODE(_2172_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5319__B1 (.DIODE(_2178_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5322__B2 (.DIODE(_2181_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6424__A2 (.DIODE(_2182_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5762__A1 (.DIODE(_2182_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5323__A1 (.DIODE(_2182_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5620__A2 (.DIODE(_2214_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5356__C_N (.DIODE(_2214_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6539__B (.DIODE(_2216_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6516__D_N (.DIODE(_2216_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5358__B (.DIODE(_2216_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6431__A2 (.DIODE(_2219_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5764__A1 (.DIODE(_2219_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5361__A1 (.DIODE(_2219_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5654__B2 (.DIODE(_2229_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5374__A2 (.DIODE(_2229_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6540__A (.DIODE(_2242_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6514__A (.DIODE(_2242_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5386__A2 (.DIODE(_2242_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5387__B2 (.DIODE(_2244_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6434__B (.DIODE(_2245_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5388__A (.DIODE(_2245_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5729__C1 (.DIODE(_2247_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5699__C1 (.DIODE(_2247_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5669__C1 (.DIODE(_2247_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5390__C1 (.DIODE(_2247_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5408__B1 (.DIODE(_2264_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5684__A1 (.DIODE(_2275_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5432__A2 (.DIODE(_2275_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5435__B2 (.DIODE(_2291_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6440__B2 (.DIODE(_2292_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5768__A1 (.DIODE(_2292_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5436__A1 (.DIODE(_2292_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5731__A2 (.DIODE(_2296_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5701__A2 (.DIODE(_2296_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5671__A2 (.DIODE(_2296_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5641__A2 (.DIODE(_2296_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5632__A2 (.DIODE(_2296_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5578__A2 (.DIODE(_2296_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5544__A2 (.DIODE(_2296_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5533__A2 (.DIODE(_2296_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5481__A2 (.DIODE(_2296_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5445__A2 (.DIODE(_2296_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5729__B1 (.DIODE(_2297_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5699__B1 (.DIODE(_2297_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5669__B1 (.DIODE(_2297_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5639__B1 (.DIODE(_2297_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5630__B1 (.DIODE(_2297_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5576__B1 (.DIODE(_2297_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5542__B1 (.DIODE(_2297_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5531__B1 (.DIODE(_2297_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5479__B1 (.DIODE(_2297_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5443__B1 (.DIODE(_2297_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5445__B1 (.DIODE(_2300_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5716__A1 (.DIODE(_2311_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5466__A2 (.DIODE(_2311_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5470__B2 (.DIODE(_2325_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6447__B2 (.DIODE(_2326_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5771__A1 (.DIODE(_2326_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5471__A1 (.DIODE(_2326_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6655__C (.DIODE(_2331_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5729__A2 (.DIODE(_2331_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5699__A2 (.DIODE(_2331_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5669__A2 (.DIODE(_2331_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5639__A2 (.DIODE(_2331_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5630__A2 (.DIODE(_2331_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5576__A2 (.DIODE(_2331_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5542__A2 (.DIODE(_2331_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5531__A2 (.DIODE(_2331_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5479__A2 (.DIODE(_2331_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6559__B (.DIODE(_2332_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5730__B1 (.DIODE(_2332_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5700__B1 (.DIODE(_2332_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5670__B1 (.DIODE(_2332_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5640__B1 (.DIODE(_2332_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5631__B1 (.DIODE(_2332_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5577__B1 (.DIODE(_2332_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5543__B1 (.DIODE(_2332_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5532__B1 (.DIODE(_2332_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5478__B1 (.DIODE(_2332_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5505__C (.DIODE(_2352_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5508__B2 (.DIODE(_2362_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6451__B1 (.DIODE(_2363_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5773__A1 (.DIODE(_2363_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5509__A1 (.DIODE(_2363_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5716__A2 (.DIODE(_2370_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5684__A2 (.DIODE(_2370_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5521__B2 (.DIODE(_2370_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5521__C1 (.DIODE(_2374_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5526__B1 (.DIODE(_2376_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5529__B2 (.DIODE(_2382_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6460__A2 (.DIODE(_2383_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5775__A1 (.DIODE(_2383_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5537__A2 (.DIODE(_2383_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5566__C1 (.DIODE(_2418_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5570__B2 (.DIODE(_2422_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6466__A2 (.DIODE(_2423_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5777__A1 (.DIODE(_2423_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5571__A1 (.DIODE(_2423_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5595__A2 (.DIODE(_2441_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5602__B2 (.DIODE(_2453_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6473__A2 (.DIODE(_2454_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5779__A1 (.DIODE(_2454_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5603__A1 (.DIODE(_2454_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5768__S (.DIODE(_2457_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5766__S (.DIODE(_2457_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5764__S (.DIODE(_2457_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5762__S (.DIODE(_2457_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5760__S (.DIODE(_2457_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5758__S (.DIODE(_2457_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5756__S (.DIODE(_2457_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5726__S (.DIODE(_2457_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5696__S (.DIODE(_2457_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5606__S (.DIODE(_2457_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5621__A2 (.DIODE(_2467_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5628__B2 (.DIODE(_2478_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6480__A2 (.DIODE(_2479_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5781__A1 (.DIODE(_2479_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5636__A2 (.DIODE(_2479_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6483__C1 (.DIODE(_2492_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5643__B1_N (.DIODE(_2492_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5659__D (.DIODE(_2508_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5662__B2 (.DIODE(_2511_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6483__B1 (.DIODE(_2512_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5663__A (.DIODE(_2512_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5689__B1 (.DIODE(_2533_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5689__C1 (.DIODE(_2537_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5693__B2 (.DIODE(_2541_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6487__B1 (.DIODE(_2542_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5785__A1 (.DIODE(_2542_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5694__A1 (.DIODE(_2542_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6495__C1 (.DIODE(_2550_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5703__B1_N (.DIODE(_2550_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5717__B1_N (.DIODE(_2564_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6551__A (.DIODE(_2566_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6519__A (.DIODE(_2566_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5720__A2 (.DIODE(_2566_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5722__B1 (.DIODE(_2568_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6495__B1 (.DIODE(_2570_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5723__A (.DIODE(_2570_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5787__A1 (.DIODE(_2571_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5724__A1 (.DIODE(_2571_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5744__B1 (.DIODE(_2586_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5748__B1 (.DIODE(_2591_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6551__B (.DIODE(_2596_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6533__A1 (.DIODE(_2596_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6527__A0 (.DIODE(_2596_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6519__B (.DIODE(_2596_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5751__A2 (.DIODE(_2596_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6506__A2 (.DIODE(_2600_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5789__A1 (.DIODE(_2600_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5754__A1 (.DIODE(_2600_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5789__S (.DIODE(_2610_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5787__S (.DIODE(_2610_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5785__S (.DIODE(_2610_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5783__S (.DIODE(_2610_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5781__S (.DIODE(_2610_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5779__S (.DIODE(_2610_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5777__S (.DIODE(_2610_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5775__S (.DIODE(_2610_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5773__S (.DIODE(_2610_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5771__S (.DIODE(_2610_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5859__A1 (.DIODE(_2634_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5854__A1 (.DIODE(_2634_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5849__A1 (.DIODE(_2634_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5844__A1 (.DIODE(_2634_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5839__A1 (.DIODE(_2634_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5834__A1 (.DIODE(_2634_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5829__A1 (.DIODE(_2634_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5823__A1 (.DIODE(_2634_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6126__A1 (.DIODE(_2637_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6088__A1 (.DIODE(_2637_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6050__A1 (.DIODE(_2637_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6013__A1 (.DIODE(_2637_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5975__A1 (.DIODE(_2637_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5938__A1 (.DIODE(_2637_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5899__A1 (.DIODE(_2637_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5823__A2 (.DIODE(_2637_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5860__A (.DIODE(_2638_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5858__B (.DIODE(_2638_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5853__B (.DIODE(_2638_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5848__B (.DIODE(_2638_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5843__B (.DIODE(_2638_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5821__A (.DIODE(_2638_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5893__A (.DIODE(_2639_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5889__A (.DIODE(_2639_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5885__A (.DIODE(_2639_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5881__A (.DIODE(_2639_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5876__A (.DIODE(_2639_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5873__A (.DIODE(_2639_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5838__B (.DIODE(_2639_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5833__B (.DIODE(_2639_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5827__B (.DIODE(_2639_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5822__B (.DIODE(_2639_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6128__A1 (.DIODE(_2643_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6090__A1 (.DIODE(_2643_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6053__A1 (.DIODE(_2643_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6015__A1 (.DIODE(_2643_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5977__A1 (.DIODE(_2643_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5940__A1 (.DIODE(_2643_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5901__A1 (.DIODE(_2643_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5829__A2 (.DIODE(_2643_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5874__C1 (.DIODE(_2645_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5870__C1 (.DIODE(_2645_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5866__C1 (.DIODE(_2645_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5859__C1 (.DIODE(_2645_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5854__C1 (.DIODE(_2645_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5849__C1 (.DIODE(_2645_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5844__C1 (.DIODE(_2645_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5839__C1 (.DIODE(_2645_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5834__C1 (.DIODE(_2645_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5829__C1 (.DIODE(_2645_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6130__A1 (.DIODE(_2648_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6092__A1 (.DIODE(_2648_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6055__A1 (.DIODE(_2648_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6017__A1 (.DIODE(_2648_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5979__A1 (.DIODE(_2648_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5942__A1 (.DIODE(_2648_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5903__A1 (.DIODE(_2648_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5834__A2 (.DIODE(_2648_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6132__A1 (.DIODE(_2652_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6094__A1 (.DIODE(_2652_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6057__A1 (.DIODE(_2652_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6019__A1 (.DIODE(_2652_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5982__A1 (.DIODE(_2652_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5944__A1 (.DIODE(_2652_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5905__A1 (.DIODE(_2652_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5839__A2 (.DIODE(_2652_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6136__A1 (.DIODE(_2660_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6099__A1 (.DIODE(_2660_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6061__A1 (.DIODE(_2660_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6023__A1 (.DIODE(_2660_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5986__A1 (.DIODE(_2660_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5948__A1 (.DIODE(_2660_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5910__A1 (.DIODE(_2660_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5849__A2 (.DIODE(_2660_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6138__A1 (.DIODE(_2664_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6101__A1 (.DIODE(_2664_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6063__A1 (.DIODE(_2664_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6025__A1 (.DIODE(_2664_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5988__A1 (.DIODE(_2664_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5950__A1 (.DIODE(_2664_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5912__A1 (.DIODE(_2664_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5854__A2 (.DIODE(_2664_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6140__A1 (.DIODE(_2668_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6103__A1 (.DIODE(_2668_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6065__A1 (.DIODE(_2668_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6028__A1 (.DIODE(_2668_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5990__A1 (.DIODE(_2668_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5952__A1 (.DIODE(_2668_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5914__A1 (.DIODE(_2668_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5859__A2 (.DIODE(_2668_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5894__A2 (.DIODE(_2670_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5890__A2 (.DIODE(_2670_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5886__A2 (.DIODE(_2670_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5882__A2 (.DIODE(_2670_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5878__A2 (.DIODE(_2670_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5874__A2 (.DIODE(_2670_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5870__A2 (.DIODE(_2670_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5869__A (.DIODE(_2670_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5866__A2 (.DIODE(_2670_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5865__A (.DIODE(_2670_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5892__A2_N (.DIODE(_2672_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5888__A2_N (.DIODE(_2672_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5884__A2_N (.DIODE(_2672_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5880__A2_N (.DIODE(_2672_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5875__A2_N (.DIODE(_2672_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5872__A2_N (.DIODE(_2672_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5868__A2_N (.DIODE(_2672_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5864__A2_N (.DIODE(_2672_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6142__A (.DIODE(_2674_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6105__A (.DIODE(_2674_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6067__A (.DIODE(_2674_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6030__A (.DIODE(_2674_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5992__A (.DIODE(_2674_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5954__A (.DIODE(_2674_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5916__A (.DIODE(_2674_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5865__B (.DIODE(_2674_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6144__A (.DIODE(_2677_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6107__A (.DIODE(_2677_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6069__A (.DIODE(_2677_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6032__A (.DIODE(_2677_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5994__A (.DIODE(_2677_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5956__A (.DIODE(_2677_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5918__A (.DIODE(_2677_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5869__B (.DIODE(_2677_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6147__A (.DIODE(_2680_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6109__A (.DIODE(_2680_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6071__A (.DIODE(_2680_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6034__A (.DIODE(_2680_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5996__A (.DIODE(_2680_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5959__A (.DIODE(_2680_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5920__A (.DIODE(_2680_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5873__B (.DIODE(_2680_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6149__A (.DIODE(_2682_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6111__A (.DIODE(_2682_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6073__A (.DIODE(_2682_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6036__A (.DIODE(_2682_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5998__A (.DIODE(_2682_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5961__A (.DIODE(_2682_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5922__A (.DIODE(_2682_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5876__B (.DIODE(_2682_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5907__C1 (.DIODE(_2684_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5905__C1 (.DIODE(_2684_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5903__C1 (.DIODE(_2684_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5901__C1 (.DIODE(_2684_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5899__C1 (.DIODE(_2684_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5894__C1 (.DIODE(_2684_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5890__C1 (.DIODE(_2684_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5886__C1 (.DIODE(_2684_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5882__C1 (.DIODE(_2684_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5878__C1 (.DIODE(_2684_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6151__A (.DIODE(_2686_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6113__A (.DIODE(_2686_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6076__A (.DIODE(_2686_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6038__A (.DIODE(_2686_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6000__A (.DIODE(_2686_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5963__A (.DIODE(_2686_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5924__A (.DIODE(_2686_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5881__B (.DIODE(_2686_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6153__A (.DIODE(_2689_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6115__A (.DIODE(_2689_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6078__A (.DIODE(_2689_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6040__A (.DIODE(_2689_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6002__A (.DIODE(_2689_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5965__A (.DIODE(_2689_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5926__A (.DIODE(_2689_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5885__B (.DIODE(_2689_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6155__A (.DIODE(_2692_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6117__A (.DIODE(_2692_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6080__A (.DIODE(_2692_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6042__A (.DIODE(_2692_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6005__A (.DIODE(_2692_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5967__A (.DIODE(_2692_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5928__A (.DIODE(_2692_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5889__B (.DIODE(_2692_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6157__A (.DIODE(_2695_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6119__A (.DIODE(_2695_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6082__A (.DIODE(_2695_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6044__A (.DIODE(_2695_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6007__A (.DIODE(_2695_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5969__A (.DIODE(_2695_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5930__A (.DIODE(_2695_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5893__B (.DIODE(_2695_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5914__A2 (.DIODE(_2697_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5912__A2 (.DIODE(_2697_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5910__A2 (.DIODE(_2697_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5907__A2 (.DIODE(_2697_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5905__A2 (.DIODE(_2697_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5903__A2 (.DIODE(_2697_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5901__A2 (.DIODE(_2697_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5899__A2 (.DIODE(_2697_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5915__A (.DIODE(_2698_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5913__B (.DIODE(_2698_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5911__B (.DIODE(_2698_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5908__B (.DIODE(_2698_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5906__B (.DIODE(_2698_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5897__A (.DIODE(_2698_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5930__B (.DIODE(_2699_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5928__B (.DIODE(_2699_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5926__B (.DIODE(_2699_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5924__B (.DIODE(_2699_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5922__B (.DIODE(_2699_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5920__B (.DIODE(_2699_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5904__B (.DIODE(_2699_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5902__B (.DIODE(_2699_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5900__B (.DIODE(_2699_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5898__B (.DIODE(_2699_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5929__C1 (.DIODE(_2706_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5927__C1 (.DIODE(_2706_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5925__C1 (.DIODE(_2706_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5923__C1 (.DIODE(_2706_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5921__C1 (.DIODE(_2706_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5919__C1 (.DIODE(_2706_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5917__C1 (.DIODE(_2706_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5914__C1 (.DIODE(_2706_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5912__C1 (.DIODE(_2706_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5910__C1 (.DIODE(_2706_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5933__A2 (.DIODE(_2709_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5929__A2 (.DIODE(_2709_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5927__A2 (.DIODE(_2709_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5925__A2 (.DIODE(_2709_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5923__A2 (.DIODE(_2709_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5921__A2 (.DIODE(_2709_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5919__A2 (.DIODE(_2709_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5918__B (.DIODE(_2709_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5917__A2 (.DIODE(_2709_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5916__B (.DIODE(_2709_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6145__A (.DIODE(_2718_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6120__A (.DIODE(_2718_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6098__A (.DIODE(_2718_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6074__A (.DIODE(_2718_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6052__A (.DIODE(_2718_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6027__A (.DIODE(_2718_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6003__A (.DIODE(_2718_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5981__A (.DIODE(_2718_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5957__A (.DIODE(_2718_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5932__A (.DIODE(_2718_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5955__C1 (.DIODE(_2719_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5952__C1 (.DIODE(_2719_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5950__C1 (.DIODE(_2719_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5948__C1 (.DIODE(_2719_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5946__C1 (.DIODE(_2719_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5944__C1 (.DIODE(_2719_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5942__C1 (.DIODE(_2719_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5940__C1 (.DIODE(_2719_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5938__C1 (.DIODE(_2719_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5933__C1 (.DIODE(_2719_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5952__A2 (.DIODE(_2720_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5950__A2 (.DIODE(_2720_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5948__A2 (.DIODE(_2720_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5946__A2 (.DIODE(_2720_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5944__A2 (.DIODE(_2720_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5942__A2 (.DIODE(_2720_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5940__A2 (.DIODE(_2720_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5938__A2 (.DIODE(_2720_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5953__A (.DIODE(_2721_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5951__B (.DIODE(_2721_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5949__B (.DIODE(_2721_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5947__B (.DIODE(_2721_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5945__B (.DIODE(_2721_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5936__A (.DIODE(_2721_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5969__B (.DIODE(_2722_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5967__B (.DIODE(_2722_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5965__B (.DIODE(_2722_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5963__B (.DIODE(_2722_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5961__B (.DIODE(_2722_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5959__B (.DIODE(_2722_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5943__B (.DIODE(_2722_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5941__B (.DIODE(_2722_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5939__B (.DIODE(_2722_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5937__B (.DIODE(_2722_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5970__A2 (.DIODE(_2731_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5968__A2 (.DIODE(_2731_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5966__A2 (.DIODE(_2731_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5964__A2 (.DIODE(_2731_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5962__A2 (.DIODE(_2731_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5960__A2 (.DIODE(_2731_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5958__A2 (.DIODE(_2731_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5956__B (.DIODE(_2731_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5955__A2 (.DIODE(_2731_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5954__B (.DIODE(_2731_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5979__C1 (.DIODE(_2734_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5977__C1 (.DIODE(_2734_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5975__C1 (.DIODE(_2734_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5970__C1 (.DIODE(_2734_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5968__C1 (.DIODE(_2734_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5966__C1 (.DIODE(_2734_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5964__C1 (.DIODE(_2734_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5962__C1 (.DIODE(_2734_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5960__C1 (.DIODE(_2734_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5958__C1 (.DIODE(_2734_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5990__A2 (.DIODE(_2741_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5988__A2 (.DIODE(_2741_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5986__A2 (.DIODE(_2741_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5984__A2 (.DIODE(_2741_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5982__A2 (.DIODE(_2741_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5979__A2 (.DIODE(_2741_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5977__A2 (.DIODE(_2741_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5975__A2 (.DIODE(_2741_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5991__A (.DIODE(_2742_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5989__B (.DIODE(_2742_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5987__B (.DIODE(_2742_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5985__B (.DIODE(_2742_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5983__B (.DIODE(_2742_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5973__A (.DIODE(_2742_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6007__B (.DIODE(_2743_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6005__B (.DIODE(_2743_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6002__B (.DIODE(_2743_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6000__B (.DIODE(_2743_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5998__B (.DIODE(_2743_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5996__B (.DIODE(_2743_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5980__B (.DIODE(_2743_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5978__B (.DIODE(_2743_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5976__B (.DIODE(_2743_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5974__B (.DIODE(_2743_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6001__C1 (.DIODE(_2748_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5999__C1 (.DIODE(_2748_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5997__C1 (.DIODE(_2748_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5995__C1 (.DIODE(_2748_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5993__C1 (.DIODE(_2748_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5990__C1 (.DIODE(_2748_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5988__C1 (.DIODE(_2748_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5986__C1 (.DIODE(_2748_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5984__C1 (.DIODE(_2748_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5982__C1 (.DIODE(_2748_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6025__C1 (.DIODE(_2760_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6023__C1 (.DIODE(_2760_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6021__C1 (.DIODE(_2760_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6019__C1 (.DIODE(_2760_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6017__C1 (.DIODE(_2760_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6015__C1 (.DIODE(_2760_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6013__C1 (.DIODE(_2760_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6008__C1 (.DIODE(_2760_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6006__C1 (.DIODE(_2760_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6004__C1 (.DIODE(_2760_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6028__A2 (.DIODE(_2763_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6025__A2 (.DIODE(_2763_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6023__A2 (.DIODE(_2763_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6021__A2 (.DIODE(_2763_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6019__A2 (.DIODE(_2763_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6017__A2 (.DIODE(_2763_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6015__A2 (.DIODE(_2763_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6013__A2 (.DIODE(_2763_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6029__A (.DIODE(_2764_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6026__B (.DIODE(_2764_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6024__B (.DIODE(_2764_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6022__B (.DIODE(_2764_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6020__B (.DIODE(_2764_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6011__A (.DIODE(_2764_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6044__B (.DIODE(_2765_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6042__B (.DIODE(_2765_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6040__B (.DIODE(_2765_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6038__B (.DIODE(_2765_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6036__B (.DIODE(_2765_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6034__B (.DIODE(_2765_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6018__B (.DIODE(_2765_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6016__B (.DIODE(_2765_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6014__B (.DIODE(_2765_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6012__B (.DIODE(_2765_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6050__C1 (.DIODE(_2774_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6045__C1 (.DIODE(_2774_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6043__C1 (.DIODE(_2774_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6041__C1 (.DIODE(_2774_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6039__C1 (.DIODE(_2774_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6037__C1 (.DIODE(_2774_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6035__C1 (.DIODE(_2774_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6033__C1 (.DIODE(_2774_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6031__C1 (.DIODE(_2774_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6028__C1 (.DIODE(_2774_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6045__A2 (.DIODE(_2775_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6043__A2 (.DIODE(_2775_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6041__A2 (.DIODE(_2775_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6039__A2 (.DIODE(_2775_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6037__A2 (.DIODE(_2775_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6035__A2 (.DIODE(_2775_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6033__A2 (.DIODE(_2775_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6032__B (.DIODE(_2775_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6031__A2 (.DIODE(_2775_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6030__B (.DIODE(_2775_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6065__A2 (.DIODE(_2784_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6063__A2 (.DIODE(_2784_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6061__A2 (.DIODE(_2784_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6059__A2 (.DIODE(_2784_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6057__A2 (.DIODE(_2784_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6055__A2 (.DIODE(_2784_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6053__A2 (.DIODE(_2784_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6050__A2 (.DIODE(_2784_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6066__A (.DIODE(_2785_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6064__B (.DIODE(_2785_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6062__B (.DIODE(_2785_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6060__B (.DIODE(_2785_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6058__B (.DIODE(_2785_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6048__A (.DIODE(_2785_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6082__B (.DIODE(_2786_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6080__B (.DIODE(_2786_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6078__B (.DIODE(_2786_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6076__B (.DIODE(_2786_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6073__B (.DIODE(_2786_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6071__B (.DIODE(_2786_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6056__B (.DIODE(_2786_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6054__B (.DIODE(_2786_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6051__B (.DIODE(_2786_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6049__B (.DIODE(_2786_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6072__C1 (.DIODE(_2789_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6070__C1 (.DIODE(_2789_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6068__C1 (.DIODE(_2789_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6065__C1 (.DIODE(_2789_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6063__C1 (.DIODE(_2789_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6061__C1 (.DIODE(_2789_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6059__C1 (.DIODE(_2789_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6057__C1 (.DIODE(_2789_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6055__C1 (.DIODE(_2789_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6053__C1 (.DIODE(_2789_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6083__A2 (.DIODE(_2796_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6081__A2 (.DIODE(_2796_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6079__A2 (.DIODE(_2796_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6077__A2 (.DIODE(_2796_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6075__A2 (.DIODE(_2796_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6072__A2 (.DIODE(_2796_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6070__A2 (.DIODE(_2796_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6069__B (.DIODE(_2796_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6068__A2 (.DIODE(_2796_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6067__B (.DIODE(_2796_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6096__C1 (.DIODE(_2801_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6094__C1 (.DIODE(_2801_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6092__C1 (.DIODE(_2801_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6090__C1 (.DIODE(_2801_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6088__C1 (.DIODE(_2801_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6083__C1 (.DIODE(_2801_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6081__C1 (.DIODE(_2801_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6079__C1 (.DIODE(_2801_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6077__C1 (.DIODE(_2801_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6075__C1 (.DIODE(_2801_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6103__A2 (.DIODE(_2806_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6101__A2 (.DIODE(_2806_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6099__A2 (.DIODE(_2806_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6096__A2 (.DIODE(_2806_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6094__A2 (.DIODE(_2806_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6092__A2 (.DIODE(_2806_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6090__A2 (.DIODE(_2806_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6088__A2 (.DIODE(_2806_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6104__A (.DIODE(_2807_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6102__B (.DIODE(_2807_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6100__B (.DIODE(_2807_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6097__B (.DIODE(_2807_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6095__B (.DIODE(_2807_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6086__A (.DIODE(_2807_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6119__B (.DIODE(_2808_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6117__B (.DIODE(_2808_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6115__B (.DIODE(_2808_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6113__B (.DIODE(_2808_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6111__B (.DIODE(_2808_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6109__B (.DIODE(_2808_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6093__B (.DIODE(_2808_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6091__B (.DIODE(_2808_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6089__B (.DIODE(_2808_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6087__B (.DIODE(_2808_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6118__C1 (.DIODE(_2815_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6116__C1 (.DIODE(_2815_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6114__C1 (.DIODE(_2815_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6112__C1 (.DIODE(_2815_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6110__C1 (.DIODE(_2815_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6108__C1 (.DIODE(_2815_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6106__C1 (.DIODE(_2815_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6103__C1 (.DIODE(_2815_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6101__C1 (.DIODE(_2815_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6099__C1 (.DIODE(_2815_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6121__A2 (.DIODE(_2818_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6118__A2 (.DIODE(_2818_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6116__A2 (.DIODE(_2818_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6114__A2 (.DIODE(_2818_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6112__A2 (.DIODE(_2818_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6110__A2 (.DIODE(_2818_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6108__A2 (.DIODE(_2818_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6107__B (.DIODE(_2818_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6106__A2 (.DIODE(_2818_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6105__B (.DIODE(_2818_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6143__C1 (.DIODE(_2827_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6140__C1 (.DIODE(_2827_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6138__C1 (.DIODE(_2827_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6136__C1 (.DIODE(_2827_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6134__C1 (.DIODE(_2827_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6132__C1 (.DIODE(_2827_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6130__C1 (.DIODE(_2827_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6128__C1 (.DIODE(_2827_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6126__C1 (.DIODE(_2827_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6121__C1 (.DIODE(_2827_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6141__A (.DIODE(_2829_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6139__B (.DIODE(_2829_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6137__B (.DIODE(_2829_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6135__B (.DIODE(_2829_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6133__B (.DIODE(_2829_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6124__A (.DIODE(_2829_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6157__B (.DIODE(_2830_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6155__B (.DIODE(_2830_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6153__B (.DIODE(_2830_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6151__B (.DIODE(_2830_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6149__B (.DIODE(_2830_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6147__B (.DIODE(_2830_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6131__B (.DIODE(_2830_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6129__B (.DIODE(_2830_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6127__B (.DIODE(_2830_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6125__B (.DIODE(_2830_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6158__A2 (.DIODE(_2839_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6156__A2 (.DIODE(_2839_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6154__A2 (.DIODE(_2839_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6152__A2 (.DIODE(_2839_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6150__A2 (.DIODE(_2839_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6148__A2 (.DIODE(_2839_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6146__A2 (.DIODE(_2839_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6144__B (.DIODE(_2839_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6143__A2 (.DIODE(_2839_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6142__B (.DIODE(_2839_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6572__C1 (.DIODE(_2842_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6568__C1 (.DIODE(_2842_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6522__C1 (.DIODE(_2842_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6158__C1 (.DIODE(_2842_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6156__C1 (.DIODE(_2842_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6154__C1 (.DIODE(_2842_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6152__C1 (.DIODE(_2842_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6150__C1 (.DIODE(_2842_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6148__C1 (.DIODE(_2842_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6146__C1 (.DIODE(_2842_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6297__A (.DIODE(_2851_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6230__A (.DIODE(_2851_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6209__A1 (.DIODE(_2851_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6163__B1 (.DIODE(_2851_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6222__A (.DIODE(_2855_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6189__B (.DIODE(_2855_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6188__B (.DIODE(_2855_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6177__A1 (.DIODE(_2855_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6175__A1 (.DIODE(_2855_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6170__A1 (.DIODE(_2855_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6168__A (.DIODE(_2855_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6198__B1 (.DIODE(_2868_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6186__B (.DIODE(_2868_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6181__B (.DIODE(_2868_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6358__S (.DIODE(_2870_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6347__S (.DIODE(_2870_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6339__S (.DIODE(_2870_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6324__S (.DIODE(_2870_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6286__S (.DIODE(_2870_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6275__S (.DIODE(_2870_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6263__S (.DIODE(_2870_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6208__B1 (.DIODE(_2870_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6183__A (.DIODE(_2870_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6312__A2 (.DIODE(_2871_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6299__A2 (.DIODE(_2871_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6298__B1 (.DIODE(_2871_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6250__S (.DIODE(_2871_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6243__A2 (.DIODE(_2871_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6232__S (.DIODE(_2871_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6219__S (.DIODE(_2871_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6210__A2 (.DIODE(_2871_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6201__A2 (.DIODE(_2871_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6192__A2 (.DIODE(_2871_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6357__B2 (.DIODE(_2872_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6346__A2 (.DIODE(_2872_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6274__B2 (.DIODE(_2872_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6262__B2 (.DIODE(_2872_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6249__A2 (.DIODE(_2872_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6185__A (.DIODE(_2872_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6338__B2 (.DIODE(_2873_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6323__B2 (.DIODE(_2873_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6298__A2 (.DIODE(_2873_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6285__B2 (.DIODE(_2873_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6243__B1 (.DIODE(_2873_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6231__A2 (.DIODE(_2873_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6218__B2 (.DIODE(_2873_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6208__A2 (.DIODE(_2873_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6201__B1 (.DIODE(_2873_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6192__B1 (.DIODE(_2873_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6406__A1 (.DIODE(_2877_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6384__A2 (.DIODE(_2877_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6352__A2 (.DIODE(_2877_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6190__A2 (.DIODE(_2877_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6357__A1 (.DIODE(_2886_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6346__B2 (.DIODE(_2886_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6338__A1 (.DIODE(_2886_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6323__A1 (.DIODE(_2886_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6311__A (.DIODE(_2886_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6285__A1 (.DIODE(_2886_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6261__A (.DIODE(_2886_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6249__B2 (.DIODE(_2886_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6218__A1 (.DIODE(_2886_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6200__C1 (.DIODE(_2886_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6301__A2 (.DIODE(_2897_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6253__A (.DIODE(_2897_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6214__A3 (.DIODE(_2897_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6213__D (.DIODE(_2897_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6315__A2 (.DIODE(_2908_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6226__A2 (.DIODE(_2908_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6225__C (.DIODE(_2908_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6327__B (.DIODE(_2920_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6239__A2 (.DIODE(_2920_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6238__A (.DIODE(_2920_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6353__A2 (.DIODE(_2936_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6257__A2 (.DIODE(_2936_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6256__C (.DIODE(_2936_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6404__B (.DIODE(_3023_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6393__A2 (.DIODE(_3023_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6382__B (.DIODE(_3023_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6370__A2 (.DIODE(_3023_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6351__A1 (.DIODE(_3023_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6401__A2 (.DIODE(_3034_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6390__A2 (.DIODE(_3034_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6379__A2 (.DIODE(_3034_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6367__A2 (.DIODE(_3034_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6506__C1 (.DIODE(_3063_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6501__S (.DIODE(_3063_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6484__B1 (.DIODE(_3063_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6480__C1 (.DIODE(_3063_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6478__B1_N (.DIODE(_3063_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6473__C1 (.DIODE(_3063_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6466__C1 (.DIODE(_3063_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6460__C1 (.DIODE(_3063_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6431__C1 (.DIODE(_3063_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6409__A (.DIODE(_3063_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6494__A1 (.DIODE(_3064_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6493__A (.DIODE(_3064_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6486__A1 (.DIODE(_3064_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6455__A1 (.DIODE(_3064_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6450__A1 (.DIODE(_3064_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6449__A (.DIODE(_3064_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6445__A1 (.DIODE(_3064_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6444__B1 (.DIODE(_3064_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6417__A1 (.DIODE(_3064_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6414__A (.DIODE(_3064_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6495__A2 (.DIODE(_3065_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6483__A2 (.DIODE(_3065_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6465__A2 (.DIODE(_3065_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6446__B (.DIODE(_3065_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6439__B (.DIODE(_3065_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6412__A2 (.DIODE(_3065_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6495__B2 (.DIODE(_3066_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6483__B2 (.DIODE(_3066_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6434__A (.DIODE(_3066_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6424__A1 (.DIODE(_3066_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6412__B2 (.DIODE(_3066_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6698__B1 (.DIODE(_3070_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6692__B1 (.DIODE(_3070_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6507__A (.DIODE(_3070_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6481__A (.DIODE(_3070_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6474__A (.DIODE(_3070_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6467__A (.DIODE(_3070_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6461__A (.DIODE(_3070_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6432__A (.DIODE(_3070_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6416__A (.DIODE(_3070_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6697__B1 (.DIODE(_3071_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6696__B1 (.DIODE(_3071_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6494__C1 (.DIODE(_3071_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6486__C1 (.DIODE(_3071_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6455__C1 (.DIODE(_3071_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6450__C1 (.DIODE(_3071_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6445__C1 (.DIODE(_3071_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6438__C1 (.DIODE(_3071_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6425__B1 (.DIODE(_3071_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6417__C1 (.DIODE(_3071_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6506__A1 (.DIODE(_3082_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6487__B2 (.DIODE(_3082_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6480__A1 (.DIODE(_3082_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6473__A1 (.DIODE(_3082_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6466__A1 (.DIODE(_3082_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6460__A1 (.DIODE(_3082_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6451__B2 (.DIODE(_3082_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6447__B1 (.DIODE(_3082_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6440__B1 (.DIODE(_3082_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6431__A1 (.DIODE(_3082_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6496__B (.DIODE(_3092_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6491__B (.DIODE(_3092_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6442__A2 (.DIODE(_3092_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6502__B (.DIODE(_3143_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6557__A1 (.DIODE(_3150_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6556__B (.DIODE(_3150_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6535__B (.DIODE(_3150_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6532__B1 (.DIODE(_3150_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6527__S (.DIODE(_3150_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6523__S (.DIODE(_3150_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6520__B (.DIODE(_3150_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6516__A (.DIODE(_3150_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6511__A2 (.DIODE(_3150_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6634__A2 (.DIODE(_3196_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6630__A2 (.DIODE(_3196_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6626__A2 (.DIODE(_3196_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6622__A2 (.DIODE(_3196_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6617__A2 (.DIODE(_3196_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6613__A2 (.DIODE(_3196_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6562__A (.DIODE(_3196_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6609__A2 (.DIODE(_3197_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6605__A2 (.DIODE(_3197_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6601__A2 (.DIODE(_3197_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6597__A2 (.DIODE(_3197_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6593__A2 (.DIODE(_3197_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6589__A2 (.DIODE(_3197_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6585__A2 (.DIODE(_3197_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6581__A2 (.DIODE(_3197_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6572__A2 (.DIODE(_3197_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6568__A2 (.DIODE(_3197_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6633__C1 (.DIODE(_3198_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6629__C1 (.DIODE(_3198_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6625__C1 (.DIODE(_3198_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6584__A (.DIODE(_3198_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6578__A (.DIODE(_3198_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6571__A (.DIODE(_3198_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6567__A (.DIODE(_3198_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6632__B (.DIODE(_3200_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6628__B (.DIODE(_3200_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6624__B (.DIODE(_3200_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6619__B (.DIODE(_3200_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6615__B (.DIODE(_3200_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6611__B (.DIODE(_3200_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6576__A (.DIODE(_3200_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6573__A (.DIODE(_3200_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6570__S (.DIODE(_3200_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6566__S (.DIODE(_3200_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6620__A1 (.DIODE(_3206_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6616__A1 (.DIODE(_3206_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6612__A1 (.DIODE(_3206_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6608__A1 (.DIODE(_3206_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6604__A1 (.DIODE(_3206_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6600__A1 (.DIODE(_3206_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6596__A1 (.DIODE(_3206_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6592__A1 (.DIODE(_3206_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6588__A1 (.DIODE(_3206_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6579__A1 (.DIODE(_3206_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6697__A1 (.DIODE(_3207_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6614__S (.DIODE(_3207_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6610__S (.DIODE(_3207_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6606__S (.DIODE(_3207_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6602__S (.DIODE(_3207_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6598__S (.DIODE(_3207_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6594__S (.DIODE(_3207_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6590__S (.DIODE(_3207_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6586__S (.DIODE(_3207_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6575__S (.DIODE(_3207_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6633__A1 (.DIODE(_3209_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6629__A1 (.DIODE(_3209_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6625__A1 (.DIODE(_3209_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6607__B (.DIODE(_3209_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6603__B (.DIODE(_3209_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6599__B (.DIODE(_3209_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6595__B (.DIODE(_3209_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6591__B (.DIODE(_3209_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6587__B (.DIODE(_3209_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6577__B (.DIODE(_3209_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6620__C1 (.DIODE(_3211_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6616__C1 (.DIODE(_3211_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6612__C1 (.DIODE(_3211_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6608__C1 (.DIODE(_3211_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6604__C1 (.DIODE(_3211_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6600__C1 (.DIODE(_3211_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6596__C1 (.DIODE(_3211_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6592__C1 (.DIODE(_3211_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6588__C1 (.DIODE(_3211_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6579__C1 (.DIODE(_3211_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6581__B1 (.DIODE(_3212_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6617__C1 (.DIODE(_3213_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6613__C1 (.DIODE(_3213_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6609__C1 (.DIODE(_3213_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6605__C1 (.DIODE(_3213_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6601__C1 (.DIODE(_3213_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6597__C1 (.DIODE(_3213_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6593__C1 (.DIODE(_3213_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6589__C1 (.DIODE(_3213_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6585__C1 (.DIODE(_3213_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6581__C1 (.DIODE(_3213_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6670__C1 (.DIODE(_3244_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6668__C1 (.DIODE(_3244_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6666__C1 (.DIODE(_3244_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6664__C1 (.DIODE(_3244_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6662__C1 (.DIODE(_3244_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6660__C1 (.DIODE(_3244_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6634__C1 (.DIODE(_3244_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6630__C1 (.DIODE(_3244_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6626__C1 (.DIODE(_3244_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6622__C1 (.DIODE(_3244_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6643__A2 (.DIODE(_3254_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6640__A2 (.DIODE(_3254_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6637__A2 (.DIODE(_3254_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6636__B (.DIODE(_3254_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6690__B (.DIODE(_3268_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6688__B (.DIODE(_3268_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6686__B (.DIODE(_3268_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6684__B (.DIODE(_3268_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6682__B (.DIODE(_3268_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6680__B (.DIODE(_3268_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6658__A (.DIODE(_3268_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6656__A (.DIODE(_3268_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6691__A2 (.DIODE(_3269_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6689__A2 (.DIODE(_3269_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6687__A2 (.DIODE(_3269_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6685__A2 (.DIODE(_3269_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6683__A2 (.DIODE(_3269_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6681__A2 (.DIODE(_3269_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6657__A (.DIODE(_3269_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6679__A2 (.DIODE(_3270_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6677__A2 (.DIODE(_3270_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6675__A2 (.DIODE(_3270_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6673__A2 (.DIODE(_3270_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6670__A2 (.DIODE(_3270_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6668__A2 (.DIODE(_3270_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6666__A2 (.DIODE(_3270_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6664__A2 (.DIODE(_3270_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6662__A2 (.DIODE(_3270_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6660__A2 (.DIODE(_3270_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6678__B (.DIODE(_3271_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6676__B (.DIODE(_3271_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6674__B (.DIODE(_3271_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6671__B (.DIODE(_3271_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6669__B (.DIODE(_3271_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6667__B (.DIODE(_3271_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6665__B (.DIODE(_3271_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6663__B (.DIODE(_3271_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6661__B (.DIODE(_3271_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6659__B (.DIODE(_3271_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6691__C1 (.DIODE(_3279_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6689__C1 (.DIODE(_3279_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6687__C1 (.DIODE(_3279_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6685__C1 (.DIODE(_3279_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6683__C1 (.DIODE(_3279_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6681__C1 (.DIODE(_3279_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6679__C1 (.DIODE(_3279_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6677__C1 (.DIODE(_3279_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6675__C1 (.DIODE(_3279_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6673__C1 (.DIODE(_3279_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6746__A2 (.DIODE(_3292_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6740__A2 (.DIODE(_3292_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6728__A2 (.DIODE(_3292_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6722__A2 (.DIODE(_3292_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6720__B1 (.DIODE(_3292_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6710__A2 (.DIODE(_3292_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6701__C1 (.DIODE(_3292_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6752__B1 (.DIODE(_3295_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6747__A2 (.DIODE(_3295_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6741__A2 (.DIODE(_3295_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6735__A2 (.DIODE(_3295_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6729__A2 (.DIODE(_3295_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6723__A2 (.DIODE(_3295_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6717__B (.DIODE(_3295_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6712__A2 (.DIODE(_3295_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6752__A2 (.DIODE(_3299_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6751__A (.DIODE(_3299_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6745__B1 (.DIODE(_3299_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6739__B1 (.DIODE(_3299_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6734__A1 (.DIODE(_3299_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6733__B (.DIODE(_3299_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6727__B1 (.DIODE(_3299_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6716__S (.DIODE(_3299_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6708__C1 (.DIODE(_3299_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6753__A2 (.DIODE(_3301_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6746__B1 (.DIODE(_3301_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6740__B1 (.DIODE(_3301_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6734__C1 (.DIODE(_3301_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6728__B1 (.DIODE(_3301_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6722__C1 (.DIODE(_3301_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6718__A1 (.DIODE(_3301_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6710__C1 (.DIODE(_3301_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6768__C1 (.DIODE(_3303_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6765__C1 (.DIODE(_3303_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6762__C1 (.DIODE(_3303_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6747__C1 (.DIODE(_3303_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6741__C1 (.DIODE(_3303_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6735__C1 (.DIODE(_3303_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6729__C1 (.DIODE(_3303_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6723__C1 (.DIODE(_3303_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6718__C1 (.DIODE(_3303_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6712__C1 (.DIODE(_3303_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6782__S (.DIODE(_3341_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6779__A (.DIODE(_3341_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6776__A (.DIODE(_3341_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6770__B1 (.DIODE(_3341_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6764__B1 (.DIODE(_3341_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6758__A (.DIODE(_3341_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6780__A2 (.DIODE(_3342_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6777__A2 (.DIODE(_3342_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6774__A2 (.DIODE(_3342_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6773__A (.DIODE(_3342_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6771__A2 (.DIODE(_3342_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6768__A2 (.DIODE(_3342_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6767__A (.DIODE(_3342_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6765__A2 (.DIODE(_3342_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6762__A2 (.DIODE(_3342_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6761__A (.DIODE(_3342_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6781__S (.DIODE(_3343_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6778__S (.DIODE(_3343_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6775__S (.DIODE(_3343_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6772__S (.DIODE(_3343_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6770__A2 (.DIODE(_3343_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6769__B (.DIODE(_3343_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6766__S (.DIODE(_3343_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6764__A2 (.DIODE(_3343_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6763__B (.DIODE(_3343_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6760__S (.DIODE(_3343_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5401__S (.DIODE(\core_1.dec_mem_access ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4110__A (.DIODE(\core_1.dec_mem_access ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5811__B (.DIODE(\core_1.dec_mem_long ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4132__A1 (.DIODE(\core_1.dec_mem_long ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3579__C1 (.DIODE(\core_1.dec_mem_long ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5809__A0 (.DIODE(\core_1.dec_mem_width ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4131__A1 (.DIODE(\core_1.dec_mem_width ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4457__A (.DIODE(\core_1.dec_r_bus_imm ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4454__A (.DIODE(\core_1.dec_r_bus_imm ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4417__A (.DIODE(\core_1.dec_r_bus_imm ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4399__A (.DIODE(\core_1.dec_r_bus_imm ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4395__A (.DIODE(\core_1.dec_r_bus_imm ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4002__A (.DIODE(\core_1.dec_r_bus_imm ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5545__B (.DIODE(\core_1.dec_sreg_irt ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5482__B (.DIODE(\core_1.dec_sreg_irt ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5409__B (.DIODE(\core_1.dec_sreg_irt ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5281__B1 (.DIODE(\core_1.dec_sreg_irt ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5215__B1 (.DIODE(\core_1.dec_sreg_irt ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4898__B (.DIODE(\core_1.dec_sreg_irt ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4894__A (.DIODE(\core_1.dec_sreg_irt ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3979__A (.DIODE(\core_1.dec_sreg_irt ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6755__A2 (.DIODE(\core_1.dec_sreg_jal_over ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5273__C1 (.DIODE(\core_1.dec_sreg_jal_over ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5261__B1 (.DIODE(\core_1.dec_sreg_jal_over ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5253__A (.DIODE(\core_1.dec_sreg_jal_over ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5217__A (.DIODE(\core_1.dec_sreg_jal_over ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5205__B1 (.DIODE(\core_1.dec_sreg_jal_over ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5192__A (.DIODE(\core_1.dec_sreg_jal_over ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4125__B2 (.DIODE(\core_1.dec_sreg_jal_over ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6700__A (.DIODE(\core_1.dec_sreg_store ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6509__A (.DIODE(\core_1.dec_sreg_store ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4122__A (.DIODE(\core_1.dec_sreg_store ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3996__B (.DIODE(\core_1.dec_sreg_store ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3983__D (.DIODE(\core_1.dec_sreg_store ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3980__A1 (.DIODE(\core_1.dec_sreg_store ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4117__A (.DIODE(\core_1.dec_used_operands[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3589__B1 (.DIODE(\core_1.dec_used_operands[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4120__A1 (.DIODE(\core_1.dec_used_operands[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3559__C1 (.DIODE(\core_1.dec_used_operands[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4345__A1 (.DIODE(\core_1.decode.i_imm_pass[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4077__A1 (.DIODE(\core_1.decode.i_imm_pass[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4347__A1 (.DIODE(\core_1.decode.i_imm_pass[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4079__A1 (.DIODE(\core_1.decode.i_imm_pass[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4349__A1 (.DIODE(\core_1.decode.i_imm_pass[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4081__A1 (.DIODE(\core_1.decode.i_imm_pass[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4351__A1 (.DIODE(\core_1.decode.i_imm_pass[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4083__A1 (.DIODE(\core_1.decode.i_imm_pass[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4307__A1 (.DIODE(\core_1.decode.i_instr_l[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4025__A1 (.DIODE(\core_1.decode.i_instr_l[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3902__B (.DIODE(\core_1.decode.i_instr_l[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3889__A1 (.DIODE(\core_1.decode.i_instr_l[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3852__B (.DIODE(\core_1.decode.i_instr_l[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3832__A (.DIODE(\core_1.decode.i_instr_l[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3823__B (.DIODE(\core_1.decode.i_instr_l[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3820__A (.DIODE(\core_1.decode.i_instr_l[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3813__B (.DIODE(\core_1.decode.i_instr_l[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3806__B (.DIODE(\core_1.decode.i_instr_l[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4328__A1 (.DIODE(\core_1.decode.i_instr_l[10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4074__A1 (.DIODE(\core_1.decode.i_instr_l[10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4043__A1 (.DIODE(\core_1.decode.i_instr_l[10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4031__B2 (.DIODE(\core_1.decode.i_instr_l[10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4331__A1 (.DIODE(\core_1.decode.i_instr_l[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4045__A1 (.DIODE(\core_1.decode.i_instr_l[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4033__B2 (.DIODE(\core_1.decode.i_instr_l[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4334__A1 (.DIODE(\core_1.decode.i_instr_l[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4048__A1 (.DIODE(\core_1.decode.i_instr_l[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4035__B2 (.DIODE(\core_1.decode.i_instr_l[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4337__A1 (.DIODE(\core_1.decode.i_instr_l[13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4043__B2 (.DIODE(\core_1.decode.i_instr_l[13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4031__A1 (.DIODE(\core_1.decode.i_instr_l[13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4340__A1 (.DIODE(\core_1.decode.i_instr_l[14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4045__B2 (.DIODE(\core_1.decode.i_instr_l[14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4033__A1 (.DIODE(\core_1.decode.i_instr_l[14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4343__A1 (.DIODE(\core_1.decode.i_instr_l[15] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4048__B2 (.DIODE(\core_1.decode.i_instr_l[15] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4035__A1 (.DIODE(\core_1.decode.i_instr_l[15] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4309__A1 (.DIODE(\core_1.decode.i_instr_l[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4130__A1 (.DIODE(\core_1.decode.i_instr_l[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3902__A (.DIODE(\core_1.decode.i_instr_l[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3877__A1 (.DIODE(\core_1.decode.i_instr_l[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3852__A (.DIODE(\core_1.decode.i_instr_l[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3831__A (.DIODE(\core_1.decode.i_instr_l[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3823__A (.DIODE(\core_1.decode.i_instr_l[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3821__A (.DIODE(\core_1.decode.i_instr_l[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3813__A (.DIODE(\core_1.decode.i_instr_l[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3805__A (.DIODE(\core_1.decode.i_instr_l[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4321__A1 (.DIODE(\core_1.decode.i_instr_l[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4071__A1 (.DIODE(\core_1.decode.i_instr_l[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4064__B (.DIODE(\core_1.decode.i_instr_l[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4062__A_N (.DIODE(\core_1.decode.i_instr_l[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4060__A (.DIODE(\core_1.decode.i_instr_l[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4055__A_N (.DIODE(\core_1.decode.i_instr_l[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4915__A1 (.DIODE(\core_1.decode.i_jmp_pred_pass ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4393__A0 (.DIODE(\core_1.decode.i_jmp_pred_pass ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6186__A (.DIODE(\core_1.decode.o_submit ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6162__A (.DIODE(\core_1.decode.o_submit ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4605__A (.DIODE(\core_1.decode.o_submit ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3595__A (.DIODE(\core_1.decode.o_submit ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3594__A (.DIODE(\core_1.decode.o_submit ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3552__B (.DIODE(\core_1.decode.o_submit ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5108__A1 (.DIODE(\core_1.decode.oc_alu_mode[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5100__A (.DIODE(\core_1.decode.oc_alu_mode[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5096__A1 (.DIODE(\core_1.decode.oc_alu_mode[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5094__A (.DIODE(\core_1.decode.oc_alu_mode[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4880__D (.DIODE(\core_1.decode.oc_alu_mode[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4846__A (.DIODE(\core_1.decode.oc_alu_mode[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4838__A (.DIODE(\core_1.decode.oc_alu_mode[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4835__A1 (.DIODE(\core_1.decode.oc_alu_mode[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3883__A (.DIODE(\core_1.decode.oc_alu_mode[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5736__A1 (.DIODE(\core_1.decode.oc_alu_mode[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5714__A1 (.DIODE(\core_1.decode.oc_alu_mode[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5681__B2 (.DIODE(\core_1.decode.oc_alu_mode[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5619__A1 (.DIODE(\core_1.decode.oc_alu_mode[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5592__A1 (.DIODE(\core_1.decode.oc_alu_mode[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5236__A1 (.DIODE(\core_1.decode.oc_alu_mode[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4887__A1 (.DIODE(\core_1.decode.oc_alu_mode[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4879__D (.DIODE(\core_1.decode.oc_alu_mode[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3899__A (.DIODE(\core_1.decode.oc_alu_mode[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5518__A (.DIODE(\core_1.decode.oc_alu_mode[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4884__A (.DIODE(\core_1.decode.oc_alu_mode[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4879__C (.DIODE(\core_1.decode.oc_alu_mode[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3898__A1 (.DIODE(\core_1.decode.oc_alu_mode[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5714__B2 (.DIODE(\core_1.decode.oc_alu_mode[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5682__A1 (.DIODE(\core_1.decode.oc_alu_mode[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5619__B2 (.DIODE(\core_1.decode.oc_alu_mode[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5590__A (.DIODE(\core_1.decode.oc_alu_mode[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5342__C1 (.DIODE(\core_1.decode.oc_alu_mode[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5236__B2 (.DIODE(\core_1.decode.oc_alu_mode[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4887__B2 (.DIODE(\core_1.decode.oc_alu_mode[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4880__B (.DIODE(\core_1.decode.oc_alu_mode[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3819__A (.DIODE(\core_1.decode.oc_alu_mode[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5713__A1 (.DIODE(\core_1.decode.oc_alu_mode[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5680__A1 (.DIODE(\core_1.decode.oc_alu_mode[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5618__A1 (.DIODE(\core_1.decode.oc_alu_mode[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5591__A1 (.DIODE(\core_1.decode.oc_alu_mode[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5381__A1 (.DIODE(\core_1.decode.oc_alu_mode[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5235__A1 (.DIODE(\core_1.decode.oc_alu_mode[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4886__A1 (.DIODE(\core_1.decode.oc_alu_mode[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4880__C (.DIODE(\core_1.decode.oc_alu_mode[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3826__A (.DIODE(\core_1.decode.oc_alu_mode[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5713__B2 (.DIODE(\core_1.decode.oc_alu_mode[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5681__A1 (.DIODE(\core_1.decode.oc_alu_mode[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5618__C1 (.DIODE(\core_1.decode.oc_alu_mode[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5233__A (.DIODE(\core_1.decode.oc_alu_mode[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4886__B2 (.DIODE(\core_1.decode.oc_alu_mode[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4879__A (.DIODE(\core_1.decode.oc_alu_mode[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3851__A (.DIODE(\core_1.decode.oc_alu_mode[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5818__A0 (.DIODE(\core_1.ew_data[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5259__A0 (.DIODE(\core_1.ew_data[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3927__A0 (.DIODE(\core_1.ew_data[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3911__A (.DIODE(\core_1.ew_data[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5825__A0 (.DIODE(\core_1.ew_data[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5279__A0 (.DIODE(\core_1.ew_data[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3929__A0 (.DIODE(\core_1.ew_data[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3913__A (.DIODE(\core_1.ew_data[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5831__A0 (.DIODE(\core_1.ew_data[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5325__A0 (.DIODE(\core_1.ew_data[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3931__A0 (.DIODE(\core_1.ew_data[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3915__A (.DIODE(\core_1.ew_data[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5836__A0 (.DIODE(\core_1.ew_data[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5363__A0 (.DIODE(\core_1.ew_data[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3933__A0 (.DIODE(\core_1.ew_data[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3917__A (.DIODE(\core_1.ew_data[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5841__A0 (.DIODE(\core_1.ew_data[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5403__A0 (.DIODE(\core_1.ew_data[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3935__A0 (.DIODE(\core_1.ew_data[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3919__A (.DIODE(\core_1.ew_data[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5846__A0 (.DIODE(\core_1.ew_data[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5438__A0 (.DIODE(\core_1.ew_data[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3937__A0 (.DIODE(\core_1.ew_data[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3921__A (.DIODE(\core_1.ew_data[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5851__A0 (.DIODE(\core_1.ew_data[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5473__A0 (.DIODE(\core_1.ew_data[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3939__A0 (.DIODE(\core_1.ew_data[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3923__A (.DIODE(\core_1.ew_data[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5856__A0 (.DIODE(\core_1.ew_data[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5511__A0 (.DIODE(\core_1.ew_data[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3941__A0 (.DIODE(\core_1.ew_data[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3925__A (.DIODE(\core_1.ew_data[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5861__A_N (.DIODE(\core_1.ew_mem_width ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5809__A1 (.DIODE(\core_1.ew_mem_width ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3943__B_N (.DIODE(\core_1.ew_mem_width ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3908__B (.DIODE(\core_1.ew_mem_width ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6085__A (.DIODE(\core_1.ew_reg_ie[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6084__A (.DIODE(\core_1.ew_reg_ie[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5793__A1 (.DIODE(\core_1.ew_reg_ie[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3584__B2 (.DIODE(\core_1.ew_reg_ie[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3575__A1 (.DIODE(\core_1.ew_reg_ie[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3555__A1 (.DIODE(\core_1.ew_reg_ie[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6047__A (.DIODE(\core_1.ew_reg_ie[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6046__A (.DIODE(\core_1.ew_reg_ie[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5795__A1 (.DIODE(\core_1.ew_reg_ie[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3583__B (.DIODE(\core_1.ew_reg_ie[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3574__B (.DIODE(\core_1.ew_reg_ie[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3555__A2 (.DIODE(\core_1.ew_reg_ie[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6010__A (.DIODE(\core_1.ew_reg_ie[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6009__A (.DIODE(\core_1.ew_reg_ie[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5797__A1 (.DIODE(\core_1.ew_reg_ie[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3585__A1 (.DIODE(\core_1.ew_reg_ie[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3572__B (.DIODE(\core_1.ew_reg_ie[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3555__A3 (.DIODE(\core_1.ew_reg_ie[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5972__A (.DIODE(\core_1.ew_reg_ie[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5971__A (.DIODE(\core_1.ew_reg_ie[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5799__A1 (.DIODE(\core_1.ew_reg_ie[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3587__A1 (.DIODE(\core_1.ew_reg_ie[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3578__A3 (.DIODE(\core_1.ew_reg_ie[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3557__A0 (.DIODE(\core_1.ew_reg_ie[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5935__A (.DIODE(\core_1.ew_reg_ie[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5934__A (.DIODE(\core_1.ew_reg_ie[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5801__A1 (.DIODE(\core_1.ew_reg_ie[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3587__B2 (.DIODE(\core_1.ew_reg_ie[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3578__A0 (.DIODE(\core_1.ew_reg_ie[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3557__A1 (.DIODE(\core_1.ew_reg_ie[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5896__A (.DIODE(\core_1.ew_reg_ie[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5895__A (.DIODE(\core_1.ew_reg_ie[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5803__A1 (.DIODE(\core_1.ew_reg_ie[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3586__B (.DIODE(\core_1.ew_reg_ie[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3578__A1 (.DIODE(\core_1.ew_reg_ie[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3557__A2 (.DIODE(\core_1.ew_reg_ie[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5820__A (.DIODE(\core_1.ew_reg_ie[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5816__A (.DIODE(\core_1.ew_reg_ie[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5805__A1 (.DIODE(\core_1.ew_reg_ie[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3588__A1 (.DIODE(\core_1.ew_reg_ie[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3578__A2 (.DIODE(\core_1.ew_reg_ie[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3557__A3 (.DIODE(\core_1.ew_reg_ie[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6522__A1 (.DIODE(\core_1.execute.alu_flag_reg.o_d[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5207__A (.DIODE(\core_1.execute.alu_flag_reg.o_d[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3966__B (.DIODE(\core_1.execute.alu_flag_reg.o_d[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3963__A1 (.DIODE(\core_1.execute.alu_flag_reg.o_d[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3958__B (.DIODE(\core_1.execute.alu_flag_reg.o_d[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3955__A (.DIODE(\core_1.execute.alu_flag_reg.o_d[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6524__A0 (.DIODE(\core_1.execute.alu_flag_reg.o_d[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5263__A (.DIODE(\core_1.execute.alu_flag_reg.o_d[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4862__A (.DIODE(\core_1.execute.alu_flag_reg.o_d[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3966__A (.DIODE(\core_1.execute.alu_flag_reg.o_d[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3963__B1 (.DIODE(\core_1.execute.alu_flag_reg.o_d[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3960__A0 (.DIODE(\core_1.execute.alu_flag_reg.o_d[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6528__A0 (.DIODE(\core_1.execute.alu_flag_reg.o_d[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5288__A1 (.DIODE(\core_1.execute.alu_flag_reg.o_d[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3960__A1 (.DIODE(\core_1.execute.alu_flag_reg.o_d[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3958__A (.DIODE(\core_1.execute.alu_flag_reg.o_d[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3953__A (.DIODE(\core_1.execute.alu_flag_reg.o_d[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6537__A1 (.DIODE(\core_1.execute.alu_flag_reg.o_d[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5331__A1 (.DIODE(\core_1.execute.alu_flag_reg.o_d[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3964__A (.DIODE(\core_1.execute.alu_flag_reg.o_d[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6212__S0 (.DIODE(\core_1.execute.alu_mul_div.cbit[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6193__C1 (.DIODE(\core_1.execute.alu_mul_div.cbit[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6167__A (.DIODE(\core_1.execute.alu_mul_div.cbit[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4712__B1 (.DIODE(\core_1.execute.alu_mul_div.cbit[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4660__A (.DIODE(\core_1.execute.alu_mul_div.cbit[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4194__A (.DIODE(\core_1.execute.alu_mul_div.cbit[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6223__A (.DIODE(\core_1.execute.alu_mul_div.cbit[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6213__B (.DIODE(\core_1.execute.alu_mul_div.cbit[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6187__B (.DIODE(\core_1.execute.alu_mul_div.cbit[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4665__A (.DIODE(\core_1.execute.alu_mul_div.cbit[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4192__A (.DIODE(\core_1.execute.alu_mul_div.cbit[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6213__A (.DIODE(\core_1.execute.alu_mul_div.cbit[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6204__A1 (.DIODE(\core_1.execute.alu_mul_div.cbit[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6187__A (.DIODE(\core_1.execute.alu_mul_div.cbit[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4664__A (.DIODE(\core_1.execute.alu_mul_div.cbit[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4190__A (.DIODE(\core_1.execute.alu_mul_div.cbit[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6180__B (.DIODE(\core_1.execute.alu_mul_div.comp ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4488__A (.DIODE(\core_1.execute.alu_mul_div.comp ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4200__A (.DIODE(\core_1.execute.alu_mul_div.comp ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3597__A (.DIODE(\core_1.execute.alu_mul_div.comp ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5360__A1 (.DIODE(\core_1.execute.alu_mul_div.div_cur[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4530__A1 (.DIODE(\core_1.execute.alu_mul_div.div_cur[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4525__A1 (.DIODE(\core_1.execute.alu_mul_div.div_cur[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4518__A (.DIODE(\core_1.execute.alu_mul_div.div_cur[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4462__A (.DIODE(\core_1.execute.alu_mul_div.div_cur[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4450__A (.DIODE(\core_1.execute.alu_mul_div.div_cur[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4537__A1 (.DIODE(\core_1.execute.alu_mul_div.div_cur[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4531__A1 (.DIODE(\core_1.execute.alu_mul_div.div_cur[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4445__A (.DIODE(\core_1.execute.alu_mul_div.div_cur[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4439__A (.DIODE(\core_1.execute.alu_mul_div.div_cur[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5470__A1 (.DIODE(\core_1.execute.alu_mul_div.div_cur[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4552__A1 (.DIODE(\core_1.execute.alu_mul_div.div_cur[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4545__A1 (.DIODE(\core_1.execute.alu_mul_div.div_cur[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4434__A (.DIODE(\core_1.execute.alu_mul_div.div_cur[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4433__A (.DIODE(\core_1.execute.alu_mul_div.div_cur[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5508__A1 (.DIODE(\core_1.execute.alu_mul_div.div_cur[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4558__A1 (.DIODE(\core_1.execute.alu_mul_div.div_cur[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4553__A1 (.DIODE(\core_1.execute.alu_mul_div.div_cur[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4547__A (.DIODE(\core_1.execute.alu_mul_div.div_cur[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4469__A (.DIODE(\core_1.execute.alu_mul_div.div_cur[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4430__A (.DIODE(\core_1.execute.alu_mul_div.div_cur[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5529__A1 (.DIODE(\core_1.execute.alu_mul_div.div_cur[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4564__A1 (.DIODE(\core_1.execute.alu_mul_div.div_cur[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4559__A1 (.DIODE(\core_1.execute.alu_mul_div.div_cur[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4471__A (.DIODE(\core_1.execute.alu_mul_div.div_cur[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4425__A (.DIODE(\core_1.execute.alu_mul_div.div_cur[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5750__B1 (.DIODE(\core_1.execute.alu_mul_div.i_div ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5719__B1 (.DIODE(\core_1.execute.alu_mul_div.i_div ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5600__B1 (.DIODE(\core_1.execute.alu_mul_div.i_div ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5506__B1 (.DIODE(\core_1.execute.alu_mul_div.i_div ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5468__B1 (.DIODE(\core_1.execute.alu_mul_div.i_div ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5433__B1 (.DIODE(\core_1.execute.alu_mul_div.i_div ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5385__B1 (.DIODE(\core_1.execute.alu_mul_div.i_div ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5250__B1 (.DIODE(\core_1.execute.alu_mul_div.i_div ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3888__A (.DIODE(\core_1.execute.alu_mul_div.i_div ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3593__A (.DIODE(\core_1.execute.alu_mul_div.i_div ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5753__A2 (.DIODE(\core_1.execute.alu_mul_div.i_mod ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5722__A2_N (.DIODE(\core_1.execute.alu_mul_div.i_mod ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5602__A2 (.DIODE(\core_1.execute.alu_mul_div.i_mod ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5570__A2 (.DIODE(\core_1.execute.alu_mul_div.i_mod ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5322__A2 (.DIODE(\core_1.execute.alu_mul_div.i_mod ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5218__B1 (.DIODE(\core_1.execute.alu_mul_div.i_mod ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4781__A (.DIODE(\core_1.execute.alu_mul_div.i_mod ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3856__A (.DIODE(\core_1.execute.alu_mul_div.i_mod ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3593__B (.DIODE(\core_1.execute.alu_mul_div.i_mod ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6312__A1 (.DIODE(\core_1.execute.alu_mul_div.mul_res[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6308__B1 (.DIODE(\core_1.execute.alu_mul_div.mul_res[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6307__A (.DIODE(\core_1.execute.alu_mul_div.mul_res[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5627__A2 (.DIODE(\core_1.execute.alu_mul_div.mul_res[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6219__A1 (.DIODE(\core_1.execute.alu_mul_div.mul_res[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6211__A (.DIODE(\core_1.execute.alu_mul_div.mul_res[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5359__A2 (.DIODE(\core_1.execute.alu_mul_div.mul_res[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6232__A1 (.DIODE(\core_1.execute.alu_mul_div.mul_res[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6226__B1 (.DIODE(\core_1.execute.alu_mul_div.mul_res[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6225__B (.DIODE(\core_1.execute.alu_mul_div.mul_res[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5385__A2 (.DIODE(\core_1.execute.alu_mul_div.mul_res[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6275__A1 (.DIODE(\core_1.execute.alu_mul_div.mul_res[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6270__A (.DIODE(\core_1.execute.alu_mul_div.mul_res[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6269__A (.DIODE(\core_1.execute.alu_mul_div.mul_res[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5528__A2 (.DIODE(\core_1.execute.alu_mul_div.mul_res[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6698__A1 (.DIODE(\core_1.execute.irq_en ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6692__A1 (.DIODE(\core_1.execute.irq_en ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6159__B1 (.DIODE(\core_1.execute.irq_en ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5287__B2 (.DIODE(\core_1.execute.irq_en ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3528__B1 (.DIODE(\core_1.execute.irq_en ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6627__A1 (.DIODE(\core_1.execute.mem_stage_pc[14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4958__A1 (.DIODE(\core_1.execute.mem_stage_pc[14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6762__A1 (.DIODE(\core_1.execute.pc_high_buff_out[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6708__A1 (.DIODE(\core_1.execute.pc_high_buff_out[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5208__A1 (.DIODE(\core_1.execute.pc_high_buff_out[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6765__A1 (.DIODE(\core_1.execute.pc_high_buff_out[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6715__A1 (.DIODE(\core_1.execute.pc_high_buff_out[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5265__A1 (.DIODE(\core_1.execute.pc_high_buff_out[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6771__A1 (.DIODE(\core_1.execute.pc_high_buff_out[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6727__A1 (.DIODE(\core_1.execute.pc_high_buff_out[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5329__B2 (.DIODE(\core_1.execute.pc_high_buff_out[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6774__A1 (.DIODE(\core_1.execute.pc_high_buff_out[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6732__A1 (.DIODE(\core_1.execute.pc_high_buff_out[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5390__B2 (.DIODE(\core_1.execute.pc_high_buff_out[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6780__A1 (.DIODE(\core_1.execute.pc_high_buff_out[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6745__A1 (.DIODE(\core_1.execute.pc_high_buff_out[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5442__B2 (.DIODE(\core_1.execute.pc_high_buff_out[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6748__A (.DIODE(\core_1.execute.pc_high_buff_out[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5480__B2 (.DIODE(\core_1.execute.pc_high_buff_out[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6725__A3 (.DIODE(\core_1.execute.pc_high_out[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6724__D (.DIODE(\core_1.execute.pc_high_out[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6714__A2 (.DIODE(\core_1.execute.pc_high_out[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6713__B (.DIODE(\core_1.execute.pc_high_out[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6712__A1 (.DIODE(\core_1.execute.pc_high_out[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6706__A (.DIODE(\core_1.execute.pc_high_out[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5211__A (.DIODE(\core_1.execute.pc_high_out[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3546__A (.DIODE(\core_1.execute.pc_high_out[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6725__A2 (.DIODE(\core_1.execute.pc_high_out[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6724__C (.DIODE(\core_1.execute.pc_high_out[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6717__A (.DIODE(\core_1.execute.pc_high_out[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6714__A1 (.DIODE(\core_1.execute.pc_high_out[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6713__A (.DIODE(\core_1.execute.pc_high_out[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5270__B2 (.DIODE(\core_1.execute.pc_high_out[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3544__A (.DIODE(\core_1.execute.pc_high_out[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6725__A1 (.DIODE(\core_1.execute.pc_high_out[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6724__B (.DIODE(\core_1.execute.pc_high_out[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6723__A1 (.DIODE(\core_1.execute.pc_high_out[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6719__A (.DIODE(\core_1.execute.pc_high_out[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5284__A1 (.DIODE(\core_1.execute.pc_high_out[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3533__A (.DIODE(\core_1.execute.pc_high_out[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6729__A1 (.DIODE(\core_1.execute.pc_high_out[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6725__B1 (.DIODE(\core_1.execute.pc_high_out[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6724__A (.DIODE(\core_1.execute.pc_high_out[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5331__B2 (.DIODE(\core_1.execute.pc_high_out[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3535__A (.DIODE(\core_1.execute.pc_high_out[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6737__A1 (.DIODE(\core_1.execute.pc_high_out[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6736__B (.DIODE(\core_1.execute.pc_high_out[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6735__A1 (.DIODE(\core_1.execute.pc_high_out[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6731__A1 (.DIODE(\core_1.execute.pc_high_out[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6730__A (.DIODE(\core_1.execute.pc_high_out[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5393__B2 (.DIODE(\core_1.execute.pc_high_out[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3539__A (.DIODE(\core_1.execute.pc_high_out[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6741__A1 (.DIODE(\core_1.execute.pc_high_out[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6737__B1 (.DIODE(\core_1.execute.pc_high_out[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6736__A (.DIODE(\core_1.execute.pc_high_out[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5405__A1 (.DIODE(\core_1.execute.pc_high_out[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3542__A (.DIODE(\core_1.execute.pc_high_out[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6747__A1 (.DIODE(\core_1.execute.pc_high_out[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6743__A (.DIODE(\core_1.execute.pc_high_out[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6742__A (.DIODE(\core_1.execute.pc_high_out[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5444__B2 (.DIODE(\core_1.execute.pc_high_out[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3538__A (.DIODE(\core_1.execute.pc_high_out[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6753__A1 (.DIODE(\core_1.execute.pc_high_out[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6749__A (.DIODE(\core_1.execute.pc_high_out[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5478__A1 (.DIODE(\core_1.execute.pc_high_out[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3534__A (.DIODE(\core_1.execute.pc_high_out[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6112__A1 (.DIODE(\core_1.execute.rf.reg_outputs[1][11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4680__A1 (.DIODE(\core_1.execute.rf.reg_outputs[1][11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3429__D (.DIODE(\core_1.execute.rf.reg_outputs[1][11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6093__A (.DIODE(\core_1.execute.rf.reg_outputs[1][3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5163__A1 (.DIODE(\core_1.execute.rf.reg_outputs[1][3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4735__A1 (.DIODE(\core_1.execute.rf.reg_outputs[1][3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3492__B2 (.DIODE(\core_1.execute.rf.reg_outputs[1][3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6095__A (.DIODE(\core_1.execute.rf.reg_outputs[1][4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5167__A1 (.DIODE(\core_1.execute.rf.reg_outputs[1][4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4740__A1 (.DIODE(\core_1.execute.rf.reg_outputs[1][4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3485__A1 (.DIODE(\core_1.execute.rf.reg_outputs[1][4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6100__A (.DIODE(\core_1.execute.rf.reg_outputs[1][6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5179__A1 (.DIODE(\core_1.execute.rf.reg_outputs[1][6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4747__A1 (.DIODE(\core_1.execute.rf.reg_outputs[1][6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3469__B2 (.DIODE(\core_1.execute.rf.reg_outputs[1][6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6079__A1 (.DIODE(\core_1.execute.rf.reg_outputs[2][13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4694__A1 (.DIODE(\core_1.execute.rf.reg_outputs[2][13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3417__A1 (.DIODE(\core_1.execute.rf.reg_outputs[2][13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6041__A1 (.DIODE(\core_1.execute.rf.reg_outputs[3][13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4693__B2 (.DIODE(\core_1.execute.rf.reg_outputs[3][13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3413__D (.DIODE(\core_1.execute.rf.reg_outputs[3][13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6033__A1 (.DIODE(\core_1.execute.rf.reg_outputs[3][9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4625__A (.DIODE(\core_1.execute.rf.reg_outputs[3][9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3448__D (.DIODE(\core_1.execute.rf.reg_outputs[3][9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5999__A1 (.DIODE(\core_1.execute.rf.reg_outputs[4][11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4679__A (.DIODE(\core_1.execute.rf.reg_outputs[4][11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3430__A1 (.DIODE(\core_1.execute.rf.reg_outputs[4][11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6008__A1 (.DIODE(\core_1.execute.rf.reg_outputs[4][15] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4615__A1 (.DIODE(\core_1.execute.rf.reg_outputs[4][15] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3380__A (.DIODE(\core_1.execute.rf.reg_outputs[4][15] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5993__A1 (.DIODE(\core_1.execute.rf.reg_outputs[4][8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4655__A (.DIODE(\core_1.execute.rf.reg_outputs[4][8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3454__B2 (.DIODE(\core_1.execute.rf.reg_outputs[4][8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5995__A1 (.DIODE(\core_1.execute.rf.reg_outputs[4][9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4627__A (.DIODE(\core_1.execute.rf.reg_outputs[4][9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3445__B2 (.DIODE(\core_1.execute.rf.reg_outputs[4][9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5937__A (.DIODE(\core_1.execute.rf.reg_outputs[5][0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4723__C (.DIODE(\core_1.execute.rf.reg_outputs[5][0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3518__C (.DIODE(\core_1.execute.rf.reg_outputs[5][0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5962__A1 (.DIODE(\core_1.execute.rf.reg_outputs[5][11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4678__A1 (.DIODE(\core_1.execute.rf.reg_outputs[5][11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3427__C (.DIODE(\core_1.execute.rf.reg_outputs[5][11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5966__A1 (.DIODE(\core_1.execute.rf.reg_outputs[5][13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4691__A1 (.DIODE(\core_1.execute.rf.reg_outputs[5][13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3412__A1 (.DIODE(\core_1.execute.rf.reg_outputs[5][13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5968__A1 (.DIODE(\core_1.execute.rf.reg_outputs[5][14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4687__A1 (.DIODE(\core_1.execute.rf.reg_outputs[5][14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3393__C (.DIODE(\core_1.execute.rf.reg_outputs[5][14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5958__A1 (.DIODE(\core_1.execute.rf.reg_outputs[5][9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4626__A1 (.DIODE(\core_1.execute.rf.reg_outputs[5][9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3445__A1 (.DIODE(\core_1.execute.rf.reg_outputs[5][9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5923__A1 (.DIODE(\core_1.execute.rf.reg_outputs[6][11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4677__A1 (.DIODE(\core_1.execute.rf.reg_outputs[6][11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3428__D (.DIODE(\core_1.execute.rf.reg_outputs[6][11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5925__A1 (.DIODE(\core_1.execute.rf.reg_outputs[6][12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4673__B2 (.DIODE(\core_1.execute.rf.reg_outputs[6][12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3420__B2 (.DIODE(\core_1.execute.rf.reg_outputs[6][12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5927__A1 (.DIODE(\core_1.execute.rf.reg_outputs[6][13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4691__B2 (.DIODE(\core_1.execute.rf.reg_outputs[6][13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3407__B2 (.DIODE(\core_1.execute.rf.reg_outputs[6][13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5917__A1 (.DIODE(\core_1.execute.rf.reg_outputs[6][8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4656__A1 (.DIODE(\core_1.execute.rf.reg_outputs[6][8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3453__B2 (.DIODE(\core_1.execute.rf.reg_outputs[6][8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5919__A1 (.DIODE(\core_1.execute.rf.reg_outputs[6][9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4629__B2 (.DIODE(\core_1.execute.rf.reg_outputs[6][9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3446__B2 (.DIODE(\core_1.execute.rf.reg_outputs[6][9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5886__A1 (.DIODE(\core_1.execute.rf.reg_outputs[7][13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4695__A1 (.DIODE(\core_1.execute.rf.reg_outputs[7][13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3414__A (.DIODE(\core_1.execute.rf.reg_outputs[7][13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6696__A1 (.DIODE(\core_1.execute.sreg_irq_flags.i_d[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3529__B (.DIODE(\core_1.execute.sreg_irq_flags.i_d[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6692__B2 (.DIODE(\core_1.execute.sreg_irq_flags.o_d[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5200__A (.DIODE(\core_1.execute.sreg_irq_flags.o_d[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6693__A (.DIODE(\core_1.execute.sreg_irq_flags.o_d[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5264__A (.DIODE(\core_1.execute.sreg_irq_flags.o_d[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6698__B2 (.DIODE(\core_1.execute.sreg_irq_flags.o_d[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5392__A (.DIODE(\core_1.execute.sreg_irq_flags.o_d[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6568__A1 (.DIODE(\core_1.execute.sreg_irq_pc.o_d[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5201__A1 (.DIODE(\core_1.execute.sreg_irq_pc.o_d[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5191__A (.DIODE(\core_1.execute.sreg_irq_pc.o_d[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6572__A1 (.DIODE(\core_1.execute.sreg_irq_pc.o_d[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5267__A1 (.DIODE(\core_1.execute.sreg_irq_pc.o_d[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4898__A (.DIODE(\core_1.execute.sreg_irq_pc.o_d[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6581__A1 (.DIODE(\core_1.execute.sreg_irq_pc.o_d[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6422__A (.DIODE(\core_1.execute.sreg_irq_pc.o_d[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5290__A1 (.DIODE(\core_1.execute.sreg_irq_pc.o_d[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5283__A1 (.DIODE(\core_1.execute.sreg_irq_pc.o_d[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6589__A1 (.DIODE(\core_1.execute.sreg_irq_pc.o_d[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6435__A1 (.DIODE(\core_1.execute.sreg_irq_pc.o_d[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5396__A0 (.DIODE(\core_1.execute.sreg_irq_pc.o_d[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5390__A1 (.DIODE(\core_1.execute.sreg_irq_pc.o_d[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6593__A1 (.DIODE(\core_1.execute.sreg_irq_pc.o_d[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6440__A1 (.DIODE(\core_1.execute.sreg_irq_pc.o_d[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5409__A (.DIODE(\core_1.execute.sreg_irq_pc.o_d[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5406__A1 (.DIODE(\core_1.execute.sreg_irq_pc.o_d[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6601__A1 (.DIODE(\core_1.execute.sreg_irq_pc.o_d[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5482__A (.DIODE(\core_1.execute.sreg_irq_pc.o_d[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5478__B2 (.DIODE(\core_1.execute.sreg_irq_pc.o_d[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5811__A (.DIODE(\core_1.execute.sreg_long_ptr_en ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5328__A1 (.DIODE(\core_1.execute.sreg_long_ptr_en ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4150__B2 (.DIODE(\core_1.execute.sreg_long_ptr_en ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3579__B1 (.DIODE(\core_1.execute.sreg_long_ptr_en ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6649__B2 (.DIODE(\core_1.execute.trap_flag ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5267__B2 (.DIODE(\core_1.execute.trap_flag ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4969__A (.DIODE(\core_1.execute.trap_flag ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3632__B_N (.DIODE(\core_1.fetch.out_buffer_valid ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3627__B_N (.DIODE(\core_1.fetch.out_buffer_valid ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3625__B_N (.DIODE(\core_1.fetch.out_buffer_valid ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3624__S (.DIODE(\core_1.fetch.out_buffer_valid ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3623__S (.DIODE(\core_1.fetch.out_buffer_valid ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3621__S (.DIODE(\core_1.fetch.out_buffer_valid ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3618__B_N (.DIODE(\core_1.fetch.out_buffer_valid ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3613__A (.DIODE(\core_1.fetch.out_buffer_valid ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3610__S (.DIODE(\core_1.fetch.out_buffer_valid ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3525__A (.DIODE(\core_1.fetch.out_buffer_valid ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4280__C_N (.DIODE(\core_1.fetch.prev_request_pc[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3778__B1 (.DIODE(\core_1.fetch.prev_request_pc[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3715__A (.DIODE(\core_1.fetch.prev_request_pc[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3688__B2 (.DIODE(\core_1.fetch.prev_request_pc[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3677__A (.DIODE(\core_1.fetch.prev_request_pc[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4282__A (.DIODE(\core_1.fetch.prev_request_pc[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3774__A (.DIODE(\core_1.fetch.prev_request_pc[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3716__A (.DIODE(\core_1.fetch.prev_request_pc[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3688__A1 (.DIODE(\core_1.fetch.prev_request_pc[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3685__A1_N (.DIODE(\core_1.fetch.prev_request_pc[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4296__B2 (.DIODE(\core_1.fetch.prev_request_pc[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3753__A (.DIODE(\core_1.fetch.prev_request_pc[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3748__A (.DIODE(\core_1.fetch.prev_request_pc[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3719__B (.DIODE(\core_1.fetch.prev_request_pc[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3663__A1 (.DIODE(\core_1.fetch.prev_request_pc[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3652__B2 (.DIODE(\core_1.fetch.prev_request_pc[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4297__B2 (.DIODE(\core_1.fetch.prev_request_pc[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3749__A (.DIODE(\core_1.fetch.prev_request_pc[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3719__A (.DIODE(\core_1.fetch.prev_request_pc[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3655__A1_N (.DIODE(\core_1.fetch.prev_request_pc[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3652__A1 (.DIODE(\core_1.fetch.prev_request_pc[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_i_clk_A (.DIODE(i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_input1_A (.DIODE(i_core_int_sreg[0]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input2_A (.DIODE(i_core_int_sreg[10]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input3_A (.DIODE(i_core_int_sreg[11]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input4_A (.DIODE(i_core_int_sreg[12]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input5_A (.DIODE(i_core_int_sreg[13]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input6_A (.DIODE(i_core_int_sreg[14]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input7_A (.DIODE(i_core_int_sreg[15]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input8_A (.DIODE(i_core_int_sreg[1]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input9_A (.DIODE(i_core_int_sreg[2]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input10_A (.DIODE(i_core_int_sreg[3]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input11_A (.DIODE(i_core_int_sreg[4]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input12_A (.DIODE(i_core_int_sreg[5]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input13_A (.DIODE(i_core_int_sreg[6]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input14_A (.DIODE(i_core_int_sreg[7]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input15_A (.DIODE(i_core_int_sreg[8]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input16_A (.DIODE(i_core_int_sreg[9]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input17_A (.DIODE(i_disable));
 sky130_fd_sc_hd__diode_2 ANTENNA_input18_A (.DIODE(i_irq));
 sky130_fd_sc_hd__diode_2 ANTENNA_input19_A (.DIODE(i_mc_core_int));
 sky130_fd_sc_hd__diode_2 ANTENNA_input20_A (.DIODE(i_mem_ack));
 sky130_fd_sc_hd__diode_2 ANTENNA_input21_A (.DIODE(i_mem_data[0]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input22_A (.DIODE(i_mem_data[10]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input23_A (.DIODE(i_mem_data[11]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input24_A (.DIODE(i_mem_data[12]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input25_A (.DIODE(i_mem_data[13]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input26_A (.DIODE(i_mem_data[14]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input27_A (.DIODE(i_mem_data[15]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input28_A (.DIODE(i_mem_data[1]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input29_A (.DIODE(i_mem_data[2]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input30_A (.DIODE(i_mem_data[3]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input31_A (.DIODE(i_mem_data[4]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input32_A (.DIODE(i_mem_data[5]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input33_A (.DIODE(i_mem_data[6]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input34_A (.DIODE(i_mem_data[7]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input35_A (.DIODE(i_mem_data[8]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input36_A (.DIODE(i_mem_data[9]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input37_A (.DIODE(i_mem_exception));
 sky130_fd_sc_hd__diode_2 ANTENNA_input38_A (.DIODE(i_req_data[0]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input39_A (.DIODE(i_req_data[10]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input40_A (.DIODE(i_req_data[11]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input41_A (.DIODE(i_req_data[12]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input42_A (.DIODE(i_req_data[13]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input43_A (.DIODE(i_req_data[14]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input44_A (.DIODE(i_req_data[15]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input45_A (.DIODE(i_req_data[16]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input46_A (.DIODE(i_req_data[17]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input47_A (.DIODE(i_req_data[18]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input48_A (.DIODE(i_req_data[19]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input49_A (.DIODE(i_req_data[1]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input50_A (.DIODE(i_req_data[20]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input51_A (.DIODE(i_req_data[21]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input52_A (.DIODE(i_req_data[22]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input53_A (.DIODE(i_req_data[23]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input54_A (.DIODE(i_req_data[24]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input55_A (.DIODE(i_req_data[25]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input56_A (.DIODE(i_req_data[26]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input57_A (.DIODE(i_req_data[27]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input58_A (.DIODE(i_req_data[28]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input59_A (.DIODE(i_req_data[29]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input60_A (.DIODE(i_req_data[2]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input61_A (.DIODE(i_req_data[30]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input62_A (.DIODE(i_req_data[31]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input63_A (.DIODE(i_req_data[3]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input64_A (.DIODE(i_req_data[4]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input65_A (.DIODE(i_req_data[5]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input66_A (.DIODE(i_req_data[6]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input67_A (.DIODE(i_req_data[7]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input68_A (.DIODE(i_req_data[8]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input69_A (.DIODE(i_req_data[9]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input70_A (.DIODE(i_req_data_valid));
 sky130_fd_sc_hd__diode_2 ANTENNA_input71_A (.DIODE(i_rst));
 sky130_fd_sc_hd__diode_2 ANTENNA__7188__CLK (.DIODE(clknet_leaf_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6972__CLK (.DIODE(clknet_leaf_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7190__CLK (.DIODE(clknet_leaf_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__5699__B2 (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 ANTENNA__5729__B2 (.DIODE(net7));
 sky130_fd_sc_hd__diode_2 ANTENNA__5405__B2 (.DIODE(net12));
 sky130_fd_sc_hd__diode_2 ANTENNA__5479__B2 (.DIODE(net14));
 sky130_fd_sc_hd__diode_2 ANTENNA__5814__A1 (.DIODE(net20));
 sky130_fd_sc_hd__diode_2 ANTENNA__3591__A (.DIODE(net20));
 sky130_fd_sc_hd__diode_2 ANTENNA__5817__A1 (.DIODE(net21));
 sky130_fd_sc_hd__diode_2 ANTENNA__5875__A1_N (.DIODE(net23));
 sky130_fd_sc_hd__diode_2 ANTENNA__5835__A0 (.DIODE(net23));
 sky130_fd_sc_hd__diode_2 ANTENNA__5880__A1_N (.DIODE(net24));
 sky130_fd_sc_hd__diode_2 ANTENNA__5840__A0 (.DIODE(net24));
 sky130_fd_sc_hd__diode_2 ANTENNA__5884__A1_N (.DIODE(net25));
 sky130_fd_sc_hd__diode_2 ANTENNA__5845__A0 (.DIODE(net25));
 sky130_fd_sc_hd__diode_2 ANTENNA__5888__A1_N (.DIODE(net26));
 sky130_fd_sc_hd__diode_2 ANTENNA__5850__A0 (.DIODE(net26));
 sky130_fd_sc_hd__diode_2 ANTENNA__5892__A1_N (.DIODE(net27));
 sky130_fd_sc_hd__diode_2 ANTENNA__5855__A0 (.DIODE(net27));
 sky130_fd_sc_hd__diode_2 ANTENNA__5824__A1 (.DIODE(net28));
 sky130_fd_sc_hd__diode_2 ANTENNA__5830__A1 (.DIODE(net29));
 sky130_fd_sc_hd__diode_2 ANTENNA__5835__A1 (.DIODE(net30));
 sky130_fd_sc_hd__diode_2 ANTENNA__5840__A1 (.DIODE(net31));
 sky130_fd_sc_hd__diode_2 ANTENNA__5845__A1 (.DIODE(net32));
 sky130_fd_sc_hd__diode_2 ANTENNA__5850__A1 (.DIODE(net33));
 sky130_fd_sc_hd__diode_2 ANTENNA__5855__A1 (.DIODE(net34));
 sky130_fd_sc_hd__diode_2 ANTENNA__6631__S (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA__6627__S (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA__6623__S (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA__6618__S (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA__6582__S (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA__6574__A (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA__6569__S (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA__6564__S (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA__4386__A (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA__3529__A (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA__4225__A0 (.DIODE(net69));
 sky130_fd_sc_hd__diode_2 ANTENNA__3704__A0 (.DIODE(net69));
 sky130_fd_sc_hd__diode_2 ANTENNA__4378__B (.DIODE(net70));
 sky130_fd_sc_hd__diode_2 ANTENNA__4273__A1 (.DIODE(net70));
 sky130_fd_sc_hd__diode_2 ANTENNA__4204__D_N (.DIODE(net70));
 sky130_fd_sc_hd__diode_2 ANTENNA__3947__A2 (.DIODE(net70));
 sky130_fd_sc_hd__diode_2 ANTENNA__3906__S (.DIODE(net70));
 sky130_fd_sc_hd__diode_2 ANTENNA__3642__A2 (.DIODE(net70));
 sky130_fd_sc_hd__diode_2 ANTENNA__6415__A (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA__4902__B (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA__4295__A (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA__4204__A (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA__4201__B (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA__4144__A (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA__4056__A (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA__3802__A (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA__3799__A (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA__3523__A (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA_output73_A (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA__6610__A0 (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA__6489__C (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA__6470__A (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA__6469__B1 (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA__5578__A1 (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA__4949__A (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA__3747__A1 (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA_output74_A (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA__6614__A0 (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA__6489__B (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA__6477__A (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA__6476__A (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA__5632__A1 (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA__4951__A (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA__3744__A1 (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA_output75_A (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA__6618__A0 (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA__6489__A (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA__6485__A1 (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA__6484__A1 (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA__5641__A1 (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA__4953__A (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA__3740__A1 (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA_output76_A (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA__6623__A0 (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA__6497__A (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA__6492__A (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA__5671__A1 (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA__4955__A (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA__3736__A1 (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA_output77_A (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA__6701__A2 (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA__6627__A0 (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA__6499__A (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA__6498__A (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA__5701__A1 (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA__4957__A (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA__3733__A1 (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA_output78_A (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA__6631__A0 (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA__6503__A (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA__5731__A1 (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA__4959__A (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA__3729__A1 (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA_output79_A (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA__6569__A0 (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA__6419__C (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA__6418__A2 (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA__5262__A (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA__4925__A (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA__4778__B (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA__4771__B1 (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA__3785__A1 (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA_output80_A (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA__6575__A0 (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA__6419__A (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA__6418__B1 (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA__5281__A1 (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA__4927__A (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA__3781__A1 (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA_output81_A (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA__6582__A0 (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA__6441__B (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA__5333__A1 (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA__4929__A (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA__3777__A1 (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA_output82_A (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA__6586__A0 (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA__6443__B (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA__6441__A (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA__5395__A1 (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA__4933__A (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA__3773__A1 (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA_output83_A (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA__6590__A0 (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA__6496__A (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA__6490__A (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA__6443__A (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA__6442__B1 (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA__5408__A1 (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA__4936__A (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA__3769__A1 (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA_output84_A (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA__6594__A0 (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA__6488__C (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA__6453__B (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA__6452__A1 (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA__6448__A (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA__5445__A1 (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA__4938__A (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA__3765__A1 (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA_output85_A (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA__6598__A0 (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA__6488__B (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA__6453__A (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA__6452__B1 (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA__5481__A1 (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA__4941__A (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA__3761__A1 (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA_output86_A (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA__6602__A0 (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA__6488__A (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA__6457__A (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA__6456__A (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA__5533__A1 (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA__4945__A (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA__3756__A1 (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA_output87_A (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA__6606__A0 (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA__6489__D (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA__6470__B (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA__6469__A1 (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA__6463__A (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA__5544__A1 (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA__4947__A (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA__3752__A1 (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA_output88_A (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA__6125__A (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA__4729__A (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA__3520__A (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA_output89_A (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA__6148__A1 (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA__4637__A1 (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA__4418__A1 (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA__3443__A1 (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA_output90_A (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA__6150__A1 (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA__4681__B2 (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA__4414__A1 (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA__3434__A1 (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA_output91_A (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA__6152__A1 (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA__4674__A1 (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA__3425__B2 (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA_output92_A (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA__6154__A1 (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA__4696__A1 (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA__3418__B2 (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA_output93_A (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA__6156__A1 (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA__4688__A1 (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA__4401__A1 (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA__3402__A1 (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA_output94_A (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA__6158__A1 (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA__4791__A1 (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA__4624__A1 (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA__4396__A1 (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA__3390__A1 (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA_output95_A (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA__6127__A (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA__4713__A (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA__3512__A (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA_output96_A (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA__6129__A (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA__4711__A (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA__3505__A1 (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA_output97_A (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 ANTENNA__6131__A (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 ANTENNA__4819__A1 (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 ANTENNA__4738__A1 (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 ANTENNA__3496__B2 (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 ANTENNA_output98_A (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA__6133__A (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA__4820__A1 (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA__4745__A1 (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA__3489__B2 (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA_output99_A (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 ANTENNA__6135__A (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 ANTENNA__4759__B2 (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 ANTENNA__3482__B2 (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 ANTENNA_output100_A (.DIODE(net100));
 sky130_fd_sc_hd__diode_2 ANTENNA__6137__A (.DIODE(net100));
 sky130_fd_sc_hd__diode_2 ANTENNA__4751__A1 (.DIODE(net100));
 sky130_fd_sc_hd__diode_2 ANTENNA__3474__A (.DIODE(net100));
 sky130_fd_sc_hd__diode_2 ANTENNA_output101_A (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA__6139__A (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA__4651__A1 (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA__3466__A (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA_output102_A (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA__6143__A1 (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA__4658__A1 (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA__3458__B2 (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA_output103_A (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA__6146__A1 (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA__4630__A1 (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA__3450__A (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA_output104_A (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA__4917__A1 (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA_output106_A (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA__6647__A (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA__5210__A (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA__3988__A1 (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA__3987__A (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA_output109_A (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 ANTENNA_output110_A (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA_output111_A (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA_output112_A (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA_output115_A (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA_output132_A (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA__5148__A0 (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA_output133_A (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 ANTENNA__5160__A1 (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 ANTENNA_output134_A (.DIODE(net134));
 sky130_fd_sc_hd__diode_2 ANTENNA__5165__A0 (.DIODE(net134));
 sky130_fd_sc_hd__diode_2 ANTENNA_output135_A (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA__5172__A0 (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA_output136_A (.DIODE(net136));
 sky130_fd_sc_hd__diode_2 ANTENNA__5177__A0 (.DIODE(net136));
 sky130_fd_sc_hd__diode_2 ANTENNA_output137_A (.DIODE(net137));
 sky130_fd_sc_hd__diode_2 ANTENNA__5183__A0 (.DIODE(net137));
 sky130_fd_sc_hd__diode_2 ANTENNA_output138_A (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA__5189__A (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA_output155_A (.DIODE(net155));
 sky130_fd_sc_hd__diode_2 ANTENNA__5812__A1 (.DIODE(net155));
 sky130_fd_sc_hd__diode_2 ANTENNA__3949__A (.DIODE(net155));
 sky130_fd_sc_hd__diode_2 ANTENNA_output156_A (.DIODE(net156));
 sky130_fd_sc_hd__diode_2 ANTENNA__3592__A1 (.DIODE(net156));
 sky130_fd_sc_hd__diode_2 ANTENNA_output157_A (.DIODE(net157));
 sky130_fd_sc_hd__diode_2 ANTENNA__3927__S (.DIODE(net157));
 sky130_fd_sc_hd__diode_2 ANTENNA__3925__B (.DIODE(net157));
 sky130_fd_sc_hd__diode_2 ANTENNA__3923__B (.DIODE(net157));
 sky130_fd_sc_hd__diode_2 ANTENNA__3921__B (.DIODE(net157));
 sky130_fd_sc_hd__diode_2 ANTENNA__3919__B (.DIODE(net157));
 sky130_fd_sc_hd__diode_2 ANTENNA__3917__B (.DIODE(net157));
 sky130_fd_sc_hd__diode_2 ANTENNA__3915__B (.DIODE(net157));
 sky130_fd_sc_hd__diode_2 ANTENNA__3913__B (.DIODE(net157));
 sky130_fd_sc_hd__diode_2 ANTENNA__3911__B (.DIODE(net157));
 sky130_fd_sc_hd__diode_2 ANTENNA_output161_A (.DIODE(net161));
 sky130_fd_sc_hd__diode_2 ANTENNA__4276__A1 (.DIODE(net161));
 sky130_fd_sc_hd__diode_2 ANTENNA_output162_A (.DIODE(net162));
 sky130_fd_sc_hd__diode_2 ANTENNA__4298__A2 (.DIODE(net162));
 sky130_fd_sc_hd__diode_2 ANTENNA_output168_A (.DIODE(net168));
 sky130_fd_sc_hd__diode_2 ANTENNA__4279__A2 (.DIODE(net168));
 sky130_fd_sc_hd__diode_2 ANTENNA_output169_A (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 ANTENNA__4281__A2 (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 ANTENNA_output170_A (.DIODE(net170));
 sky130_fd_sc_hd__diode_2 ANTENNA__4283__A1 (.DIODE(net170));
 sky130_fd_sc_hd__diode_2 ANTENNA_output171_A (.DIODE(net171));
 sky130_fd_sc_hd__diode_2 ANTENNA__4286__A2 (.DIODE(net171));
 sky130_fd_sc_hd__diode_2 ANTENNA_output172_A (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 ANTENNA__4288__A2 (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 ANTENNA_output173_A (.DIODE(net173));
 sky130_fd_sc_hd__diode_2 ANTENNA__4290__A1 (.DIODE(net173));
 sky130_fd_sc_hd__diode_2 ANTENNA_output174_A (.DIODE(net174));
 sky130_fd_sc_hd__diode_2 ANTENNA__4293__A1 (.DIODE(net174));
 sky130_fd_sc_hd__diode_2 ANTENNA_output175_A (.DIODE(net175));
 sky130_fd_sc_hd__diode_2 ANTENNA__4296__A2 (.DIODE(net175));
 sky130_fd_sc_hd__diode_2 ANTENNA_output176_A (.DIODE(net176));
 sky130_fd_sc_hd__diode_2 ANTENNA__4297__A2 (.DIODE(net176));
 sky130_fd_sc_hd__diode_2 ANTENNA_output177_A (.DIODE(net177));
 sky130_fd_sc_hd__diode_2 ANTENNA__4379__B1 (.DIODE(net177));
 sky130_fd_sc_hd__diode_2 ANTENNA__4299__A1 (.DIODE(net177));
 sky130_fd_sc_hd__diode_2 ANTENNA__4298__A1 (.DIODE(net177));
 sky130_fd_sc_hd__diode_2 ANTENNA__4297__A1 (.DIODE(net177));
 sky130_fd_sc_hd__diode_2 ANTENNA__4296__A1 (.DIODE(net177));
 sky130_fd_sc_hd__diode_2 ANTENNA__4288__A1 (.DIODE(net177));
 sky130_fd_sc_hd__diode_2 ANTENNA__4286__A1 (.DIODE(net177));
 sky130_fd_sc_hd__diode_2 ANTENNA__4281__A1 (.DIODE(net177));
 sky130_fd_sc_hd__diode_2 ANTENNA__4279__A1 (.DIODE(net177));
 sky130_fd_sc_hd__diode_2 ANTENNA_output178_A (.DIODE(net178));
 sky130_fd_sc_hd__diode_2 ANTENNA__5198__A_N (.DIODE(net178));
 sky130_fd_sc_hd__diode_2 ANTENNA__5194__B (.DIODE(net178));
 sky130_fd_sc_hd__diode_2 ANTENNA__4457__B (.DIODE(net178));
 sky130_fd_sc_hd__diode_2 ANTENNA__4135__B (.DIODE(net178));
 sky130_fd_sc_hd__diode_2 ANTENNA__4077__A0 (.DIODE(net178));
 sky130_fd_sc_hd__diode_2 ANTENNA__3977__B_N (.DIODE(net178));
 sky130_fd_sc_hd__diode_2 ANTENNA_output179_A (.DIODE(net179));
 sky130_fd_sc_hd__diode_2 ANTENNA__4417__B (.DIODE(net179));
 sky130_fd_sc_hd__diode_2 ANTENNA__4098__A0 (.DIODE(net179));
 sky130_fd_sc_hd__diode_2 ANTENNA__3982__B (.DIODE(net179));
 sky130_fd_sc_hd__diode_2 ANTENNA__3976__D (.DIODE(net179));
 sky130_fd_sc_hd__diode_2 ANTENNA_output180_A (.DIODE(net180));
 sky130_fd_sc_hd__diode_2 ANTENNA__4995__A2 (.DIODE(net180));
 sky130_fd_sc_hd__diode_2 ANTENNA__4797__A2 (.DIODE(net180));
 sky130_fd_sc_hd__diode_2 ANTENNA__4415__A2 (.DIODE(net180));
 sky130_fd_sc_hd__diode_2 ANTENNA__4100__A0 (.DIODE(net180));
 sky130_fd_sc_hd__diode_2 ANTENNA__3982__A (.DIODE(net180));
 sky130_fd_sc_hd__diode_2 ANTENNA__3976__C (.DIODE(net180));
 sky130_fd_sc_hd__diode_2 ANTENNA_output181_A (.DIODE(net181));
 sky130_fd_sc_hd__diode_2 ANTENNA__4408__B (.DIODE(net181));
 sky130_fd_sc_hd__diode_2 ANTENNA__4102__A0 (.DIODE(net181));
 sky130_fd_sc_hd__diode_2 ANTENNA__3975__B (.DIODE(net181));
 sky130_fd_sc_hd__diode_2 ANTENNA_output182_A (.DIODE(net182));
 sky130_fd_sc_hd__diode_2 ANTENNA__4795__A0 (.DIODE(net182));
 sky130_fd_sc_hd__diode_2 ANTENNA__4405__A (.DIODE(net182));
 sky130_fd_sc_hd__diode_2 ANTENNA__4104__A0 (.DIODE(net182));
 sky130_fd_sc_hd__diode_2 ANTENNA__3975__A (.DIODE(net182));
 sky130_fd_sc_hd__diode_2 ANTENNA_output183_A (.DIODE(net183));
 sky130_fd_sc_hd__diode_2 ANTENNA__4399__B (.DIODE(net183));
 sky130_fd_sc_hd__diode_2 ANTENNA__4106__A0 (.DIODE(net183));
 sky130_fd_sc_hd__diode_2 ANTENNA__3975__D (.DIODE(net183));
 sky130_fd_sc_hd__diode_2 ANTENNA_output184_A (.DIODE(net184));
 sky130_fd_sc_hd__diode_2 ANTENNA__4978__A2 (.DIODE(net184));
 sky130_fd_sc_hd__diode_2 ANTENNA__4796__A2 (.DIODE(net184));
 sky130_fd_sc_hd__diode_2 ANTENNA__4397__A2 (.DIODE(net184));
 sky130_fd_sc_hd__diode_2 ANTENNA__4108__A0 (.DIODE(net184));
 sky130_fd_sc_hd__diode_2 ANTENNA__3975__C (.DIODE(net184));
 sky130_fd_sc_hd__diode_2 ANTENNA_output185_A (.DIODE(net185));
 sky130_fd_sc_hd__diode_2 ANTENNA__5198__D (.DIODE(net185));
 sky130_fd_sc_hd__diode_2 ANTENNA__5194__A (.DIODE(net185));
 sky130_fd_sc_hd__diode_2 ANTENNA__4454__B (.DIODE(net185));
 sky130_fd_sc_hd__diode_2 ANTENNA__4135__A_N (.DIODE(net185));
 sky130_fd_sc_hd__diode_2 ANTENNA__4079__A0 (.DIODE(net185));
 sky130_fd_sc_hd__diode_2 ANTENNA__3977__A_N (.DIODE(net185));
 sky130_fd_sc_hd__diode_2 ANTENNA_output186_A (.DIODE(net186));
 sky130_fd_sc_hd__diode_2 ANTENNA__5202__B (.DIODE(net186));
 sky130_fd_sc_hd__diode_2 ANTENNA__5197__B (.DIODE(net186));
 sky130_fd_sc_hd__diode_2 ANTENNA__4451__A0 (.DIODE(net186));
 sky130_fd_sc_hd__diode_2 ANTENNA__4081__A0 (.DIODE(net186));
 sky130_fd_sc_hd__diode_2 ANTENNA__3972__A (.DIODE(net186));
 sky130_fd_sc_hd__diode_2 ANTENNA_output187_A (.DIODE(net187));
 sky130_fd_sc_hd__diode_2 ANTENNA__5209__A (.DIODE(net187));
 sky130_fd_sc_hd__diode_2 ANTENNA__5206__A (.DIODE(net187));
 sky130_fd_sc_hd__diode_2 ANTENNA__5202__A (.DIODE(net187));
 sky130_fd_sc_hd__diode_2 ANTENNA__5197__A_N (.DIODE(net187));
 sky130_fd_sc_hd__diode_2 ANTENNA__4447__B (.DIODE(net187));
 sky130_fd_sc_hd__diode_2 ANTENNA__4083__A0 (.DIODE(net187));
 sky130_fd_sc_hd__diode_2 ANTENNA__3974__A_N (.DIODE(net187));
 sky130_fd_sc_hd__diode_2 ANTENNA_output188_A (.DIODE(net188));
 sky130_fd_sc_hd__diode_2 ANTENNA__4443__A (.DIODE(net188));
 sky130_fd_sc_hd__diode_2 ANTENNA__4440__A0 (.DIODE(net188));
 sky130_fd_sc_hd__diode_2 ANTENNA__4086__A0 (.DIODE(net188));
 sky130_fd_sc_hd__diode_2 ANTENNA__3973__B (.DIODE(net188));
 sky130_fd_sc_hd__diode_2 ANTENNA_output189_A (.DIODE(net189));
 sky130_fd_sc_hd__diode_2 ANTENNA__4436__B (.DIODE(net189));
 sky130_fd_sc_hd__diode_2 ANTENNA__4088__A0 (.DIODE(net189));
 sky130_fd_sc_hd__diode_2 ANTENNA__3973__A (.DIODE(net189));
 sky130_fd_sc_hd__diode_2 ANTENNA_output190_A (.DIODE(net190));
 sky130_fd_sc_hd__diode_2 ANTENNA__4431__A0 (.DIODE(net190));
 sky130_fd_sc_hd__diode_2 ANTENNA__4090__A0 (.DIODE(net190));
 sky130_fd_sc_hd__diode_2 ANTENNA__3973__D (.DIODE(net190));
 sky130_fd_sc_hd__diode_2 ANTENNA_output191_A (.DIODE(net191));
 sky130_fd_sc_hd__diode_2 ANTENNA__4428__B (.DIODE(net191));
 sky130_fd_sc_hd__diode_2 ANTENNA__4092__A0 (.DIODE(net191));
 sky130_fd_sc_hd__diode_2 ANTENNA__3973__C (.DIODE(net191));
 sky130_fd_sc_hd__diode_2 ANTENNA_output192_A (.DIODE(net192));
 sky130_fd_sc_hd__diode_2 ANTENNA__4426__A0 (.DIODE(net192));
 sky130_fd_sc_hd__diode_2 ANTENNA__4094__A0 (.DIODE(net192));
 sky130_fd_sc_hd__diode_2 ANTENNA__3983__B (.DIODE(net192));
 sky130_fd_sc_hd__diode_2 ANTENNA__3976__B (.DIODE(net192));
 sky130_fd_sc_hd__diode_2 ANTENNA_output193_A (.DIODE(net193));
 sky130_fd_sc_hd__diode_2 ANTENNA__4422__B (.DIODE(net193));
 sky130_fd_sc_hd__diode_2 ANTENNA__4096__A0 (.DIODE(net193));
 sky130_fd_sc_hd__diode_2 ANTENNA__3983__A_N (.DIODE(net193));
 sky130_fd_sc_hd__diode_2 ANTENNA__3976__A (.DIODE(net193));
 sky130_fd_sc_hd__diode_2 ANTENNA_output194_A (.DIODE(net194));
 sky130_fd_sc_hd__diode_2 ANTENNA__6710__A1 (.DIODE(net194));
 sky130_fd_sc_hd__diode_2 ANTENNA__6660__A1 (.DIODE(net194));
 sky130_fd_sc_hd__diode_2 ANTENNA__6637__A1 (.DIODE(net194));
 sky130_fd_sc_hd__diode_2 ANTENNA__6566__A0 (.DIODE(net194));
 sky130_fd_sc_hd__diode_2 ANTENNA__6520__A (.DIODE(net194));
 sky130_fd_sc_hd__diode_2 ANTENNA__6412__A1 (.DIODE(net194));
 sky130_fd_sc_hd__diode_2 ANTENNA__5257__A1 (.DIODE(net194));
 sky130_fd_sc_hd__diode_2 ANTENNA__4145__A1 (.DIODE(net194));
 sky130_fd_sc_hd__diode_2 ANTENNA_output195_A (.DIODE(net195));
 sky130_fd_sc_hd__diode_2 ANTENNA__6681__A1 (.DIODE(net195));
 sky130_fd_sc_hd__diode_2 ANTENNA__6472__A1 (.DIODE(net195));
 sky130_fd_sc_hd__diode_2 ANTENNA__5604__A1 (.DIODE(net195));
 sky130_fd_sc_hd__diode_2 ANTENNA__4172__A1 (.DIODE(net195));
 sky130_fd_sc_hd__diode_2 ANTENNA_output196_A (.DIODE(net196));
 sky130_fd_sc_hd__diode_2 ANTENNA__6683__A1 (.DIODE(net196));
 sky130_fd_sc_hd__diode_2 ANTENNA__6479__B1 (.DIODE(net196));
 sky130_fd_sc_hd__diode_2 ANTENNA__4175__A1 (.DIODE(net196));
 sky130_fd_sc_hd__diode_2 ANTENNA_output198_A (.DIODE(net198));
 sky130_fd_sc_hd__diode_2 ANTENNA__6687__A1 (.DIODE(net198));
 sky130_fd_sc_hd__diode_2 ANTENNA__6487__A1 (.DIODE(net198));
 sky130_fd_sc_hd__diode_2 ANTENNA__5695__A1 (.DIODE(net198));
 sky130_fd_sc_hd__diode_2 ANTENNA__4795__A1 (.DIODE(net198));
 sky130_fd_sc_hd__diode_2 ANTENNA__4181__A1 (.DIODE(net198));
 sky130_fd_sc_hd__diode_2 ANTENNA_output199_A (.DIODE(net199));
 sky130_fd_sc_hd__diode_2 ANTENNA__6689__A1 (.DIODE(net199));
 sky130_fd_sc_hd__diode_2 ANTENNA__5725__A1 (.DIODE(net199));
 sky130_fd_sc_hd__diode_2 ANTENNA__4184__A1 (.DIODE(net199));
 sky130_fd_sc_hd__diode_2 ANTENNA_output200_A (.DIODE(net200));
 sky130_fd_sc_hd__diode_2 ANTENNA__6691__A1 (.DIODE(net200));
 sky130_fd_sc_hd__diode_2 ANTENNA__6505__B1 (.DIODE(net200));
 sky130_fd_sc_hd__diode_2 ANTENNA__5755__A1 (.DIODE(net200));
 sky130_fd_sc_hd__diode_2 ANTENNA__4187__A1 (.DIODE(net200));
 sky130_fd_sc_hd__diode_2 ANTENNA_output201_A (.DIODE(net201));
 sky130_fd_sc_hd__diode_2 ANTENNA__6763__A (.DIODE(net201));
 sky130_fd_sc_hd__diode_2 ANTENNA__6716__A0 (.DIODE(net201));
 sky130_fd_sc_hd__diode_2 ANTENNA__6662__A1 (.DIODE(net201));
 sky130_fd_sc_hd__diode_2 ANTENNA__6640__A1 (.DIODE(net201));
 sky130_fd_sc_hd__diode_2 ANTENNA__6570__A0 (.DIODE(net201));
 sky130_fd_sc_hd__diode_2 ANTENNA__6523__A1 (.DIODE(net201));
 sky130_fd_sc_hd__diode_2 ANTENNA__5278__A1 (.DIODE(net201));
 sky130_fd_sc_hd__diode_2 ANTENNA__4899__B2 (.DIODE(net201));
 sky130_fd_sc_hd__diode_2 ANTENNA__4147__A1 (.DIODE(net201));
 sky130_fd_sc_hd__diode_2 ANTENNA_output202_A (.DIODE(net202));
 sky130_fd_sc_hd__diode_2 ANTENNA__6722__A1 (.DIODE(net202));
 sky130_fd_sc_hd__diode_2 ANTENNA__6664__A1 (.DIODE(net202));
 sky130_fd_sc_hd__diode_2 ANTENNA__6643__A1 (.DIODE(net202));
 sky130_fd_sc_hd__diode_2 ANTENNA__6527__A1 (.DIODE(net202));
 sky130_fd_sc_hd__diode_2 ANTENNA__6161__A2 (.DIODE(net202));
 sky130_fd_sc_hd__diode_2 ANTENNA__5324__A1 (.DIODE(net202));
 sky130_fd_sc_hd__diode_2 ANTENNA__4451__A1 (.DIODE(net202));
 sky130_fd_sc_hd__diode_2 ANTENNA_output203_A (.DIODE(net203));
 sky130_fd_sc_hd__diode_2 ANTENNA__6769__A (.DIODE(net203));
 sky130_fd_sc_hd__diode_2 ANTENNA__6728__A1 (.DIODE(net203));
 sky130_fd_sc_hd__diode_2 ANTENNA__6666__A1 (.DIODE(net203));
 sky130_fd_sc_hd__diode_2 ANTENNA__6583__A0 (.DIODE(net203));
 sky130_fd_sc_hd__diode_2 ANTENNA__6535__A (.DIODE(net203));
 sky130_fd_sc_hd__diode_2 ANTENNA__6430__B1 (.DIODE(net203));
 sky130_fd_sc_hd__diode_2 ANTENNA__5362__A1 (.DIODE(net203));
 sky130_fd_sc_hd__diode_2 ANTENNA__4448__A2 (.DIODE(net203));
 sky130_fd_sc_hd__diode_2 ANTENNA__4150__A1 (.DIODE(net203));
 sky130_fd_sc_hd__diode_2 ANTENNA_output204_A (.DIODE(net204));
 sky130_fd_sc_hd__diode_2 ANTENNA__6668__A1 (.DIODE(net204));
 sky130_fd_sc_hd__diode_2 ANTENNA__6556__A (.DIODE(net204));
 sky130_fd_sc_hd__diode_2 ANTENNA__6435__B1 (.DIODE(net204));
 sky130_fd_sc_hd__diode_2 ANTENNA__4440__A1 (.DIODE(net204));
 sky130_fd_sc_hd__diode_2 ANTENNA__4153__A1 (.DIODE(net204));
 sky130_fd_sc_hd__diode_2 ANTENNA_output205_A (.DIODE(net205));
 sky130_fd_sc_hd__diode_2 ANTENNA__6740__A1 (.DIODE(net205));
 sky130_fd_sc_hd__diode_2 ANTENNA__6670__A1 (.DIODE(net205));
 sky130_fd_sc_hd__diode_2 ANTENNA__5437__A1 (.DIODE(net205));
 sky130_fd_sc_hd__diode_2 ANTENNA__4156__A1 (.DIODE(net205));
 sky130_fd_sc_hd__diode_2 ANTENNA_output206_A (.DIODE(net206));
 sky130_fd_sc_hd__diode_2 ANTENNA__6746__A1 (.DIODE(net206));
 sky130_fd_sc_hd__diode_2 ANTENNA__6673__A1 (.DIODE(net206));
 sky130_fd_sc_hd__diode_2 ANTENNA__5472__A1 (.DIODE(net206));
 sky130_fd_sc_hd__diode_2 ANTENNA__4431__A1 (.DIODE(net206));
 sky130_fd_sc_hd__diode_2 ANTENNA__4159__A1 (.DIODE(net206));
 sky130_fd_sc_hd__diode_2 ANTENNA_output207_A (.DIODE(net207));
 sky130_fd_sc_hd__diode_2 ANTENNA__6752__A1 (.DIODE(net207));
 sky130_fd_sc_hd__diode_2 ANTENNA__6675__A1 (.DIODE(net207));
 sky130_fd_sc_hd__diode_2 ANTENNA__6451__A1 (.DIODE(net207));
 sky130_fd_sc_hd__diode_2 ANTENNA__5510__A1 (.DIODE(net207));
 sky130_fd_sc_hd__diode_2 ANTENNA__4162__A1 (.DIODE(net207));
 sky130_fd_sc_hd__diode_2 ANTENNA_output208_A (.DIODE(net208));
 sky130_fd_sc_hd__diode_2 ANTENNA__6677__A1 (.DIODE(net208));
 sky130_fd_sc_hd__diode_2 ANTENNA__6459__B1 (.DIODE(net208));
 sky130_fd_sc_hd__diode_2 ANTENNA__5538__A1 (.DIODE(net208));
 sky130_fd_sc_hd__diode_2 ANTENNA__4426__A1 (.DIODE(net208));
 sky130_fd_sc_hd__diode_2 ANTENNA__4165__A1 (.DIODE(net208));
 sky130_fd_sc_hd__diode_2 ANTENNA_output209_A (.DIODE(net209));
 sky130_fd_sc_hd__diode_2 ANTENNA__6679__A1 (.DIODE(net209));
 sky130_fd_sc_hd__diode_2 ANTENNA__5572__A1 (.DIODE(net209));
 sky130_fd_sc_hd__diode_2 ANTENNA__4169__A1 (.DIODE(net209));
 sky130_fd_sc_hd__diode_2 ANTENNA_output210_A (.DIODE(net210));
 sky130_fd_sc_hd__diode_2 ANTENNA__4139__A (.DIODE(net210));
 sky130_fd_sc_hd__diode_2 ANTENNA__3788__A1 (.DIODE(net211));
 sky130_fd_sc_hd__diode_2 ANTENNA_output72_A (.DIODE(net211));
 sky130_fd_sc_hd__diode_2 ANTENNA__6564__A0 (.DIODE(net211));
 sky130_fd_sc_hd__diode_2 ANTENNA__6419__B (.DIODE(net211));
 sky130_fd_sc_hd__diode_2 ANTENNA__6418__A1 (.DIODE(net211));
 sky130_fd_sc_hd__diode_2 ANTENNA__6413__A (.DIODE(net211));
 sky130_fd_sc_hd__diode_2 ANTENNA__5196__A (.DIODE(net211));
 sky130_fd_sc_hd__diode_2 ANTENNA__5193__A (.DIODE(net211));
 sky130_fd_sc_hd__diode_2 ANTENNA__4778__A (.DIODE(net211));
 sky130_fd_sc_hd__diode_2 ANTENNA__4771__A1 (.DIODE(net211));
 sky130_fd_sc_hd__diode_2 ANTENNA__6974__CLK (.DIODE(clknet_leaf_1_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6973__CLK (.DIODE(clknet_leaf_1_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7204__CLK (.DIODE(clknet_leaf_1_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7202__CLK (.DIODE(clknet_leaf_1_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7201__CLK (.DIODE(clknet_leaf_1_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7213__CLK (.DIODE(clknet_leaf_2_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6970__CLK (.DIODE(clknet_leaf_2_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7206__CLK (.DIODE(clknet_leaf_2_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7221__CLK (.DIODE(clknet_leaf_2_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7214__CLK (.DIODE(clknet_leaf_2_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7218__CLK (.DIODE(clknet_leaf_2_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7219__CLK (.DIODE(clknet_leaf_2_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7217__CLK (.DIODE(clknet_leaf_2_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7208__CLK (.DIODE(clknet_leaf_2_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7207__CLK (.DIODE(clknet_leaf_2_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7203__CLK (.DIODE(clknet_leaf_2_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7209__CLK (.DIODE(clknet_leaf_2_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7210__CLK (.DIODE(clknet_leaf_2_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6969__CLK (.DIODE(clknet_leaf_3_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6851__CLK (.DIODE(clknet_leaf_3_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6957__CLK (.DIODE(clknet_leaf_3_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6956__CLK (.DIODE(clknet_leaf_3_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6955__CLK (.DIODE(clknet_leaf_3_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6958__CLK (.DIODE(clknet_leaf_3_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7124__CLK (.DIODE(clknet_leaf_5_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7155__CLK (.DIODE(clknet_leaf_5_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7060__CLK (.DIODE(clknet_leaf_5_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7156__CLK (.DIODE(clknet_leaf_5_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7123__CLK (.DIODE(clknet_leaf_5_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7128__CLK (.DIODE(clknet_leaf_5_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7064__CLK (.DIODE(clknet_leaf_5_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7129__CLK (.DIODE(clknet_leaf_5_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7065__CLK (.DIODE(clknet_leaf_5_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7140__CLK (.DIODE(clknet_leaf_6_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7076__CLK (.DIODE(clknet_leaf_6_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7078__CLK (.DIODE(clknet_leaf_6_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7142__CLK (.DIODE(clknet_leaf_6_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7141__CLK (.DIODE(clknet_leaf_6_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7077__CLK (.DIODE(clknet_leaf_6_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7093__CLK (.DIODE(clknet_leaf_6_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7125__CLK (.DIODE(clknet_leaf_6_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7094__CLK (.DIODE(clknet_leaf_6_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7062__CLK (.DIODE(clknet_leaf_6_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7157__CLK (.DIODE(clknet_leaf_6_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7126__CLK (.DIODE(clknet_leaf_6_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7110__CLK (.DIODE(clknet_leaf_6_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7107__CLK (.DIODE(clknet_leaf_6_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7108__CLK (.DIODE(clknet_leaf_6_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7139__CLK (.DIODE(clknet_leaf_6_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7075__CLK (.DIODE(clknet_leaf_6_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7091__CLK (.DIODE(clknet_leaf_6_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7092__CLK (.DIODE(clknet_leaf_6_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7212__CLK (.DIODE(clknet_leaf_7_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6962__CLK (.DIODE(clknet_leaf_7_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6961__CLK (.DIODE(clknet_leaf_7_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6960__CLK (.DIODE(clknet_leaf_7_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6959__CLK (.DIODE(clknet_leaf_7_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6965__CLK (.DIODE(clknet_leaf_7_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6966__CLK (.DIODE(clknet_leaf_7_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6964__CLK (.DIODE(clknet_leaf_7_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6963__CLK (.DIODE(clknet_leaf_7_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7137__CLK (.DIODE(clknet_leaf_9_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7070__CLK (.DIODE(clknet_leaf_9_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7153__CLK (.DIODE(clknet_leaf_9_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7149__CLK (.DIODE(clknet_leaf_9_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7069__CLK (.DIODE(clknet_leaf_9_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7150__CLK (.DIODE(clknet_leaf_9_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7148__CLK (.DIODE(clknet_leaf_9_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7068__CLK (.DIODE(clknet_leaf_9_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7089__CLK (.DIODE(clknet_leaf_10_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7116__CLK (.DIODE(clknet_leaf_10_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7117__CLK (.DIODE(clknet_leaf_10_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7121__CLK (.DIODE(clknet_leaf_10_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7122__CLK (.DIODE(clknet_leaf_10_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7118__CLK (.DIODE(clknet_leaf_10_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7101__CLK (.DIODE(clknet_leaf_10_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7085__CLK (.DIODE(clknet_leaf_10_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7105__CLK (.DIODE(clknet_leaf_10_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7086__CLK (.DIODE(clknet_leaf_10_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7102__CLK (.DIODE(clknet_leaf_10_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7133__CLK (.DIODE(clknet_leaf_10_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7073__CLK (.DIODE(clknet_leaf_10_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7134__CLK (.DIODE(clknet_leaf_10_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7132__CLK (.DIODE(clknet_leaf_10_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7071__CLK (.DIODE(clknet_leaf_11_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7135__CLK (.DIODE(clknet_leaf_11_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7151__CLK (.DIODE(clknet_leaf_11_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7072__CLK (.DIODE(clknet_leaf_11_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7136__CLK (.DIODE(clknet_leaf_11_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7083__CLK (.DIODE(clknet_leaf_11_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7088__CLK (.DIODE(clknet_leaf_11_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7104__CLK (.DIODE(clknet_leaf_11_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7087__CLK (.DIODE(clknet_leaf_11_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7103__CLK (.DIODE(clknet_leaf_11_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7084__CLK (.DIODE(clknet_leaf_11_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7100__CLK (.DIODE(clknet_leaf_11_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7080__CLK (.DIODE(clknet_leaf_14_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7144__CLK (.DIODE(clknet_leaf_14_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7098__CLK (.DIODE(clknet_leaf_14_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7066__CLK (.DIODE(clknet_leaf_14_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7130__CLK (.DIODE(clknet_leaf_14_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7145__CLK (.DIODE(clknet_leaf_14_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7081__CLK (.DIODE(clknet_leaf_14_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7095__CLK (.DIODE(clknet_leaf_15_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7063__CLK (.DIODE(clknet_leaf_15_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7143__CLK (.DIODE(clknet_leaf_15_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7111__CLK (.DIODE(clknet_leaf_15_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7159__CLK (.DIODE(clknet_leaf_15_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7160__CLK (.DIODE(clknet_leaf_15_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7079__CLK (.DIODE(clknet_leaf_15_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7096__CLK (.DIODE(clknet_leaf_15_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6885__CLK (.DIODE(clknet_leaf_16_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6863__CLK (.DIODE(clknet_leaf_16_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6864__CLK (.DIODE(clknet_leaf_16_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6916__CLK (.DIODE(clknet_leaf_16_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7113__CLK (.DIODE(clknet_leaf_16_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6914__CLK (.DIODE(clknet_leaf_16_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7255__CLK (.DIODE(clknet_leaf_16_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7173__CLK (.DIODE(clknet_leaf_16_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7175__CLK (.DIODE(clknet_leaf_16_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7178__CLK (.DIODE(clknet_leaf_16_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7174__CLK (.DIODE(clknet_leaf_16_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7162__CLK (.DIODE(clknet_leaf_16_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7161__CLK (.DIODE(clknet_leaf_16_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7127__CLK (.DIODE(clknet_leaf_16_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7114__CLK (.DIODE(clknet_leaf_16_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6915__CLK (.DIODE(clknet_leaf_16_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6794__CLK (.DIODE(clknet_leaf_16_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6792__CLK (.DIODE(clknet_leaf_16_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6793__CLK (.DIODE(clknet_leaf_16_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7182__CLK (.DIODE(clknet_leaf_17_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7183__CLK (.DIODE(clknet_leaf_17_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6866__CLK (.DIODE(clknet_leaf_17_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6918__CLK (.DIODE(clknet_leaf_17_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6923__CLK (.DIODE(clknet_leaf_17_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6865__CLK (.DIODE(clknet_leaf_17_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6917__CLK (.DIODE(clknet_leaf_17_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7179__CLK (.DIODE(clknet_leaf_17_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6903__CLK (.DIODE(clknet_leaf_17_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6937__CLK (.DIODE(clknet_leaf_17_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6939__CLK (.DIODE(clknet_leaf_17_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7166__CLK (.DIODE(clknet_leaf_18_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7185__CLK (.DIODE(clknet_leaf_18_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7167__CLK (.DIODE(clknet_leaf_18_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7168__CLK (.DIODE(clknet_leaf_18_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7147__CLK (.DIODE(clknet_leaf_18_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7067__CLK (.DIODE(clknet_leaf_18_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7099__CLK (.DIODE(clknet_leaf_18_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7170__CLK (.DIODE(clknet_leaf_18_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7180__CLK (.DIODE(clknet_leaf_18_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7184__CLK (.DIODE(clknet_leaf_18_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7164__CLK (.DIODE(clknet_leaf_18_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7163__CLK (.DIODE(clknet_leaf_18_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7186__CLK (.DIODE(clknet_leaf_18_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6818__CLK (.DIODE(clknet_leaf_19_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6815__CLK (.DIODE(clknet_leaf_19_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6812__CLK (.DIODE(clknet_leaf_19_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6934__CLK (.DIODE(clknet_leaf_19_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6822__CLK (.DIODE(clknet_leaf_19_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7181__CLK (.DIODE(clknet_leaf_19_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7169__CLK (.DIODE(clknet_leaf_19_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6823__CLK (.DIODE(clknet_leaf_19_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6935__CLK (.DIODE(clknet_leaf_19_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7115__CLK (.DIODE(clknet_leaf_19_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7119__CLK (.DIODE(clknet_leaf_19_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7152__CLK (.DIODE(clknet_leaf_19_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7165__CLK (.DIODE(clknet_leaf_19_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7120__CLK (.DIODE(clknet_leaf_19_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6867__CLK (.DIODE(clknet_leaf_20_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6813__CLK (.DIODE(clknet_leaf_20_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6884__CLK (.DIODE(clknet_leaf_20_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6817__CLK (.DIODE(clknet_leaf_20_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6925__CLK (.DIODE(clknet_leaf_20_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6924__CLK (.DIODE(clknet_leaf_20_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6820__CLK (.DIODE(clknet_leaf_20_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6932__CLK (.DIODE(clknet_leaf_20_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6928__CLK (.DIODE(clknet_leaf_20_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6816__CLK (.DIODE(clknet_leaf_20_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6814__CLK (.DIODE(clknet_leaf_20_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6927__CLK (.DIODE(clknet_leaf_20_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6930__CLK (.DIODE(clknet_leaf_20_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6888__CLK (.DIODE(clknet_leaf_21_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6887__CLK (.DIODE(clknet_leaf_21_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6936__CLK (.DIODE(clknet_leaf_21_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6938__CLK (.DIODE(clknet_leaf_21_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6889__CLK (.DIODE(clknet_leaf_21_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6886__CLK (.DIODE(clknet_leaf_21_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6922__CLK (.DIODE(clknet_leaf_21_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6920__CLK (.DIODE(clknet_leaf_21_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6921__CLK (.DIODE(clknet_leaf_21_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6919__CLK (.DIODE(clknet_leaf_21_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6931__CLK (.DIODE(clknet_leaf_22_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6926__CLK (.DIODE(clknet_leaf_22_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6819__CLK (.DIODE(clknet_leaf_22_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6929__CLK (.DIODE(clknet_leaf_22_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6868__CLK (.DIODE(clknet_leaf_22_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6892__CLK (.DIODE(clknet_leaf_22_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6893__CLK (.DIODE(clknet_leaf_22_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6890__CLK (.DIODE(clknet_leaf_22_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6894__CLK (.DIODE(clknet_leaf_24_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6895__CLK (.DIODE(clknet_leaf_24_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7045__CLK (.DIODE(clknet_leaf_24_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7044__CLK (.DIODE(clknet_leaf_24_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6896__CLK (.DIODE(clknet_leaf_24_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6897__CLK (.DIODE(clknet_leaf_24_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6898__CLK (.DIODE(clknet_leaf_24_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6900__CLK (.DIODE(clknet_leaf_24_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6899__CLK (.DIODE(clknet_leaf_24_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6869__CLK (.DIODE(clknet_leaf_24_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6901__CLK (.DIODE(clknet_leaf_24_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6872__CLK (.DIODE(clknet_leaf_24_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6874__CLK (.DIODE(clknet_leaf_24_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7029__CLK (.DIODE(clknet_leaf_25_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7028__CLK (.DIODE(clknet_leaf_25_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7027__CLK (.DIODE(clknet_leaf_25_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7274__CLK (.DIODE(clknet_leaf_25_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7275__CLK (.DIODE(clknet_leaf_25_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7277__CLK (.DIODE(clknet_leaf_25_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6849__CLK (.DIODE(clknet_leaf_25_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7278__CLK (.DIODE(clknet_leaf_25_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6846__CLK (.DIODE(clknet_leaf_25_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6891__CLK (.DIODE(clknet_leaf_25_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7279__CLK (.DIODE(clknet_leaf_25_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7276__CLK (.DIODE(clknet_leaf_25_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6861__CLK (.DIODE(clknet_leaf_25_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6860__CLK (.DIODE(clknet_leaf_26_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7040__CLK (.DIODE(clknet_leaf_26_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7024__CLK (.DIODE(clknet_leaf_26_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7025__CLK (.DIODE(clknet_leaf_26_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7041__CLK (.DIODE(clknet_leaf_26_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7042__CLK (.DIODE(clknet_leaf_26_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6862__CLK (.DIODE(clknet_leaf_26_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7043__CLK (.DIODE(clknet_leaf_26_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7234__CLK (.DIODE(clknet_leaf_27_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7230__CLK (.DIODE(clknet_leaf_27_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7273__CLK (.DIODE(clknet_leaf_27_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6845__CLK (.DIODE(clknet_leaf_27_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7272__CLK (.DIODE(clknet_leaf_27_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7023__CLK (.DIODE(clknet_leaf_27_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6844__CLK (.DIODE(clknet_leaf_27_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7022__CLK (.DIODE(clknet_leaf_27_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7039__CLK (.DIODE(clknet_leaf_27_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6850__CLK (.DIODE(clknet_leaf_28_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6848__CLK (.DIODE(clknet_leaf_28_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7026__CLK (.DIODE(clknet_leaf_28_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7232__CLK (.DIODE(clknet_leaf_28_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7231__CLK (.DIODE(clknet_leaf_28_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7233__CLK (.DIODE(clknet_leaf_28_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7236__CLK (.DIODE(clknet_leaf_28_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6990__CLK (.DIODE(clknet_leaf_29_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6991__CLK (.DIODE(clknet_leaf_29_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7253__CLK (.DIODE(clknet_leaf_29_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7254__CLK (.DIODE(clknet_leaf_29_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7257__CLK (.DIODE(clknet_leaf_29_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7256__CLK (.DIODE(clknet_leaf_29_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6847__CLK (.DIODE(clknet_leaf_29_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7171__CLK (.DIODE(clknet_leaf_30_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7172__CLK (.DIODE(clknet_leaf_30_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6993__CLK (.DIODE(clknet_leaf_30_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7176__CLK (.DIODE(clknet_leaf_30_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6992__CLK (.DIODE(clknet_leaf_30_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7013__CLK (.DIODE(clknet_leaf_30_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6987__CLK (.DIODE(clknet_leaf_30_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6986__CLK (.DIODE(clknet_leaf_30_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7250__CLK (.DIODE(clknet_leaf_30_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7251__CLK (.DIODE(clknet_leaf_30_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6989__CLK (.DIODE(clknet_leaf_30_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7252__CLK (.DIODE(clknet_leaf_30_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6988__CLK (.DIODE(clknet_leaf_30_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6796__CLK (.DIODE(clknet_leaf_31_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6800__CLK (.DIODE(clknet_leaf_31_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7005__CLK (.DIODE(clknet_leaf_31_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7205__CLK (.DIODE(clknet_leaf_31_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7046__CLK (.DIODE(clknet_leaf_31_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7051__CLK (.DIODE(clknet_leaf_31_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7050__CLK (.DIODE(clknet_leaf_31_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7097__CLK (.DIODE(clknet_leaf_31_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6791__CLK (.DIODE(clknet_leaf_31_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7177__CLK (.DIODE(clknet_leaf_31_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7112__CLK (.DIODE(clknet_leaf_31_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7248__CLK (.DIODE(clknet_leaf_32_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7249__CLK (.DIODE(clknet_leaf_32_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6985__CLK (.DIODE(clknet_leaf_32_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6983__CLK (.DIODE(clknet_leaf_32_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6980__CLK (.DIODE(clknet_leaf_32_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7054__CLK (.DIODE(clknet_leaf_32_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6940__CLK (.DIODE(clknet_leaf_32_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6902__CLK (.DIODE(clknet_leaf_32_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6941__CLK (.DIODE(clknet_leaf_32_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6835__CLK (.DIODE(clknet_leaf_32_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7244__CLK (.DIODE(clknet_leaf_33_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7245__CLK (.DIODE(clknet_leaf_33_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7242__CLK (.DIODE(clknet_leaf_33_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6979__CLK (.DIODE(clknet_leaf_33_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6984__CLK (.DIODE(clknet_leaf_33_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6978__CLK (.DIODE(clknet_leaf_33_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7246__CLK (.DIODE(clknet_leaf_33_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6843__CLK (.DIODE(clknet_leaf_35_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7222__CLK (.DIODE(clknet_leaf_35_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7227__CLK (.DIODE(clknet_leaf_35_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7226__CLK (.DIODE(clknet_leaf_35_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7229__CLK (.DIODE(clknet_leaf_35_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7228__CLK (.DIODE(clknet_leaf_35_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7247__CLK (.DIODE(clknet_leaf_35_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6982__CLK (.DIODE(clknet_leaf_35_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7225__CLK (.DIODE(clknet_leaf_35_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6842__CLK (.DIODE(clknet_leaf_35_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6856__CLK (.DIODE(clknet_leaf_36_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7030__CLK (.DIODE(clknet_leaf_36_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7014__CLK (.DIODE(clknet_leaf_36_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7015__CLK (.DIODE(clknet_leaf_36_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7018__CLK (.DIODE(clknet_leaf_36_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7270__CLK (.DIODE(clknet_leaf_36_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7271__CLK (.DIODE(clknet_leaf_36_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7019__CLK (.DIODE(clknet_leaf_36_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6857__CLK (.DIODE(clknet_leaf_36_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7035__CLK (.DIODE(clknet_leaf_36_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7036__CLK (.DIODE(clknet_leaf_36_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6858__CLK (.DIODE(clknet_leaf_36_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7037__CLK (.DIODE(clknet_leaf_36_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6859__CLK (.DIODE(clknet_leaf_36_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7038__CLK (.DIODE(clknet_leaf_36_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7020__CLK (.DIODE(clknet_leaf_36_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7021__CLK (.DIODE(clknet_leaf_36_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6852__CLK (.DIODE(clknet_leaf_39_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6999__CLK (.DIODE(clknet_leaf_39_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6994__CLK (.DIODE(clknet_leaf_39_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7289__CLK (.DIODE(clknet_leaf_39_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7290__CLK (.DIODE(clknet_leaf_39_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6837__CLK (.DIODE(clknet_leaf_39_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6976__CLK (.DIODE(clknet_leaf_39_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7291__CLK (.DIODE(clknet_leaf_39_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6853__CLK (.DIODE(clknet_leaf_39_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7031__CLK (.DIODE(clknet_leaf_39_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7267__CLK (.DIODE(clknet_leaf_39_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7032__CLK (.DIODE(clknet_leaf_39_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6854__CLK (.DIODE(clknet_leaf_39_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7269__CLK (.DIODE(clknet_leaf_39_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6840__CLK (.DIODE(clknet_leaf_39_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6838__CLK (.DIODE(clknet_leaf_39_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7266__CLK (.DIODE(clknet_leaf_39_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7264__CLK (.DIODE(clknet_leaf_39_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7265__CLK (.DIODE(clknet_leaf_39_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7285__CLK (.DIODE(clknet_leaf_40_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7294__CLK (.DIODE(clknet_leaf_40_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7287__CLK (.DIODE(clknet_leaf_40_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7298__CLK (.DIODE(clknet_leaf_40_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7288__CLK (.DIODE(clknet_leaf_40_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7286__CLK (.DIODE(clknet_leaf_40_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7296__CLK (.DIODE(clknet_leaf_40_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6996__CLK (.DIODE(clknet_leaf_40_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7001__CLK (.DIODE(clknet_leaf_40_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7000__CLK (.DIODE(clknet_leaf_40_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6997__CLK (.DIODE(clknet_leaf_40_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6995__CLK (.DIODE(clknet_leaf_40_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6998__CLK (.DIODE(clknet_leaf_40_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6977__CLK (.DIODE(clknet_leaf_40_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7299__CLK (.DIODE(clknet_leaf_41_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7292__CLK (.DIODE(clknet_leaf_41_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7297__CLK (.DIODE(clknet_leaf_41_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7295__CLK (.DIODE(clknet_leaf_41_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7293__CLK (.DIODE(clknet_leaf_41_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7263__CLK (.DIODE(clknet_leaf_41_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7002__CLK (.DIODE(clknet_leaf_41_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7280__CLK (.DIODE(clknet_leaf_41_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7284__CLK (.DIODE(clknet_leaf_41_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7281__CLK (.DIODE(clknet_leaf_42_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7261__CLK (.DIODE(clknet_leaf_42_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7258__CLK (.DIODE(clknet_leaf_42_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6910__CLK (.DIODE(clknet_leaf_42_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6909__CLK (.DIODE(clknet_leaf_42_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6904__CLK (.DIODE(clknet_leaf_42_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7004__CLK (.DIODE(clknet_leaf_42_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6825__CLK (.DIODE(clknet_leaf_42_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6828__CLK (.DIODE(clknet_leaf_42_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6829__CLK (.DIODE(clknet_leaf_42_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6908__CLK (.DIODE(clknet_leaf_42_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6905__CLK (.DIODE(clknet_leaf_42_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7300__CLK (.DIODE(clknet_leaf_42_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6836__CLK (.DIODE(clknet_leaf_42_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6831__CLK (.DIODE(clknet_leaf_42_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6833__CLK (.DIODE(clknet_leaf_45_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6785__CLK (.DIODE(clknet_leaf_45_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6807__CLK (.DIODE(clknet_leaf_45_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6830__CLK (.DIODE(clknet_leaf_45_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6827__CLK (.DIODE(clknet_leaf_45_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6803__CLK (.DIODE(clknet_leaf_45_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6826__CLK (.DIODE(clknet_leaf_45_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6787__CLK (.DIODE(clknet_leaf_45_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7239__CLK (.DIODE(clknet_leaf_45_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6786__CLK (.DIODE(clknet_leaf_45_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6784__CLK (.DIODE(clknet_leaf_45_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6946__CLK (.DIODE(clknet_leaf_45_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6788__CLK (.DIODE(clknet_leaf_45_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6948__CLK (.DIODE(clknet_leaf_45_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6943__CLK (.DIODE(clknet_leaf_45_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6944__CLK (.DIODE(clknet_leaf_45_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7240__CLK (.DIODE(clknet_leaf_46_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7241__CLK (.DIODE(clknet_leaf_46_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6804__CLK (.DIODE(clknet_leaf_46_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6805__CLK (.DIODE(clknet_leaf_46_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7237__CLK (.DIODE(clknet_leaf_46_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6802__CLK (.DIODE(clknet_leaf_46_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6913__CLK (.DIODE(clknet_leaf_46_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6912__CLK (.DIODE(clknet_leaf_46_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7056__CLK (.DIODE(clknet_leaf_46_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7057__CLK (.DIODE(clknet_leaf_46_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7055__CLK (.DIODE(clknet_leaf_46_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6824__CLK (.DIODE(clknet_leaf_46_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6806__CLK (.DIODE(clknet_leaf_46_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6975__CLK (.DIODE(clknet_leaf_46_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6810__CLK (.DIODE(clknet_leaf_46_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6811__CLK (.DIODE(clknet_leaf_46_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7243__CLK (.DIODE(clknet_leaf_46_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6808__CLK (.DIODE(clknet_leaf_46_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6809__CLK (.DIODE(clknet_leaf_46_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7006__CLK (.DIODE(clknet_leaf_47_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7009__CLK (.DIODE(clknet_leaf_47_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7008__CLK (.DIODE(clknet_leaf_47_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7007__CLK (.DIODE(clknet_leaf_47_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7012__CLK (.DIODE(clknet_leaf_47_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7047__CLK (.DIODE(clknet_leaf_47_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7048__CLK (.DIODE(clknet_leaf_47_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7011__CLK (.DIODE(clknet_leaf_47_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7010__CLK (.DIODE(clknet_leaf_47_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6797__CLK (.DIODE(clknet_leaf_47_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6799__CLK (.DIODE(clknet_leaf_47_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6795__CLK (.DIODE(clknet_leaf_47_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6911__CLK (.DIODE(clknet_leaf_47_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7058__CLK (.DIODE(clknet_leaf_47_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6801__CLK (.DIODE(clknet_leaf_47_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6798__CLK (.DIODE(clknet_leaf_47_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7052__CLK (.DIODE(clknet_leaf_47_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7053__CLK (.DIODE(clknet_leaf_47_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7049__CLK (.DIODE(clknet_leaf_47_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6951__CLK (.DIODE(clknet_leaf_47_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7238__CLK (.DIODE(clknet_leaf_47_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7192__CLK (.DIODE(clknet_leaf_49_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7193__CLK (.DIODE(clknet_leaf_49_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7194__CLK (.DIODE(clknet_leaf_49_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7191__CLK (.DIODE(clknet_leaf_49_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6949__CLK (.DIODE(clknet_leaf_49_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7189__CLK (.DIODE(clknet_leaf_50_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7199__CLK (.DIODE(clknet_leaf_50_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7198__CLK (.DIODE(clknet_leaf_50_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7197__CLK (.DIODE(clknet_leaf_50_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7196__CLK (.DIODE(clknet_leaf_50_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7200__CLK (.DIODE(clknet_leaf_50_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7195__CLK (.DIODE(clknet_leaf_50_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_1_0_i_clk_A (.DIODE(clknet_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0_0_i_clk_A (.DIODE(clknet_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_2_1_0_i_clk_A (.DIODE(clknet_1_0_1_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_2_0_0_i_clk_A (.DIODE(clknet_1_0_1_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_2_3_0_i_clk_A (.DIODE(clknet_1_1_1_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_2_2_0_i_clk_A (.DIODE(clknet_1_1_1_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_50_i_clk_A (.DIODE(clknet_2_0_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_49_i_clk_A (.DIODE(clknet_2_0_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_opt_1_0_i_clk_A (.DIODE(clknet_2_0_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_47_i_clk_A (.DIODE(clknet_2_0_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_44_i_clk_A (.DIODE(clknet_2_0_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_4_i_clk_A (.DIODE(clknet_2_0_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_3_i_clk_A (.DIODE(clknet_2_0_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_2_i_clk_A (.DIODE(clknet_2_0_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_1_i_clk_A (.DIODE(clknet_2_0_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_0_i_clk_A (.DIODE(clknet_2_0_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_46_i_clk_A (.DIODE(clknet_2_1_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_45_i_clk_A (.DIODE(clknet_2_1_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_43_i_clk_A (.DIODE(clknet_2_1_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_42_i_clk_A (.DIODE(clknet_2_1_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_41_i_clk_A (.DIODE(clknet_2_1_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_40_i_clk_A (.DIODE(clknet_2_1_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_39_i_clk_A (.DIODE(clknet_2_1_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_38_i_clk_A (.DIODE(clknet_2_1_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_37_i_clk_A (.DIODE(clknet_2_1_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_36_i_clk_A (.DIODE(clknet_2_1_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_35_i_clk_A (.DIODE(clknet_2_1_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_34_i_clk_A (.DIODE(clknet_2_1_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_33_i_clk_A (.DIODE(clknet_2_1_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_32_i_clk_A (.DIODE(clknet_2_1_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_31_i_clk_A (.DIODE(clknet_2_1_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_15_i_clk_A (.DIODE(clknet_2_2_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_14_i_clk_A (.DIODE(clknet_2_2_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_13_i_clk_A (.DIODE(clknet_2_2_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_12_i_clk_A (.DIODE(clknet_2_2_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_11_i_clk_A (.DIODE(clknet_2_2_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_10_i_clk_A (.DIODE(clknet_2_2_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_9_i_clk_A (.DIODE(clknet_2_2_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_8_i_clk_A (.DIODE(clknet_2_2_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_7_i_clk_A (.DIODE(clknet_2_2_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_6_i_clk_A (.DIODE(clknet_2_2_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_5_i_clk_A (.DIODE(clknet_2_2_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_30_i_clk_A (.DIODE(clknet_2_3_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_29_i_clk_A (.DIODE(clknet_2_3_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_28_i_clk_A (.DIODE(clknet_2_3_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_27_i_clk_A (.DIODE(clknet_2_3_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_26_i_clk_A (.DIODE(clknet_2_3_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_25_i_clk_A (.DIODE(clknet_2_3_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_24_i_clk_A (.DIODE(clknet_2_3_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_opt_2_0_i_clk_A (.DIODE(clknet_2_3_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_22_i_clk_A (.DIODE(clknet_2_3_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_21_i_clk_A (.DIODE(clknet_2_3_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_20_i_clk_A (.DIODE(clknet_2_3_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_19_i_clk_A (.DIODE(clknet_2_3_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_18_i_clk_A (.DIODE(clknet_2_3_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_17_i_clk_A (.DIODE(clknet_2_3_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_16_i_clk_A (.DIODE(clknet_2_3_0_i_clk));
 sky130_ef_sc_hd__decap_12 FILLER_0_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_685 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_769 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_797 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_825 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_447 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_457 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_486 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_492 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_521 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_525 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_537 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_839 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_433 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_494 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_500 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_506 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_512 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_518 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_537 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_543 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_555 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_567 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_417 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_463 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_519 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_525 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_538 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_544 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_558 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_570 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_576 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_588 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_612 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_839 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_436 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_459 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_514 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_523 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_538 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_550 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_557 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_417 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_462 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_470 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_484 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_495 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_519 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_524 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_565 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_571 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_747 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_753 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_774 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_780 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_797 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_815 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_827 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_839 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_419 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_442 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_486 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_495 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_512 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_525 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_539 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_547 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_555 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_580 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_719 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_739 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_745 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_753 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_767 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_773 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_797 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_831 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_424 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_447 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_467 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_481 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_487 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_495 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_518 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_530 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_536 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_542 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_558 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_567 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_685 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_697 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_704 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_712 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_716 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_720 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_741 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_749 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_753 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_759 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_771 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_803 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_811 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_815 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_823 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_827 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_839 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_439 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_448 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_454 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_487 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_493 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_504 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_522 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_537 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_549 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_563 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_672 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_684 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_696 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_708 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_717 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_723 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_735 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_741 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_744 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_754 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_763 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_773 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_791 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_797 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_803 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_813 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_817 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_823 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_435 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_470 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_476 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_482 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_494 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_515 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_521 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_553 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_558 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_567 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_574 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_594 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_637 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_641 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_661 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_678 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_690 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_702 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_726 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_735 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_738 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_748 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_762 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_775 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_793 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_799 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_819 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_825 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_833 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_551 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_563 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_642 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_654 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_660 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_664 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_670 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_678 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_699 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_708 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_714 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_726 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_738 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_746 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_754 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_769 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_775 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_778 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_791 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_799 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_806 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_813 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_831 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_834 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_417 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_437 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_461 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_500 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_513 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_526 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_536 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_544 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_577 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_583 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_595 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_625 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_635 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_641 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_649 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_666 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_695 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_720 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_745 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_766 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_772 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_797 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_803 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_811 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_815 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_823 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_826 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_440 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_452 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_464 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_468 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_472 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_491 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_508 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_514 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_518 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_521 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_549 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_559 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_566 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_578 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_607 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_625 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_643 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_651 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_659 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_683 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_689 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_699 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_707 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_724 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_731 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_735 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_744 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_750 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_777 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_783 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_795 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_803 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_808 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_833 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_471 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_494 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_512 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_519 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_526 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_532 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_538 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_555 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_575 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_581 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_587 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_605 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_621 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_633 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_643 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_647 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_654 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_660 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_666 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_682 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_691 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_697 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_706 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_714 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_720 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_747 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_759 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_771 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_797 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_800 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_806 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_814 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_823 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_829 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_833 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_419 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_431 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_435 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_440 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_463 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_498 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_509 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_542 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_553 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_567 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_577 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_598 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_605 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_609 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_619 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_625 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_635 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_641 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_650 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_662 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_680 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_684 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_687 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_710 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_716 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_732 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_736 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_745 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_761 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_767 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_773 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_779 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_791 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_813 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_823 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_829 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_833 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_413 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_424 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_527 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_540 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_548 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_576 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_582 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_590 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_625 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_632 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_639 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_648 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_654 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_666 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_685 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_697 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_700 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_708 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_712 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_715 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_743 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_749 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_755 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_761 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_767 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_804 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_811 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_817 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_823 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_831 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_419 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_499 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_514 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_523 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_529 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_541 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_551 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_558 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_579 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_585 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_623 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_633 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_652 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_658 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_670 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_682 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_706 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_719 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_734 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_740 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_746 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_754 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_772 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_778 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_786 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_817 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_823 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_435 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_453 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_466 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_478 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_502 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_522 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_528 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_534 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_538 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_544 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_552 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_565 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_571 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_577 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_585 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_591 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_603 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_631 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_640 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_647 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_658 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_678 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_690 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_702 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_710 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_722 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_741 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_753 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_761 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_766 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_792 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_798 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_804 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_810 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_814 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_822 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_828 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_419 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_439 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_501 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_513 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_537 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_540 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_552 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_560 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_576 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_598 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_604 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_614 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_623 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_632 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_649 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_655 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_675 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_725 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_738 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_742 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_745 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_753 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_763 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_771 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_777 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_783 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_789 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_800 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_806 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_820 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_433 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_473 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_485 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_509 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_515 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_518 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_526 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_529 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_535 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_575 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_595 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_621 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_634 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_640 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_646 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_652 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_664 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_673 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_681 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_686 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_692 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_706 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_710 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_714 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_717 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_725 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_734 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_743 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_749 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_764 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_772 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_792 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_800 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_434 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_440 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_448 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_464 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_507 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_519 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_543 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_557 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_562 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_566 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_593 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_599 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_602 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_616 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_628 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_649 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_655 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_661 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_680 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_705 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_709 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_715 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_719 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_723 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_744 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_750 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_767 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_774 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_780 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_786 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_792 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_798 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_804 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_810 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_819 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_823 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_413 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_475 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_516 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_520 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_527 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_534 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_541 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_547 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_578 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_584 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_596 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_608 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_637 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_644 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_655 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_661 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_684 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_691 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_702 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_719 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_725 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_733 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_739 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_753 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_766 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_772 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_778 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_789 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_795 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_807 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_829 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_833 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_428 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_436 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_500 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_512 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_538 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_545 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_551 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_577 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_625 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_628 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_632 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_635 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_652 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_661 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_668 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_674 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_684 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_690 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_706 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_714 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_718 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_735 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_743 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_746 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_752 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_763 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_779 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_782 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_798 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_804 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_818 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_428 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_472 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_484 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_492 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_515 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_521 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_525 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_538 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_570 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_605 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_621 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_637 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_670 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_673 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_681 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_686 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_692 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_698 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_702 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_726 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_737 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_743 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_748 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_760 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_766 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_772 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_778 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_789 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_793 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_811 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_817 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_825 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_839 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_377 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_430 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_436 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_440 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_443 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_455 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_463 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_487 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_490 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_499 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_506 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_523 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_549 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_562 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_571 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_603 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_612 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_620 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_626 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_660 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_664 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_667 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_679 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_699 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_705 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_708 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_720 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_728 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_742 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_761 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_767 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_776 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_784 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_793 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_804 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_810 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_821 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_824 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_413 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_473 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_495 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_523 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_528 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_534 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_540 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_558 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_567 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_574 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_578 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_599 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_605 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_622 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_628 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_634 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_646 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_652 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_658 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_685 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_691 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_694 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_706 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_726 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_755 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_761 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_791 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_797 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_803 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_809 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_821 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_824 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_377 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_389 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_397 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_403 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_497 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_500 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_527 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_555 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_559 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_565 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_611 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_620 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_626 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_630 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_638 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_645 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_653 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_662 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_670 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_698 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_725 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_735 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_743 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_761 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_767 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_773 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_779 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_791 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_801 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_817 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_828 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_373 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_390 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_415 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_427 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_459 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_471 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_483 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_521 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_527 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_539 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_576 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_590 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_596 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_602 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_635 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_643 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_651 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_661 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_669 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_681 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_687 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_699 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_707 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_747 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_754 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_760 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_766 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_778 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_797 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_809 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_815 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_818 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_377 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_429 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_432 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_440 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_443 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_463 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_482 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_551 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_554 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_560 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_584 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_605 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_610 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_616 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_628 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_669 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_690 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_723 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_745 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_761 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_772 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_776 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_779 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_787 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_791 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_799 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_803 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_831 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_838 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_367 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_370 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_390 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_430 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_434 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_447 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_459 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_465 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_482 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_492 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_529 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_541 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_550 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_565 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_571 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_583 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_595 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_639 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_651 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_657 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_664 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_677 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_694 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_700 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_706 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_712 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_740 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_746 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_756 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_768 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_771 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_789 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_795 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_807 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_815 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_821 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_827 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_369 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_386 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_394 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_400 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_412 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_441 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_454 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_466 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_472 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_502 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_508 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_516 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_553 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_559 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_571 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_625 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_633 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_641 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_667 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_677 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_693 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_713 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_722 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_728 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_731 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_743 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_752 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_761 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_770 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_776 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_780 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_789 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_817 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_829 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_835 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_367 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_424 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_466 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_472 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_510 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_527 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_541 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_550 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_557 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_567 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_574 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_583 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_591 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_603 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_625 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_633 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_644 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_658 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_677 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_683 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_695 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_703 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_707 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_713 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_722 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_733 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_745 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_759 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_790 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_796 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_807 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_821 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_824 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_439 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_472 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_497 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_510 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_545 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_557 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_575 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_595 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_603 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_610 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_619 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_627 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_653 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_660 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_666 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_678 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_698 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_707 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_711 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_717 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_723 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_735 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_743 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_747 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_766 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_783 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_788 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_794 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_800 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_818 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_824 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_828 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_373 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_381 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_386 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_404 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_424 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_435 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_470 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_476 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_500 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_541 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_547 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_582 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_592 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_604 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_614 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_628 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_637 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_646 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_670 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_685 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_697 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_707 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_714 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_741 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_745 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_765 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_771 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_792 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_798 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_804 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_814 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_820 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_831 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_380 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_386 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_396 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_418 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_445 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_463 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_482 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_494 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_506 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_512 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_520 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_549 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_555 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_567 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_621 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_633 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_699 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_714 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_720 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_726 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_730 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_747 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_767 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_773 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_789 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_793 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_796 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_831 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_835 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_361 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_382 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_388 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_398 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_420 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_426 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_485 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_491 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_509 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_527 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_536 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_542 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_548 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_585 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_605 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_625 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_631 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_643 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_655 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_663 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_688 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_700 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_715 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_726 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_740 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_746 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_752 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_758 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_764 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_776 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_797 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_805 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_810 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_823 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_827 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_384 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_406 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_412 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_434 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_450 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_456 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_517 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_551 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_587 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_603 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_610 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_616 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_623 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_629 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_643 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_645 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_653 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_660 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_671 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_679 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_732 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_738 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_744 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_769 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_789 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_792 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_798 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_823 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_830 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_361 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_386 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_400 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_406 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_410 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_432 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_446 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_459 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_469 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_522 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_528 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_542 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_550 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_573 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_585 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_598 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_604 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_624 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_631 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_644 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_650 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_659 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_670 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_695 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_702 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_708 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_714 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_718 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_765 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_777 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_795 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_816 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_822 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_377 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_385 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_402 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_415 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_443 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_497 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_506 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_540 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_549 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_564 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_570 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_576 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_593 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_597 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_639 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_650 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_663 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_683 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_712 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_718 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_730 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_742 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_754 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_757 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_765 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_770 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_790 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_802 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_808 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_819 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_403 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_412 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_420 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_423 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_436 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_457 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_463 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_487 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_521 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_530 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_599 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_605 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_637 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_647 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_654 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_661 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_685 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_707 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_721 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_745 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_751 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_759 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_763 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_769 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_781 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_791 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_799 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_805 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_811 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_817 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_378 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_407 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_435 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_454 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_460 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_497 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_508 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_514 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_520 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_539 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_551 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_560 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_567 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_573 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_593 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_599 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_607 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_627 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_642 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_653 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_656 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_668 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_680 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_698 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_707 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_717 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_723 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_748 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_768 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_776 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_780 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_786 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_792 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_798 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_806 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_810 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_361 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_373 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_409 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_412 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_426 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_434 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_473 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_476 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_495 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_509 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_521 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_550 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_568 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_574 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_580 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_600 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_614 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_631 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_641 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_644 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_651 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_685 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_697 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_700 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_734 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_741 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_747 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_756 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_767 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_773 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_789 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_795 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_801 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_815 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_818 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_825 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_345 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_357 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_369 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_378 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_387 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_415 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_435 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_441 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_453 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_486 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_492 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_498 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_504 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_527 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_551 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_567 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_625 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_633 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_650 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_656 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_659 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_683 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_695 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_698 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_708 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_716 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_720 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_723 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_731 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_737 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_745 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_748 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_767 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_776 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_782 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_788 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_800 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_806 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_818 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_824 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_364 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_370 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_397 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_409 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_431 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_457 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_468 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_489 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_528 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_534 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_540 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_548 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_578 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_595 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_625 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_631 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_644 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_650 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_658 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_677 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_683 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_686 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_694 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_699 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_703 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_706 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_719 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_742 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_750 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_758 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_766 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_772 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_778 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_792 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_796 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_814 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_820 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_826 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_333 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_350 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_374 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_382 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_394 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_406 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_412 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_439 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_452 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_464 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_495 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_501 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_507 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_521 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_543 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_555 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_564 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_576 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_609 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_612 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_625 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_633 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_645 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_676 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_682 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_705 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_711 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_714 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_727 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_748 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_776 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_784 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_795 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_802 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_808 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_819 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_822 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_830 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_838 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_335 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_354 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_366 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_381 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_391 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_417 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_435 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_439 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_456 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_462 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_466 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_469 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_515 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_519 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_527 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_538 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_546 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_565 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_571 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_579 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_591 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_603 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_636 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_650 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_654 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_671 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_679 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_697 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_703 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_711 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_722 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_743 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_749 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_755 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_761 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_768 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_776 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_795 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_805 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_833 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_333 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_375 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_384 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_396 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_409 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_433 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_443 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_454 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_494 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_506 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_516 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_520 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_523 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_547 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_553 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_566 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_575 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_593 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_607 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_624 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_656 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_662 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_679 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_683 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_687 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_698 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_735 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_781 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_787 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_801 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_804 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_823 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_364 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_398 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_406 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_410 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_418 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_430 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_438 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_453 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_469 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_475 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_487 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_509 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_521 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_536 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_542 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_546 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_549 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_586 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_592 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_625 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_637 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_647 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_655 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_658 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_670 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_681 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_691 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_703 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_715 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_733 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_739 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_751 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_763 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_779 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_782 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_797 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_801 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_807 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_811 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_815 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_818 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_824 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_385 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_397 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_406 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_439 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_456 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_496 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_514 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_549 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_557 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_566 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_575 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_593 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_603 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_609 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_633 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_637 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_652 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_664 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_676 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_688 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_706 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_718 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_721 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_745 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_761 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_773 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_778 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_791 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_797 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_806 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_813 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_821 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_827 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_831 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_835 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_381 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_412 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_420 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_426 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_465 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_471 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_494 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_527 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_539 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_559 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_568 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_574 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_580 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_595 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_607 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_638 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_647 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_689 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_693 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_696 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_702 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_711 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_717 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_724 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_736 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_747 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_756 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_762 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_770 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_789 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_795 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_819 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_825 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_373 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_387 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_408 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_426 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_434 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_439 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_455 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_458 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_487 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_493 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_523 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_549 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_555 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_567 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_610 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_616 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_622 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_628 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_642 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_658 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_664 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_667 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_679 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_688 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_719 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_725 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_737 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_741 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_755 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_770 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_783 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_789 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_793 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_810 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_372 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_397 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_406 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_430 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_442 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_466 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_472 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_478 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_502 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_514 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_518 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_521 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_538 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_544 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_568 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_580 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_592 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_604 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_633 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_639 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_651 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_655 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_659 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_697 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_703 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_715 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_725 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_746 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_759 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_789 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_793 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_799 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_806 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_812 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_818 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_355 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_375 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_379 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_382 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_388 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_394 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_400 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_403 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_409 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_454 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_466 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_486 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_492 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_498 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_512 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_519 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_551 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_565 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_642 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_653 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_663 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_669 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_709 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_719 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_728 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_736 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_742 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_754 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_761 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_764 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_774 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_784 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_795 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_801 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_807 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_813 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_341 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_351 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_379 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_407 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_415 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_447 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_469 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_482 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_495 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_509 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_529 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_539 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_567 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_575 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_599 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_611 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_633 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_639 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_647 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_670 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_684 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_699 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_711 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_717 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_733 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_742 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_754 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_760 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_772 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_778 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_789 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_799 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_805 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_811 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_823 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_333 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_340 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_346 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_372 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_378 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_388 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_399 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_419 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_444 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_450 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_475 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_486 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_494 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_498 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_506 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_518 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_539 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_551 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_564 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_603 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_635 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_649 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_655 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_665 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_671 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_683 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_719 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_725 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_737 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_742 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_761 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_778 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_784 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_790 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_798 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_802 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_808 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_821 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_829 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_355 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_374 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_399 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_415 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_435 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_466 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_484 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_488 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_496 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_500 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_510 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_535 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_547 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_568 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_574 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_582 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_596 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_631 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_640 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_646 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_650 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_663 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_687 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_699 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_707 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_715 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_733 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_746 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_758 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_770 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_776 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_789 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_795 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_801 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_807 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_823 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_357 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_381 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_384 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_388 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_399 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_409 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_415 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_432 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_442 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_450 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_463 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_510 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_516 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_530 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_541 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_548 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_560 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_566 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_578 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_585 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_611 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_649 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_655 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_661 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_667 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_679 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_699 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_712 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_718 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_724 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_730 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_736 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_748 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_768 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_774 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_780 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_786 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_806 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_819 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_836 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_345 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_353 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_364 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_377 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_411 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_431 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_453 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_459 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_471 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_483 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_495 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_516 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_540 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_552 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_565 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_571 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_577 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_580 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_598 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_610 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_622 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_628 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_653 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_663 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_684 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_708 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_712 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_718 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_724 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_749 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_759 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_769 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_781 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_789 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_798 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_802 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_819 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_826 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_372 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_384 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_396 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_407 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_443 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_464 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_496 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_500 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_507 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_517 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_531 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_550 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_556 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_560 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_566 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_584 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_663 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_677 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_689 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_695 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_712 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_725 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_731 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_737 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_745 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_750 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_765 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_794 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_798 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_811 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_828 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_335 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_352 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_358 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_364 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_370 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_409 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_415 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_426 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_467 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_479 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_522 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_528 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_551 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_565 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_571 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_583 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_591 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_621 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_633 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_639 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_642 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_648 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_654 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_683 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_710 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_722 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_738 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_755 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_761 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_767 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_773 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_794 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_803 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_809 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_818 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_333 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_351 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_381 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_399 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_409 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_417 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_426 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_436 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_442 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_448 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_460 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_494 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_506 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_542 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_548 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_554 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_562 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_575 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_613 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_625 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_649 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_661 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_666 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_686 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_692 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_709 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_715 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_721 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_733 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_752 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_761 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_767 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_781 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_787 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_793 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_799 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_811 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_818 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_831 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_835 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_373 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_400 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_407 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_413 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_462 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_476 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_482 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_491 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_526 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_536 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_542 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_554 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_570 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_582 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_592 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_604 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_636 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_642 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_654 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_660 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_663 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_684 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_696 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_702 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_710 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_756 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_762 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_768 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_780 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_793 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_809 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_812 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_818 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_824 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_375 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_394 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_402 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_408 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_441 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_459 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_473 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_485 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_491 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_515 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_523 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_546 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_552 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_560 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_563 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_625 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_635 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_660 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_680 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_686 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_710 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_716 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_725 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_741 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_750 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_761 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_773 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_788 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_794 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_800 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_810 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_819 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_348 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_354 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_366 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_370 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_379 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_398 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_410 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_423 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_473 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_485 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_493 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_509 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_521 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_529 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_544 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_569 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_577 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_583 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_595 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_639 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_651 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_677 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_689 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_697 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_700 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_706 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_712 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_742 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_748 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_754 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_766 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_772 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_778 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_789 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_795 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_801 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_807 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_823 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_327 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_344 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_373 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_381 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_397 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_409 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_415 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_435 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_489 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_496 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_512 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_518 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_545 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_554 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_560 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_575 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_593 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_605 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_622 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_628 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_640 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_669 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_681 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_689 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_718 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_724 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_739 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_745 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_753 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_768 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_782 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_788 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_801 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_808 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_823 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_334 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_355 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_361 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_387 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_409 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_418 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_426 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_433 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_473 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_522 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_566 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_572 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_584 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_588 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_594 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_600 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_626 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_632 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_642 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_649 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_655 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_661 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_669 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_681 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_689 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_703 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_709 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_712 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_718 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_724 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_733 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_739 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_759 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_762 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_782 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_789 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_797 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_820 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_826 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_346 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_415 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_439 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_451 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_510 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_522 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_530 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_539 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_548 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_554 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_562 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_566 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_572 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_598 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_610 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_616 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_622 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_634 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_653 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_663 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_675 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_695 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_710 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_716 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_728 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_734 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_744 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_766 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_777 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_786 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_790 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_798 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_818 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_824 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_357 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_366 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_373 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_400 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_407 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_413 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_430 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_454 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_463 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_469 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_484 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_492 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_530 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_542 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_568 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_576 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_584 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_607 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_638 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_644 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_648 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_656 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_677 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_689 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_697 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_704 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_719 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_741 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_745 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_754 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_766 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_772 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_778 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_795 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_801 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_818 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_826 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_387 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_396 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_402 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_408 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_434 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_455 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_494 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_514 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_540 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_547 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_553 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_568 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_574 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_600 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_604 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_607 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_623 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_635 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_656 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_667 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_679 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_709 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_720 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_761 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_765 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_768 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_776 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_779 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_791 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_797 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_803 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_809 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_819 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_373 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_407 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_419 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_436 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_458 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_469 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_481 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_534 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_546 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_550 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_565 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_585 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_603 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_637 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_643 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_650 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_682 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_690 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_696 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_702 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_710 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_718 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_722 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_739 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_743 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_746 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_769 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_781 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_791 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_803 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_806 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_812 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_818 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_825 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_378 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_402 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_481 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_484 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_496 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_508 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_564 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_574 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_580 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_589 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_597 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_602 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_614 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_633 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_649 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_661 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_685 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_697 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_711 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_721 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_732 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_738 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_750 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_781 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_795 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_801 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_807 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_810 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_361 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_378 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_416 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_428 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_453 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_459 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_471 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_482 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_486 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_513 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_518 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_528 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_532 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_536 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_542 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_545 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_559 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_566 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_572 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_596 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_633 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_647 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_659 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_667 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_692 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_698 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_710 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_718 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_747 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_759 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_771 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_774 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_780 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_794 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_800 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_806 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_812 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_333 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_345 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_369 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_376 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_382 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_385 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_392 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_400 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_404 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_443 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_497 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_504 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_510 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_526 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_553 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_559 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_579 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_585 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_595 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_608 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_626 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_638 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_645 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_653 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_659 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_667 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_672 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_685 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_698 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_701 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_713 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_718 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_724 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_727 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_731 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_745 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_761 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_772 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_784 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_790 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_796 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_811 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_818 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_824 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_828 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_356 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_364 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_370 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_378 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_404 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_431 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_453 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_465 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_510 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_516 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_528 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_540 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_544 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_573 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_585 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_605 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_629 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_641 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_647 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_651 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_664 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_673 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_681 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_686 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_709 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_717 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_751 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_762 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_768 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_782 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_796 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_816 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_820 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_823 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_827 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_340 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_374 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_378 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_388 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_399 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_439 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_452 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_458 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_470 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_483 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_487 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_499 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_517 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_549 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_555 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_570 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_582 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_621 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_633 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_641 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_653 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_659 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_683 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_705 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_730 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_736 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_742 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_746 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_752 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_761 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_767 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_773 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_779 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_791 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_797 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_803 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_807 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_810 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_819 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_371 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_380 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_399 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_413 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_420 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_438 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_473 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_491 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_521 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_527 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_539 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_551 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_565 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_609 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_635 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_641 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_652 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_664 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_685 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_693 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_698 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_708 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_714 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_720 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_745 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_751 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_789 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_795 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_801 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_807 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_818 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_369 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_381 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_417 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_440 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_446 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_496 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_511 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_549 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_555 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_563 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_598 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_610 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_618 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_624 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_653 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_665 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_677 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_689 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_697 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_712 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_718 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_724 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_736 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_744 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_754 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_770 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_781 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_787 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_797 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_806 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_817 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_821 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_824 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_390 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_413 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_425 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_446 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_464 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_470 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_482 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_494 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_498 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_517 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_536 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_542 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_551 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_557 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_571 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_582 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_588 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_591 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_595 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_598 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_605 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_621 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_625 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_649 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_661 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_685 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_691 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_711 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_741 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_749 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_752 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_761 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_767 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_794 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_816 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_822 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_831 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_350 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_356 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_383 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_386 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_399 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_441 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_501 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_504 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_512 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_523 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_530 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_546 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_554 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_564 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_606 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_612 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_618 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_630 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_649 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_661 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_665 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_668 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_689 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_695 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_709 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_715 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_773 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_779 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_796 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_811 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_820 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_826 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_355 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_367 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_377 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_398 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_410 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_414 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_443 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_458 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_464 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_470 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_491 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_510 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_524 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_541 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_580 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_592 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_604 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_655 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_671 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_679 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_689 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_703 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_733 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_739 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_751 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_763 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_789 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_795 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_801 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_807 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_819 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_824 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_325 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_342 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_354 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_383 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_408 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_444 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_465 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_486 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_543 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_568 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_580 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_669 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_672 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_676 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_680 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_688 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_705 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_717 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_722 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_728 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_735 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_741 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_751 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_761 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_767 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_773 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_783 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_794 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_800 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_806 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_817 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_823 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_829 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_335 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_342 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_355 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_358 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_370 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_375 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_402 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_408 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_416 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_420 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_426 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_453 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_472 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_478 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_484 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_509 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_523 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_532 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_541 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_547 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_577 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_583 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_595 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_625 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_643 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_649 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_677 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_689 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_715 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_721 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_748 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_754 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_758 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_772 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_778 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_782 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_799 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_820 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_826 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_353 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_360 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_378 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_390 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_396 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_418 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_426 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_432 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_452 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_464 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_538 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_544 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_550 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_562 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_578 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_584 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_594 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_606 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_624 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_632 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_649 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_656 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_669 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_675 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_681 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_713 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_720 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_726 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_734 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_745 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_749 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_766 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_774 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_791 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_797 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_818 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_838 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_345 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_397 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_403 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_415 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_420 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_424 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_427 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_485 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_497 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_521 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_527 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_557 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_566 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_578 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_582 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_592 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_599 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_605 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_611 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_627 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_633 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_641 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_677 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_683 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_691 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_709 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_721 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_735 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_741 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_745 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_762 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_768 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_789 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_381 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_384 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_390 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_396 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_410 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_416 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_427 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_441 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_493 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_514 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_520 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_549 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_553 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_559 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_579 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_585 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_610 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_616 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_628 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_642 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_659 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_669 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_675 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_679 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_689 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_717 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_730 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_740 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_764 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_770 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_778 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_786 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_792 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_817 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_821 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_824 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_415 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_439 ();
 sky130_fd_sc_hd__decap_3 FILLER_85_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_458 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_464 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_476 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_495 ();
 sky130_fd_sc_hd__decap_3 FILLER_85_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_515 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_521 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_527 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_530 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_536 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_540 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_543 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_568 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_574 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_594 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_607 ();
 sky130_fd_sc_hd__decap_3 FILLER_85_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_633 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_643 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_649 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_655 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_661 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_671 ();
 sky130_fd_sc_hd__decap_3 FILLER_85_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_733 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_739 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_751 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_763 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_767 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_773 ();
 sky130_fd_sc_hd__decap_3 FILLER_85_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_800 ();
 sky130_fd_sc_hd__decap_3 FILLER_85_812 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_823 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_333 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_345 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_86_361 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_371 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_374 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_386 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_400 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_407 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_428 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_440 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_474 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_495 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_504 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_510 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_522 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_543 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_555 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_563 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_567 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_575 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_587 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_593 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_610 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_616 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_622 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_649 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_660 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_670 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_674 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_678 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_698 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_713 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_717 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_720 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_733 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_750 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_811 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_819 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_335 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_351 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_357 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_372 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_378 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_382 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_391 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_407 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_423 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_430 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_454 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_472 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_476 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_480 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_486 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_509 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_526 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_532 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_541 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_575 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_581 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_587 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_623 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_644 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_683 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_689 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_699 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_723 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_745 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_751 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_763 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_769 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_799 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_811 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_823 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_827 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_351 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_383 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_395 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_443 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_500 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_509 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_519 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_530 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_541 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_553 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_563 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_575 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_616 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_620 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_633 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_649 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_655 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_659 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_666 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_672 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_684 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_696 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_701 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_709 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_714 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_720 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_736 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_746 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_752 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_766 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_772 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_778 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_782 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_791 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_804 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_810 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_813 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_831 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_835 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_329 ();
 sky130_fd_sc_hd__decap_3 FILLER_89_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_348 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_382 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_429 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_454 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_466 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_478 ();
 sky130_fd_sc_hd__decap_3 FILLER_89_486 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_515 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_521 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_530 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_540 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_571 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_577 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_89_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_630 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_636 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_644 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_652 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_677 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_683 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_693 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_699 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_709 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_715 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_740 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_750 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_761 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_767 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_780 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_794 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_798 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_808 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_815 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_821 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_352 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_375 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_389 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_409 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_425 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_452 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_464 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_495 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_510 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_516 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_549 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_564 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_570 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_576 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_661 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_678 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_682 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_691 ();
 sky130_fd_sc_hd__decap_3 FILLER_90_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_711 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_715 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_721 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_734 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_740 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_746 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_752 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_766 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_772 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_782 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_792 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_335 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_355 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_372 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_378 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_91_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_409 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_427 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_463 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_510 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_527 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_539 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_551 ();
 sky130_fd_sc_hd__decap_3 FILLER_91_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_579 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_671 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_680 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_686 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_692 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_695 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_707 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_719 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_726 ();
 sky130_fd_sc_hd__decap_3 FILLER_91_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_751 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_763 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_794 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_800 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_804 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_814 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_820 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_826 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_836 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_341 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_92_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_370 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_376 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_385 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_394 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_400 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_406 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_435 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_443 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_92_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_462 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_481 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_493 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_525 ();
 sky130_fd_sc_hd__decap_3 FILLER_92_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_537 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_557 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_560 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_593 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_599 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_607 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_610 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_616 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_628 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_632 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_638 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_663 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_666 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_709 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_717 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_732 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_738 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_744 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_750 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_761 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_767 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_779 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_791 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_795 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_798 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_804 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_810 ();
 sky130_fd_sc_hd__decap_3 FILLER_92_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_818 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_824 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_833 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_367 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_370 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_93_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_403 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_412 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_420 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_428 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_438 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_476 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_484 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_529 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_549 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_573 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_592 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_635 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_641 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_649 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_662 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_689 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_695 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_707 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_93_725 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_742 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_746 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_752 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_809 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_812 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_818 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_824 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_345 ();
 sky130_fd_sc_hd__decap_3 FILLER_94_357 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_375 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_383 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_390 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_398 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_419 ();
 sky130_fd_sc_hd__decap_3 FILLER_94_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_428 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_439 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_451 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_459 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_491 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_504 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_510 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_516 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_537 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_545 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_553 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_608 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_619 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_630 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_649 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_670 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_676 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_688 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_708 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_718 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_725 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_755 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_763 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_770 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_776 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_784 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_787 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_799 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_807 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_823 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_829 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_835 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_357 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_370 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_376 ();
 sky130_fd_sc_hd__decap_3 FILLER_95_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_411 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_414 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_420 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_458 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_468 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_480 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_491 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_523 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_527 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_539 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_556 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_576 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_596 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_628 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_637 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_646 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_95_669 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_684 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_690 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_698 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_708 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_737 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_743 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_754 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_760 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_770 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_776 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_794 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_802 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_807 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_828 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_357 ();
 sky130_fd_sc_hd__decap_3 FILLER_96_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_375 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_387 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_394 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_409 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_428 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_434 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_451 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_462 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_482 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_488 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_500 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_514 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_520 ();
 sky130_fd_sc_hd__decap_3 FILLER_96_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_553 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_562 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_568 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_572 ();
 sky130_fd_sc_hd__decap_3 FILLER_96_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_593 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_599 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_607 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_611 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_649 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_655 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_676 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_685 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_699 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_715 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_721 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_727 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_735 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_743 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_755 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_763 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_774 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_786 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_789 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_802 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_808 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_817 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_827 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_835 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_335 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_346 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_356 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_377 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_391 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_423 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_430 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_436 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_442 ();
 sky130_fd_sc_hd__decap_3 FILLER_97_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_454 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_471 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_97_497 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_515 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_519 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_528 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_542 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_546 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_577 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_583 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_593 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_605 ();
 sky130_fd_sc_hd__decap_3 FILLER_97_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_621 ();
 sky130_fd_sc_hd__decap_3 FILLER_97_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_635 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_648 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_654 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_660 ();
 sky130_fd_sc_hd__decap_3 FILLER_97_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_685 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_691 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_703 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_715 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_733 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_739 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_751 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_763 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_783 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_796 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_802 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_812 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_818 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_826 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_321 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_346 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_363 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_379 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_432 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_438 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_441 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_459 ();
 sky130_fd_sc_hd__decap_3 FILLER_98_467 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_499 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_520 ();
 sky130_fd_sc_hd__decap_3 FILLER_98_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_537 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_543 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_551 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_564 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_570 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_574 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_625 ();
 sky130_fd_sc_hd__decap_3 FILLER_98_637 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_649 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_659 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_665 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_671 ();
 sky130_fd_sc_hd__decap_3 FILLER_98_679 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_691 ();
 sky130_fd_sc_hd__decap_3 FILLER_98_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_709 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_721 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_733 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_755 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_767 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_773 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_787 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_795 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_813 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_817 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_823 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_335 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_364 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_370 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_473 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_512 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_518 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_524 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_530 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_536 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_542 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_548 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_554 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_585 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_603 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_611 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_628 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_634 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_647 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_668 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_688 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_694 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_698 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_707 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_737 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_745 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_765 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_776 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_782 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_798 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_804 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_825 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_385 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_394 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_406 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_425 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_437 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_100_473 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_483 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_491 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_515 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_100_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_547 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_560 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_566 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_620 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_632 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_651 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_667 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_670 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_682 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_690 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_719 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_754 ();
 sky130_fd_sc_hd__decap_3 FILLER_100_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_762 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_775 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_795 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_810 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_349 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_391 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_412 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_433 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_459 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_484 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_490 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_529 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_538 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_544 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_584 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_590 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_596 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_602 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_608 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_709 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_715 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_746 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_752 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_766 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_789 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_793 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_796 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_802 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_809 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_815 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_821 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_357 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_360 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_418 ();
 sky130_fd_sc_hd__decap_3 FILLER_102_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_426 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_466 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_494 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_500 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_523 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_549 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_555 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_586 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_607 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_619 ();
 sky130_fd_sc_hd__decap_3 FILLER_102_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_632 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_649 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_661 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_671 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_689 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_711 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_724 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_735 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_741 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_747 ();
 sky130_fd_sc_hd__decap_3 FILLER_102_753 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_765 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_768 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_778 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_790 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_804 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_810 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_819 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_335 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_360 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_371 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_402 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_412 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_420 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_424 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_462 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_471 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_503 ();
 sky130_fd_sc_hd__decap_3 FILLER_103_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_517 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_528 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_542 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_548 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_579 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_595 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_604 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_641 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_647 ();
 sky130_fd_sc_hd__decap_3 FILLER_103_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_681 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_691 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_697 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_703 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_745 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_751 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_763 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_805 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_808 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_814 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_820 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_321 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_369 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_378 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_384 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_387 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_104_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_406 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_441 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_453 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_490 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_496 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_502 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_508 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_539 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_546 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_552 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_567 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_594 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_606 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_612 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_628 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_632 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_649 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_655 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_675 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_698 ();
 sky130_fd_sc_hd__decap_3 FILLER_104_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_707 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_717 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_734 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_740 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_752 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_777 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_787 ();
 sky130_fd_sc_hd__decap_3 FILLER_104_799 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_804 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_810 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_819 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_822 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_348 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_352 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_358 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_364 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_370 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_376 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_380 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_413 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_416 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_422 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_432 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_453 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_478 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_488 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_512 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_524 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_536 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_540 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_546 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_566 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_572 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_576 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_606 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_626 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_636 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_649 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_661 ();
 sky130_fd_sc_hd__decap_3 FILLER_105_669 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_679 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_688 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_694 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_700 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_706 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_712 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_733 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_739 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_742 ();
 sky130_fd_sc_hd__decap_3 FILLER_105_750 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_755 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_761 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_767 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_779 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_796 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_806 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_812 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_818 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_352 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_370 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_382 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_394 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_408 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_431 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_437 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_448 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_472 ();
 sky130_fd_sc_hd__decap_3 FILLER_106_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_482 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_490 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_496 ();
 sky130_fd_sc_hd__decap_3 FILLER_106_504 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_509 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_106_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_538 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_544 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_568 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_587 ();
 sky130_fd_sc_hd__decap_3 FILLER_106_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_594 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_623 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_629 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_645 ();
 sky130_fd_sc_hd__decap_3 FILLER_106_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_662 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_674 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_680 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_690 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_705 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_711 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_717 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_721 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_733 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_737 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_740 ();
 sky130_fd_sc_hd__decap_3 FILLER_106_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_766 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_772 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_784 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_787 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_793 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_797 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_803 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_824 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_833 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_107_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_350 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_359 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_107_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_400 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_406 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_412 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_420 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_426 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_432 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_454 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_460 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_484 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_496 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_536 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_107_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_573 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_628 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_634 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_638 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_641 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_648 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_654 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_660 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_694 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_700 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_706 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_710 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_716 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_722 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_733 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_741 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_744 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_768 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_775 ();
 sky130_fd_sc_hd__decap_3 FILLER_107_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_789 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_795 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_816 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_836 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_108_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_392 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_407 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_425 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_437 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_481 ();
 sky130_fd_sc_hd__decap_8 FILLER_108_487 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_495 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_516 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_530 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_539 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_549 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_555 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_567 ();
 sky130_fd_sc_hd__decap_8 FILLER_108_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_587 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_595 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_619 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_643 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_651 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_658 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_671 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_677 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_683 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_695 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_711 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_717 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_723 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_735 ();
 sky130_fd_sc_hd__decap_8 FILLER_108_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_108_749 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_764 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_770 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_776 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_791 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_797 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_817 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_821 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_831 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_835 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_342 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_354 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_360 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_402 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_409 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_416 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_422 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_428 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_440 ();
 sky130_fd_sc_hd__decap_3 FILLER_109_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_455 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_476 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_482 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_486 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_489 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_510 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_523 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_529 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_538 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_544 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_580 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_598 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_610 ();
 sky130_fd_sc_hd__decap_3 FILLER_109_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_109_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_634 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_654 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_691 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_697 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_745 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_751 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_767 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_778 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_795 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_804 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_810 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_818 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_349 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_386 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_398 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_406 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_450 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_456 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_474 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_497 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_514 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_520 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_540 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_546 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_552 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_560 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_568 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_574 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_580 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_595 ();
 sky130_fd_sc_hd__decap_3 FILLER_110_603 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_608 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_620 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_628 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_632 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_638 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_649 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_653 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_664 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_670 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_676 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_682 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_694 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_713 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_719 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_727 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_731 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_740 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_746 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_761 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_767 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_773 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_781 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_798 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_811 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_819 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_823 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_836 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_369 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_111_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_430 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_456 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_468 ();
 sky130_fd_sc_hd__decap_3 FILLER_111_476 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_485 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_523 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_526 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_536 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_542 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_548 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_554 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_581 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_591 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_604 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_630 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_636 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_642 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_648 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_655 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_661 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_683 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_689 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_695 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_111_725 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_754 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_760 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_768 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_771 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_779 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_795 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_801 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_815 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_818 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_824 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_403 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_409 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_415 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_474 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_488 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_494 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_506 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_510 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_540 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_546 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_552 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_564 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_576 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_626 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_643 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_660 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_675 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_711 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_717 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_723 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_740 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_752 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_761 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_773 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_787 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_795 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_798 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_804 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_810 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_821 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_827 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_835 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_375 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_387 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_400 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_406 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_418 ();
 sky130_fd_sc_hd__decap_3 FILLER_113_426 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_454 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_467 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_480 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_486 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_498 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_528 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_543 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_554 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_579 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_596 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_614 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_624 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_644 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_688 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_700 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_706 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_712 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_737 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_743 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_749 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_761 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_767 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_789 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_801 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_815 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_818 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_824 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_373 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_387 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_397 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_409 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_415 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_438 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_451 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_114_497 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_514 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_520 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_537 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_593 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_605 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_633 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_656 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_660 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_674 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_683 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_689 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_706 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_714 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_722 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_730 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_736 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_742 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_750 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_754 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_768 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_774 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_780 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_783 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_789 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_795 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_801 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_818 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_822 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_826 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_335 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_366 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_378 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_397 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_409 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_415 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_418 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_437 ();
 sky130_fd_sc_hd__decap_8 FILLER_115_440 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_115_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_488 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_521 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_527 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_555 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_588 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_595 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_115_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_643 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_658 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_115_677 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_685 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_699 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_719 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_733 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_739 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_751 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_759 ();
 sky130_fd_sc_hd__decap_8 FILLER_115_765 ();
 sky130_fd_sc_hd__decap_3 FILLER_115_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_795 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_801 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_805 ();
 sky130_fd_sc_hd__decap_8 FILLER_115_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_833 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_333 ();
 sky130_fd_sc_hd__decap_3 FILLER_116_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_351 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_116_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_370 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_382 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_388 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_494 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_500 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_508 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_519 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_531 ();
 sky130_fd_sc_hd__decap_8 FILLER_116_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_541 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_554 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_583 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_616 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_627 ();
 sky130_fd_sc_hd__decap_8 FILLER_116_633 ();
 sky130_fd_sc_hd__decap_3 FILLER_116_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_656 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_662 ();
 sky130_fd_sc_hd__decap_8 FILLER_116_668 ();
 sky130_fd_sc_hd__decap_8 FILLER_116_682 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_705 ();
 sky130_fd_sc_hd__decap_8 FILLER_116_711 ();
 sky130_fd_sc_hd__decap_8 FILLER_116_721 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_731 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_740 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_746 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_752 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_763 ();
 sky130_fd_sc_hd__decap_8 FILLER_116_773 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_781 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_784 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_804 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_813 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_836 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_355 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_368 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_374 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_380 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_117_389 ();
 sky130_fd_sc_hd__decap_3 FILLER_117_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_400 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_422 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_485 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_521 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_532 ();
 sky130_fd_sc_hd__decap_3 FILLER_117_540 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_546 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_568 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_574 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_598 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_635 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_647 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_661 ();
 sky130_fd_sc_hd__decap_3 FILLER_117_669 ();
 sky130_fd_sc_hd__decap_3 FILLER_117_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_678 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_684 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_688 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_700 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_712 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_740 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_746 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_755 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_761 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_767 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_773 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_792 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_798 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_804 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_814 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_827 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_833 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_357 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_387 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_409 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_433 ();
 sky130_fd_sc_hd__decap_8 FILLER_118_439 ();
 sky130_fd_sc_hd__decap_3 FILLER_118_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_452 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_458 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_470 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_496 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_523 ();
 sky130_fd_sc_hd__decap_3 FILLER_118_529 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_559 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_568 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_607 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_610 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_625 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_643 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_651 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_660 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_666 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_678 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_682 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_685 ();
 sky130_fd_sc_hd__decap_3 FILLER_118_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_717 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_721 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_734 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_747 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_775 ();
 sky130_fd_sc_hd__decap_8 FILLER_118_781 ();
 sky130_fd_sc_hd__decap_3 FILLER_118_789 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_794 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_800 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_810 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_820 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_119_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_353 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_367 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_372 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_376 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_398 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_404 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_427 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_430 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_438 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_467 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_479 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_494 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_119_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_523 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_537 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_543 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_558 ();
 sky130_fd_sc_hd__decap_3 FILLER_119_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_584 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_596 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_626 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_632 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_644 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_652 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_677 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_687 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_695 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_707 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_119_725 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_733 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_736 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_746 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_752 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_760 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_764 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_770 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_776 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_789 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_795 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_799 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_802 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_808 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_321 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_355 ();
 sky130_fd_sc_hd__decap_3 FILLER_120_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_374 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_380 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_383 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_396 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_402 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_409 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_428 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_435 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_451 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_501 ();
 sky130_fd_sc_hd__decap_8 FILLER_120_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_521 ();
 sky130_fd_sc_hd__decap_8 FILLER_120_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_548 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_554 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_560 ();
 sky130_fd_sc_hd__decap_3 FILLER_120_572 ();
 sky130_fd_sc_hd__decap_8 FILLER_120_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_120_585 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_595 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_619 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_120_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_670 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_683 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_711 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_717 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_723 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_737 ();
 sky130_fd_sc_hd__decap_8 FILLER_120_743 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_751 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_754 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_767 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_778 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_784 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_794 ();
 sky130_fd_sc_hd__decap_8 FILLER_120_800 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_813 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_821 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_827 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_335 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_343 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_347 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_359 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_371 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_378 ();
 sky130_fd_sc_hd__decap_8 FILLER_121_384 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_400 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_407 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_121_430 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_456 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_462 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_466 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_483 ();
 sky130_fd_sc_hd__decap_3 FILLER_121_495 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_500 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_512 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_522 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_536 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_548 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_573 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_591 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_121_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_625 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_634 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_640 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_652 ();
 sky130_fd_sc_hd__decap_8 FILLER_121_664 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_693 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_700 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_711 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_717 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_745 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_751 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_759 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_789 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_795 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_801 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_816 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_822 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_381 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_396 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_402 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_122_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_122_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_498 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_504 ();
 sky130_fd_sc_hd__decap_8 FILLER_122_516 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_526 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_547 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_565 ();
 sky130_fd_sc_hd__decap_8 FILLER_122_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_122_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_122_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_611 ();
 sky130_fd_sc_hd__decap_3 FILLER_122_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_649 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_661 ();
 sky130_fd_sc_hd__decap_8 FILLER_122_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_681 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_705 ();
 sky130_fd_sc_hd__decap_8 FILLER_122_718 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_732 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_736 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_742 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_748 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_754 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_768 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_779 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_788 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_795 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_808 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_819 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_355 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_358 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_372 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_378 ();
 sky130_fd_sc_hd__decap_8 FILLER_123_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_123_445 ();
 sky130_fd_sc_hd__decap_8 FILLER_123_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_459 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_471 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_483 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_495 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_509 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_521 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_536 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_548 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_123_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_123_625 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_635 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_687 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_694 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_698 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_706 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_123_741 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_768 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_774 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_780 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_800 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_821 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_831 ();
 sky130_fd_sc_hd__decap_3 FILLER_123_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_333 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_374 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_383 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_439 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_457 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_124_481 ();
 sky130_fd_sc_hd__decap_3 FILLER_124_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_495 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_511 ();
 sky130_fd_sc_hd__decap_8 FILLER_124_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_548 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_562 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_594 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_606 ();
 sky130_fd_sc_hd__decap_8 FILLER_124_618 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_124_649 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_124_679 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_689 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_699 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_707 ();
 sky130_fd_sc_hd__decap_8 FILLER_124_716 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_738 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_750 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_761 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_765 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_768 ();
 sky130_fd_sc_hd__decap_8 FILLER_124_781 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_794 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_800 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_823 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_827 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_372 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_376 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_398 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_405 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_411 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_431 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_459 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_465 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_479 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_493 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_519 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_529 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_536 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_547 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_577 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_597 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_603 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_615 ();
 sky130_fd_sc_hd__decap_3 FILLER_125_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_622 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_634 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_646 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_677 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_683 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_694 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_712 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_718 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_724 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_733 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_741 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_745 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_751 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_757 ();
 sky130_fd_sc_hd__decap_3 FILLER_125_765 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_770 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_789 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_795 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_803 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_808 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_812 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_815 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_822 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_349 ();
 sky130_fd_sc_hd__decap_8 FILLER_126_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_126_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_440 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_474 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_497 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_527 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_530 ();
 sky130_fd_sc_hd__decap_3 FILLER_126_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_551 ();
 sky130_fd_sc_hd__decap_8 FILLER_126_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_620 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_633 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_643 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_665 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_672 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_678 ();
 sky130_fd_sc_hd__decap_3 FILLER_126_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_711 ();
 sky130_fd_sc_hd__decap_8 FILLER_126_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_725 ();
 sky130_fd_sc_hd__decap_8 FILLER_126_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_737 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_740 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_764 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_770 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_782 ();
 sky130_fd_sc_hd__decap_3 FILLER_126_794 ();
 sky130_fd_sc_hd__decap_8 FILLER_126_799 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_807 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_361 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_390 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_409 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_422 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_428 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_439 ();
 sky130_fd_sc_hd__decap_3 FILLER_127_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_458 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_464 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_468 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_481 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_127_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_524 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_530 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_534 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_548 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_570 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_579 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_612 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_636 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_648 ();
 sky130_fd_sc_hd__decap_8 FILLER_127_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_685 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_699 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_705 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_711 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_729 ();
 sky130_fd_sc_hd__decap_3 FILLER_127_741 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_746 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_770 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_794 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_798 ();
 sky130_fd_sc_hd__decap_8 FILLER_127_808 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_816 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_128_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_383 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_392 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_398 ();
 sky130_fd_sc_hd__decap_8 FILLER_128_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_415 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_430 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_436 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_461 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_128_486 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_500 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_512 ();
 sky130_fd_sc_hd__decap_8 FILLER_128_515 ();
 sky130_fd_sc_hd__decap_3 FILLER_128_523 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_128_537 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_552 ();
 sky130_fd_sc_hd__decap_8 FILLER_128_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_575 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_625 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_637 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_649 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_661 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_685 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_705 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_717 ();
 sky130_fd_sc_hd__decap_8 FILLER_128_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_737 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_741 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_765 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_771 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_777 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_789 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_795 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_811 ();
 sky130_fd_sc_hd__decap_3 FILLER_128_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_818 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_824 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_379 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_409 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_426 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_439 ();
 sky130_fd_sc_hd__decap_3 FILLER_129_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_456 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_470 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_129_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_509 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_521 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_549 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_552 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_583 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_595 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_607 ();
 sky130_fd_sc_hd__decap_3 FILLER_129_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_621 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_636 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_651 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_655 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_691 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_697 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_703 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_709 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_745 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_749 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_752 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_758 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_771 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_782 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_791 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_804 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_812 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_818 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_824 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_831 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_130_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_130_385 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_401 ();
 sky130_fd_sc_hd__decap_8 FILLER_130_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_415 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_418 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_427 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_430 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_436 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_439 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_445 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_451 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_462 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_484 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_496 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_508 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_520 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_539 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_551 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_557 ();
 sky130_fd_sc_hd__decap_8 FILLER_130_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_584 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_130_598 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_606 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_616 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_620 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_656 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_667 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_687 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_717 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_723 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_737 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_743 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_755 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_763 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_770 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_776 ();
 sky130_fd_sc_hd__decap_8 FILLER_130_782 ();
 sky130_fd_sc_hd__decap_3 FILLER_130_790 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_795 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_808 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_820 ();
 sky130_fd_sc_hd__decap_8 FILLER_130_826 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_131_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_368 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_374 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_400 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_406 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_412 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_415 ();
 sky130_fd_sc_hd__decap_3 FILLER_131_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_435 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_447 ();
 sky130_fd_sc_hd__decap_3 FILLER_131_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_458 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_464 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_476 ();
 sky130_fd_sc_hd__decap_8 FILLER_131_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_510 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_522 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_535 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_548 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_554 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_621 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_628 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_634 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_637 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_663 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_131_677 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_685 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_688 ();
 sky130_fd_sc_hd__decap_8 FILLER_131_696 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_704 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_707 ();
 sky130_fd_sc_hd__decap_8 FILLER_131_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_748 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_754 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_760 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_766 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_778 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_799 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_811 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_814 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_820 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_823 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_357 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_371 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_383 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_392 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_398 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_419 ();
 sky130_fd_sc_hd__decap_3 FILLER_132_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_426 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_432 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_456 ();
 sky130_fd_sc_hd__decap_8 FILLER_132_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_132_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_132_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_550 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_556 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_562 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_568 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_586 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_598 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_607 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_620 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_632 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_132_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_669 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_711 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_717 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_723 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_732 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_744 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_750 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_778 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_784 ();
 sky130_fd_sc_hd__decap_8 FILLER_132_790 ();
 sky130_fd_sc_hd__decap_3 FILLER_132_798 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_813 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_817 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_823 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_373 ();
 sky130_fd_sc_hd__decap_3 FILLER_133_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_415 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_430 ();
 sky130_fd_sc_hd__decap_8 FILLER_133_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_456 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_480 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_509 ();
 sky130_fd_sc_hd__decap_8 FILLER_133_521 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_540 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_546 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_577 ();
 sky130_fd_sc_hd__decap_8 FILLER_133_583 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_605 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_671 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_677 ();
 sky130_fd_sc_hd__decap_8 FILLER_133_680 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_704 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_718 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_724 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_733 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_748 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_754 ();
 sky130_fd_sc_hd__decap_8 FILLER_133_760 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_772 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_778 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_793 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_822 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_831 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_333 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_387 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_134_399 ();
 sky130_fd_sc_hd__decap_3 FILLER_134_407 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_434 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_440 ();
 sky130_fd_sc_hd__decap_8 FILLER_134_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_456 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_462 ();
 sky130_fd_sc_hd__decap_8 FILLER_134_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_134_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_495 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_504 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_564 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_577 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_587 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_603 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_609 ();
 sky130_fd_sc_hd__decap_8 FILLER_134_615 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_626 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_638 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_678 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_684 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_688 ();
 sky130_fd_sc_hd__decap_3 FILLER_134_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_134_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_730 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_736 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_742 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_748 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_754 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_763 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_771 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_777 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_134_795 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_803 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_808 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_819 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_135_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_361 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_372 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_378 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_409 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_415 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_426 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_438 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_135_465 ();
 sky130_fd_sc_hd__decap_8 FILLER_135_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_497 ();
 sky130_fd_sc_hd__decap_3 FILLER_135_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_135_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_527 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_539 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_566 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_578 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_584 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_590 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_596 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_602 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_621 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_631 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_641 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_644 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_650 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_654 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_660 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_683 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_689 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_695 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_710 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_717 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_135_733 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_741 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_744 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_750 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_761 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_767 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_773 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_783 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_798 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_804 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_816 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_820 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_823 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_349 ();
 sky130_fd_sc_hd__decap_8 FILLER_136_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_136_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_378 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_386 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_392 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_398 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_416 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_454 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_466 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_481 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_487 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_499 ();
 sky130_fd_sc_hd__decap_8 FILLER_136_511 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_519 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_531 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_551 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_557 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_563 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_575 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_624 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_649 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_655 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_661 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_669 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_675 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_681 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_688 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_710 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_716 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_722 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_728 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_734 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_742 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_761 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_773 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_781 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_784 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_790 ();
 sky130_fd_sc_hd__decap_8 FILLER_136_803 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_811 ();
 sky130_fd_sc_hd__decap_8 FILLER_136_813 ();
 sky130_fd_sc_hd__decap_3 FILLER_136_821 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_826 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_397 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_401 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_431 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_435 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_469 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_480 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_486 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_503 ();
 sky130_fd_sc_hd__decap_3 FILLER_137_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_573 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_590 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_598 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_606 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_621 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_625 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_642 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_662 ();
 sky130_fd_sc_hd__decap_3 FILLER_137_669 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_685 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_695 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_707 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_738 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_744 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_750 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_756 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_764 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_767 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_783 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_791 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_794 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_798 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_808 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_814 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_820 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_401 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_434 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_440 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_454 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_466 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_481 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_493 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_529 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_559 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_593 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_607 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_613 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_619 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_625 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_634 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_649 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_655 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_666 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_672 ();
 sky130_fd_sc_hd__decap_8 FILLER_138_678 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_686 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_138_705 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_718 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_728 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_737 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_743 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_752 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_761 ();
 sky130_fd_sc_hd__decap_8 FILLER_138_783 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_791 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_813 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_831 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_835 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_349 ();
 sky130_fd_sc_hd__decap_8 FILLER_139_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_369 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_372 ();
 sky130_fd_sc_hd__decap_3 FILLER_139_384 ();
 sky130_fd_sc_hd__decap_3 FILLER_139_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_447 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_458 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_470 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_482 ();
 sky130_fd_sc_hd__decap_8 FILLER_139_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_139_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_527 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_550 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_556 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_583 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_139_595 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_603 ();
 sky130_fd_sc_hd__decap_3 FILLER_139_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_139_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_649 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_662 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_683 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_689 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_695 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_707 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_710 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_716 ();
 sky130_fd_sc_hd__decap_3 FILLER_139_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_736 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_742 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_767 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_773 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_802 ();
 sky130_fd_sc_hd__decap_8 FILLER_139_814 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_824 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_140_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_353 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_362 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_374 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_378 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_381 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_387 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_399 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_140_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_445 ();
 sky130_fd_sc_hd__decap_3 FILLER_140_457 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_484 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_496 ();
 sky130_fd_sc_hd__decap_8 FILLER_140_508 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_516 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_140_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_555 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_573 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_587 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_600 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_604 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_614 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_620 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_626 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_632 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_638 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_651 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_661 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_667 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_677 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_683 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_695 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_698 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_707 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_716 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_722 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_728 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_738 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_744 ();
 sky130_fd_sc_hd__decap_8 FILLER_140_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_765 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_776 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_782 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_794 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_806 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_819 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_827 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_353 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_359 ();
 sky130_fd_sc_hd__decap_8 FILLER_141_370 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_378 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_407 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_413 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_439 ();
 sky130_fd_sc_hd__decap_3 FILLER_141_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_141_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_485 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_492 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_512 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_536 ();
 sky130_fd_sc_hd__decap_8 FILLER_141_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_567 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_577 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_583 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_604 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_621 ();
 sky130_fd_sc_hd__decap_8 FILLER_141_627 ();
 sky130_fd_sc_hd__decap_3 FILLER_141_635 ();
 sky130_fd_sc_hd__decap_8 FILLER_141_640 ();
 sky130_fd_sc_hd__decap_3 FILLER_141_648 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_654 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_660 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_689 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_695 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_703 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_735 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_747 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_759 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_763 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_780 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_809 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_812 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_818 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_383 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_395 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_407 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_419 ();
 sky130_fd_sc_hd__decap_3 FILLER_142_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_427 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_440 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_452 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_458 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_482 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_486 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_496 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_508 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_514 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_518 ();
 sky130_fd_sc_hd__decap_3 FILLER_142_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_142_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_566 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_605 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_611 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_628 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_634 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_640 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_649 ();
 sky130_fd_sc_hd__decap_8 FILLER_142_666 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_683 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_687 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_691 ();
 sky130_fd_sc_hd__decap_3 FILLER_142_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_710 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_716 ();
 sky130_fd_sc_hd__decap_8 FILLER_142_722 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_730 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_734 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_740 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_752 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_763 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_766 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_772 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_786 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_792 ();
 sky130_fd_sc_hd__decap_8 FILLER_142_798 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_806 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_831 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_835 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_356 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_362 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_366 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_378 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_399 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_143_408 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_416 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_424 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_431 ();
 sky130_fd_sc_hd__decap_3 FILLER_143_445 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_460 ();
 sky130_fd_sc_hd__decap_8 FILLER_143_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_482 ();
 sky130_fd_sc_hd__decap_8 FILLER_143_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_143_511 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_535 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_575 ();
 sky130_fd_sc_hd__decap_8 FILLER_143_587 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_604 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_638 ();
 sky130_fd_sc_hd__decap_8 FILLER_143_644 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_652 ();
 sky130_fd_sc_hd__decap_8 FILLER_143_656 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_664 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_668 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_695 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_708 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_715 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_727 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_740 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_744 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_764 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_770 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_776 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_789 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_793 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_803 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_809 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_822 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_333 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_351 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_144_374 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_382 ();
 sky130_fd_sc_hd__decap_8 FILLER_144_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_397 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_430 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_436 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_457 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_509 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_530 ();
 sky130_fd_sc_hd__decap_8 FILLER_144_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_541 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_551 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_567 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_582 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_144_607 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_623 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_635 ();
 sky130_fd_sc_hd__decap_3 FILLER_144_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_661 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_680 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_706 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_712 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_718 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_722 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_725 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_732 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_743 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_750 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_763 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_771 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_782 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_793 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_808 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_817 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_821 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_824 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_828 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_832 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_836 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_145_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_367 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_370 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_397 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_403 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_406 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_414 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_426 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_435 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_467 ();
 sky130_fd_sc_hd__decap_8 FILLER_145_478 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_522 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_532 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_536 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_543 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_145_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_145_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_595 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_606 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_627 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_633 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_646 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_652 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_670 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_145_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_693 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_697 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_709 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_712 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_726 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_742 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_748 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_754 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_760 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_772 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_778 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_145_791 ();
 sky130_fd_sc_hd__decap_8 FILLER_145_815 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_831 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_333 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_345 ();
 sky130_fd_sc_hd__decap_8 FILLER_146_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_380 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_398 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_428 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_434 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_443 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_455 ();
 sky130_fd_sc_hd__decap_8 FILLER_146_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_552 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_564 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_576 ();
 sky130_fd_sc_hd__decap_8 FILLER_146_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_603 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_609 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_633 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_699 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_707 ();
 sky130_fd_sc_hd__decap_8 FILLER_146_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_745 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_755 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_772 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_778 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_784 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_787 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_793 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_796 ();
 sky130_fd_sc_hd__decap_8 FILLER_146_803 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_827 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_833 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_391 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_412 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_424 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_430 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_436 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_541 ();
 sky130_fd_sc_hd__decap_3 FILLER_147_553 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_579 ();
 sky130_fd_sc_hd__decap_8 FILLER_147_591 ();
 sky130_fd_sc_hd__decap_3 FILLER_147_599 ();
 sky130_fd_sc_hd__decap_8 FILLER_147_604 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_636 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_648 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_660 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_677 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_683 ();
 sky130_fd_sc_hd__decap_3 FILLER_147_695 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_700 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_706 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_765 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_780 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_809 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_821 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_827 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_148_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_394 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_400 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_412 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_416 ();
 sky130_fd_sc_hd__decap_3 FILLER_148_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_426 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_450 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_455 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_148_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_483 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_553 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_559 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_565 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_586 ();
 sky130_fd_sc_hd__decap_8 FILLER_148_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_611 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_148_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_663 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_669 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_675 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_681 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_698 ();
 sky130_fd_sc_hd__decap_3 FILLER_148_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_712 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_718 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_730 ();
 sky130_fd_sc_hd__decap_8 FILLER_148_742 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_750 ();
 sky130_fd_sc_hd__decap_3 FILLER_148_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_778 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_790 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_794 ();
 sky130_fd_sc_hd__decap_8 FILLER_148_801 ();
 sky130_fd_sc_hd__decap_3 FILLER_148_809 ();
 sky130_fd_sc_hd__decap_8 FILLER_148_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_821 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_824 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_830 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_367 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_370 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_409 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_415 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_425 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_470 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_476 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_500 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_521 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_527 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_537 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_548 ();
 sky130_fd_sc_hd__decap_3 FILLER_149_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_570 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_576 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_580 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_610 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_639 ();
 sky130_fd_sc_hd__decap_8 FILLER_149_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_653 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_656 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_679 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_691 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_697 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_703 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_709 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_715 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_741 ();
 sky130_fd_sc_hd__decap_8 FILLER_149_747 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_758 ();
 sky130_fd_sc_hd__decap_8 FILLER_149_764 ();
 sky130_fd_sc_hd__decap_3 FILLER_149_772 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_782 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_803 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_806 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_821 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_345 ();
 sky130_fd_sc_hd__decap_3 FILLER_150_357 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_410 ();
 sky130_fd_sc_hd__decap_3 FILLER_150_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_425 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_437 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_481 ();
 sky130_fd_sc_hd__decap_8 FILLER_150_493 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_501 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_504 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_510 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_518 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_554 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_571 ();
 sky130_fd_sc_hd__decap_8 FILLER_150_580 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_606 ();
 sky130_fd_sc_hd__decap_8 FILLER_150_612 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_633 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_637 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_640 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_651 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_665 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_675 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_705 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_709 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_732 ();
 sky130_fd_sc_hd__decap_8 FILLER_150_738 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_746 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_755 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_761 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_770 ();
 sky130_fd_sc_hd__decap_8 FILLER_150_776 ();
 sky130_fd_sc_hd__decap_3 FILLER_150_784 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_789 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_801 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_807 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_810 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_828 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_151_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_355 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_366 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_397 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_403 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_412 ();
 sky130_fd_sc_hd__decap_8 FILLER_151_424 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_462 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_474 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_486 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_494 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_500 ();
 sky130_fd_sc_hd__decap_3 FILLER_151_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_528 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_532 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_548 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_567 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_607 ();
 sky130_fd_sc_hd__decap_3 FILLER_151_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_621 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_633 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_636 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_647 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_653 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_659 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_663 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_681 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_691 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_715 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_743 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_754 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_760 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_766 ();
 sky130_fd_sc_hd__decap_8 FILLER_151_772 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_782 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_798 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_802 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_805 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_811 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_817 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_821 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_372 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_378 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_381 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_387 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_397 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_403 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_415 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_433 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_453 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_459 ();
 sky130_fd_sc_hd__decap_8 FILLER_152_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_498 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_507 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_518 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_548 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_557 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_575 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_593 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_605 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_608 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_614 ();
 sky130_fd_sc_hd__decap_8 FILLER_152_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_625 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_628 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_654 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_660 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_664 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_667 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_679 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_711 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_717 ();
 sky130_fd_sc_hd__decap_8 FILLER_152_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_731 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_741 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_747 ();
 sky130_fd_sc_hd__decap_3 FILLER_152_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_761 ();
 sky130_fd_sc_hd__decap_8 FILLER_152_773 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_781 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_784 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_790 ();
 sky130_fd_sc_hd__decap_8 FILLER_152_799 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_807 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_824 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_366 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_379 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_416 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_153_454 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_462 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_469 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_502 ();
 sky130_fd_sc_hd__decap_3 FILLER_153_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_530 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_539 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_551 ();
 sky130_fd_sc_hd__decap_3 FILLER_153_557 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_577 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_584 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_590 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_594 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_607 ();
 sky130_fd_sc_hd__decap_3 FILLER_153_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_627 ();
 sky130_fd_sc_hd__decap_8 FILLER_153_633 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_641 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_649 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_683 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_689 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_695 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_707 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_723 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_153_738 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_750 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_756 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_762 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_768 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_774 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_780 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_791 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_801 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_814 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_820 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_824 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_827 ();
 sky130_fd_sc_hd__decap_3 FILLER_153_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_154_345 ();
 sky130_fd_sc_hd__decap_8 FILLER_154_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_383 ();
 sky130_fd_sc_hd__decap_8 FILLER_154_395 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_407 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_435 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_444 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_456 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_487 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_491 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_500 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_506 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_543 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_549 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_557 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_586 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_602 ();
 sky130_fd_sc_hd__decap_8 FILLER_154_608 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_616 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_624 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_632 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_654 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_660 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_666 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_672 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_678 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_684 ();
 sky130_fd_sc_hd__decap_8 FILLER_154_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_705 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_717 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_731 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_737 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_740 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_746 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_752 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_771 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_782 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_788 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_824 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_373 ();
 sky130_fd_sc_hd__decap_3 FILLER_155_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_390 ();
 sky130_fd_sc_hd__decap_8 FILLER_155_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_155_406 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_414 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_155_431 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_459 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_465 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_495 ();
 sky130_fd_sc_hd__decap_3 FILLER_155_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_512 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_518 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_524 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_530 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_536 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_542 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_548 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_554 ();
 sky130_fd_sc_hd__decap_3 FILLER_155_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_578 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_590 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_605 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_626 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_641 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_649 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_655 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_661 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_683 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_689 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_713 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_741 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_747 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_753 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_761 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_765 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_790 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_796 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_806 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_810 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_155_826 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_381 ();
 sky130_fd_sc_hd__decap_8 FILLER_156_388 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_418 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_430 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_436 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_442 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_448 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_454 ();
 sky130_fd_sc_hd__decap_8 FILLER_156_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_499 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_511 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_156_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_551 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_557 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_563 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_571 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_577 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_586 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_605 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_649 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_655 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_661 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_667 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_679 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_685 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_689 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_705 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_709 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_712 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_719 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_726 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_732 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_740 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_752 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_761 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_772 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_781 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_787 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_791 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_794 ();
 sky130_fd_sc_hd__decap_8 FILLER_156_800 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_810 ();
 sky130_fd_sc_hd__decap_3 FILLER_156_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_818 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_824 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_390 ();
 sky130_fd_sc_hd__decap_3 FILLER_157_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_410 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_416 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_420 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_423 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_157_529 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_534 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_554 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_157_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_578 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_584 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_596 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_602 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_640 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_646 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_652 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_658 ();
 sky130_fd_sc_hd__decap_8 FILLER_157_664 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_680 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_690 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_696 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_702 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_708 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_733 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_745 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_770 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_776 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_157_792 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_806 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_812 ();
 sky130_fd_sc_hd__decap_8 FILLER_157_815 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_385 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_411 ();
 sky130_fd_sc_hd__decap_3 FILLER_158_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_425 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_437 ();
 sky130_fd_sc_hd__decap_8 FILLER_158_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_464 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_470 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_492 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_498 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_510 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_522 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_551 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_557 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_569 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_575 ();
 sky130_fd_sc_hd__decap_8 FILLER_158_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_607 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_613 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_619 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_625 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_631 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_649 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_655 ();
 sky130_fd_sc_hd__decap_8 FILLER_158_667 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_675 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_679 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_710 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_721 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_732 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_741 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_747 ();
 sky130_fd_sc_hd__decap_3 FILLER_158_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_761 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_767 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_773 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_781 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_824 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_828 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_159_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_159_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_406 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_412 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_433 ();
 sky130_fd_sc_hd__decap_8 FILLER_159_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_509 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_542 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_548 ();
 sky130_fd_sc_hd__decap_3 FILLER_159_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_578 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_584 ();
 sky130_fd_sc_hd__decap_8 FILLER_159_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_603 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_633 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_639 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_651 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_663 ();
 sky130_fd_sc_hd__decap_3 FILLER_159_669 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_695 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_708 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_745 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_751 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_763 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_767 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_770 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_776 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_794 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_800 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_806 ();
 sky130_fd_sc_hd__decap_8 FILLER_159_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_821 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_824 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_831 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_160_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_435 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_453 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_160_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_490 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_510 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_522 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_542 ();
 sky130_fd_sc_hd__decap_8 FILLER_160_548 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_556 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_559 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_571 ();
 sky130_fd_sc_hd__decap_8 FILLER_160_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_160_585 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_595 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_610 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_616 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_622 ();
 sky130_fd_sc_hd__decap_8 FILLER_160_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_642 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_649 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_667 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_679 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_689 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_699 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_707 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_719 ();
 sky130_fd_sc_hd__decap_8 FILLER_160_725 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_736 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_745 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_752 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_757 ();
 sky130_fd_sc_hd__decap_3 FILLER_160_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_774 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_780 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_792 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_798 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_802 ();
 sky130_fd_sc_hd__decap_3 FILLER_160_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_813 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_821 ();
 sky130_fd_sc_hd__decap_3 FILLER_160_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_411 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_414 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_424 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_430 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_434 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_446 ();
 sky130_fd_sc_hd__decap_8 FILLER_161_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_465 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_471 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_502 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_520 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_549 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_577 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_583 ();
 sky130_fd_sc_hd__decap_8 FILLER_161_594 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_633 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_637 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_640 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_661 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_667 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_695 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_707 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_710 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_716 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_722 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_738 ();
 sky130_fd_sc_hd__decap_8 FILLER_161_744 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_771 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_803 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_823 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_418 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_438 ();
 sky130_fd_sc_hd__decap_8 FILLER_162_444 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_452 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_459 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_162_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_488 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_494 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_521 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_540 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_553 ();
 sky130_fd_sc_hd__decap_8 FILLER_162_563 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_578 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_608 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_614 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_620 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_626 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_632 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_652 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_658 ();
 sky130_fd_sc_hd__decap_8 FILLER_162_680 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_688 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_691 ();
 sky130_fd_sc_hd__decap_3 FILLER_162_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_162_721 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_733 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_737 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_740 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_752 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_769 ();
 sky130_fd_sc_hd__decap_8 FILLER_162_781 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_791 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_797 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_803 ();
 sky130_fd_sc_hd__decap_3 FILLER_162_809 ();
 sky130_fd_sc_hd__decap_3 FILLER_162_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_819 ();
 sky130_fd_sc_hd__decap_3 FILLER_162_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_391 ();
 sky130_fd_sc_hd__decap_3 FILLER_163_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_398 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_410 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_422 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_446 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_459 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_465 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_163_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_515 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_521 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_535 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_582 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_588 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_594 ();
 sky130_fd_sc_hd__decap_8 FILLER_163_600 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_628 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_632 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_635 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_647 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_659 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_671 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_679 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_682 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_688 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_700 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_712 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_724 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_735 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_764 ();
 sky130_fd_sc_hd__decap_8 FILLER_163_776 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_797 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_805 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_811 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_823 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_164_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_394 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_400 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_432 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_436 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_444 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_450 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_456 ();
 sky130_fd_sc_hd__decap_8 FILLER_164_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_531 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_539 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_542 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_553 ();
 sky130_fd_sc_hd__decap_8 FILLER_164_559 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_579 ();
 sky130_fd_sc_hd__decap_3 FILLER_164_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_605 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_630 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_643 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_651 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_654 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_660 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_666 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_680 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_686 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_711 ();
 sky130_fd_sc_hd__decap_8 FILLER_164_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_725 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_728 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_734 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_739 ();
 sky130_fd_sc_hd__decap_8 FILLER_164_745 ();
 sky130_fd_sc_hd__decap_3 FILLER_164_753 ();
 sky130_fd_sc_hd__decap_8 FILLER_164_757 ();
 sky130_fd_sc_hd__decap_3 FILLER_164_765 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_771 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_783 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_795 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_798 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_804 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_810 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_820 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_826 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_165_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_381 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_390 ();
 sky130_fd_sc_hd__decap_3 FILLER_165_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_438 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_453 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_487 ();
 sky130_fd_sc_hd__decap_8 FILLER_165_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_165_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_165_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_527 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_539 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_542 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_558 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_572 ();
 sky130_fd_sc_hd__decap_8 FILLER_165_578 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_588 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_603 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_165_628 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_636 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_642 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_648 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_654 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_165_678 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_686 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_693 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_699 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_726 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_741 ();
 sky130_fd_sc_hd__decap_8 FILLER_165_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_755 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_758 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_764 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_775 ();
 sky130_fd_sc_hd__decap_3 FILLER_165_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_789 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_795 ();
 sky130_fd_sc_hd__decap_8 FILLER_165_801 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_809 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_812 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_818 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_824 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_383 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_386 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_392 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_442 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_453 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_493 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_499 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_511 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_517 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_540 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_546 ();
 sky130_fd_sc_hd__decap_8 FILLER_166_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_560 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_564 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_586 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_593 ();
 sky130_fd_sc_hd__decap_8 FILLER_166_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_609 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_623 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_629 ();
 sky130_fd_sc_hd__decap_8 FILLER_166_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_643 ();
 sky130_fd_sc_hd__decap_8 FILLER_166_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_659 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_665 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_668 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_674 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_684 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_718 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_728 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_734 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_740 ();
 sky130_fd_sc_hd__decap_8 FILLER_166_746 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_754 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_777 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_788 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_794 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_800 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_166_817 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_825 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_373 ();
 sky130_fd_sc_hd__decap_3 FILLER_167_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_411 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_417 ();
 sky130_fd_sc_hd__decap_8 FILLER_167_423 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_453 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_482 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_494 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_509 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_518 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_522 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_544 ();
 sky130_fd_sc_hd__decap_8 FILLER_167_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_558 ();
 sky130_fd_sc_hd__decap_8 FILLER_167_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_167_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_574 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_625 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_631 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_637 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_643 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_647 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_654 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_681 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_687 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_707 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_718 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_724 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_735 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_747 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_759 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_765 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_774 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_780 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_795 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_801 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_814 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_820 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_168_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_168_385 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_409 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_439 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_457 ();
 sky130_fd_sc_hd__decap_3 FILLER_168_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_507 ();
 sky130_fd_sc_hd__decap_8 FILLER_168_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_168_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_537 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_543 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_555 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_558 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_564 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_584 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_595 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_602 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_635 ();
 sky130_fd_sc_hd__decap_3 FILLER_168_641 ();
 sky130_fd_sc_hd__decap_8 FILLER_168_645 ();
 sky130_fd_sc_hd__decap_3 FILLER_168_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_658 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_666 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_672 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_678 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_684 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_705 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_711 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_717 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_721 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_730 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_746 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_752 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_775 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_795 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_801 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_824 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_412 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_433 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_467 ();
 sky130_fd_sc_hd__decap_8 FILLER_169_484 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_492 ();
 sky130_fd_sc_hd__decap_3 FILLER_169_501 ();
 sky130_fd_sc_hd__decap_3 FILLER_169_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_169_516 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_524 ();
 sky130_fd_sc_hd__decap_8 FILLER_169_542 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_550 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_556 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_572 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_578 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_591 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_606 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_624 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_630 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_636 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_642 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_648 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_654 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_666 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_680 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_686 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_692 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_698 ();
 sky130_fd_sc_hd__decap_8 FILLER_169_710 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_720 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_745 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_751 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_763 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_779 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_794 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_800 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_411 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_484 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_490 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_494 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_500 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_170_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_559 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_577 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_587 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_595 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_605 ();
 sky130_fd_sc_hd__decap_8 FILLER_170_611 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_633 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_642 ();
 sky130_fd_sc_hd__decap_3 FILLER_170_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_667 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_686 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_698 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_170_713 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_734 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_740 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_781 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_787 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_791 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_794 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_804 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_170_818 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_171_405 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_415 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_423 ();
 sky130_fd_sc_hd__decap_8 FILLER_171_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_443 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_468 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_480 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_486 ();
 sky130_fd_sc_hd__decap_8 FILLER_171_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_515 ();
 sky130_fd_sc_hd__decap_8 FILLER_171_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_559 ();
 sky130_fd_sc_hd__decap_3 FILLER_171_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_581 ();
 sky130_fd_sc_hd__decap_8 FILLER_171_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_595 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_603 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_171_621 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_631 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_691 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_709 ();
 sky130_fd_sc_hd__decap_3 FILLER_171_721 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_733 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_737 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_764 ();
 sky130_fd_sc_hd__decap_8 FILLER_171_776 ();
 sky130_fd_sc_hd__decap_8 FILLER_171_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_795 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_801 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_807 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_819 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_823 ();
 sky130_fd_sc_hd__decap_8 FILLER_171_826 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_389 ();
 sky130_fd_sc_hd__decap_8 FILLER_172_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_428 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_434 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_458 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_485 ();
 sky130_fd_sc_hd__decap_8 FILLER_172_488 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_496 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_508 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_512 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_531 ();
 sky130_fd_sc_hd__decap_3 FILLER_172_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_172_538 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_546 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_549 ();
 sky130_fd_sc_hd__decap_8 FILLER_172_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_563 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_607 ();
 sky130_fd_sc_hd__decap_8 FILLER_172_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_172_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_655 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_661 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_667 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_679 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_705 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_717 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_731 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_737 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_748 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_172_761 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_771 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_783 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_789 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_792 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_798 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_804 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_810 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_819 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_826 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_833 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_173_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_173_413 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_479 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_509 ();
 sky130_fd_sc_hd__decap_8 FILLER_173_515 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_523 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_532 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_538 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_550 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_554 ();
 sky130_fd_sc_hd__decap_3 FILLER_173_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_581 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_593 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_605 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_611 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_614 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_621 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_638 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_644 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_647 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_651 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_661 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_685 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_700 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_719 ();
 sky130_fd_sc_hd__decap_3 FILLER_173_725 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_743 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_755 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_759 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_764 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_770 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_776 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_173_789 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_797 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_800 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_806 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_812 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_818 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_824 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_408 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_425 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_437 ();
 sky130_fd_sc_hd__decap_8 FILLER_174_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_174_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_174_511 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_519 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_552 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_564 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_576 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_593 ();
 sky130_fd_sc_hd__decap_8 FILLER_174_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_626 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_632 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_649 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_655 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_667 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_671 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_683 ();
 sky130_fd_sc_hd__decap_8 FILLER_174_689 ();
 sky130_fd_sc_hd__decap_3 FILLER_174_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_705 ();
 sky130_fd_sc_hd__decap_3 FILLER_174_717 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_722 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_728 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_734 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_740 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_743 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_752 ();
 sky130_fd_sc_hd__decap_3 FILLER_174_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_767 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_778 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_791 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_797 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_803 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_807 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_810 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_820 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_409 ();
 sky130_fd_sc_hd__decap_8 FILLER_175_418 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_426 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_453 ();
 sky130_fd_sc_hd__decap_3 FILLER_175_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_473 ();
 sky130_fd_sc_hd__decap_8 FILLER_175_479 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_175_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_175_509 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_526 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_532 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_546 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_565 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_607 ();
 sky130_fd_sc_hd__decap_3 FILLER_175_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_633 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_175_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_175_665 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_683 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_689 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_695 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_707 ();
 sky130_fd_sc_hd__decap_8 FILLER_175_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_175_736 ();
 sky130_fd_sc_hd__decap_8 FILLER_175_752 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_768 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_778 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_789 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_799 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_809 ();
 sky130_fd_sc_hd__decap_8 FILLER_175_812 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_822 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_839 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_389 ();
 sky130_fd_sc_hd__decap_8 FILLER_176_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_409 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_431 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_454 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_176_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_497 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_506 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_520 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_526 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_546 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_566 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_572 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_599 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_605 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_611 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_176_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_669 ();
 sky130_fd_sc_hd__decap_8 FILLER_176_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_689 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_723 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_731 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_742 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_748 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_761 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_767 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_773 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_790 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_810 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_819 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_824 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_391 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_402 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_408 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_414 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_423 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_435 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_503 ();
 sky130_fd_sc_hd__decap_3 FILLER_177_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_522 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_528 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_534 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_540 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_548 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_577 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_587 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_593 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_599 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_636 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_642 ();
 sky130_fd_sc_hd__decap_8 FILLER_177_648 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_660 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_691 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_697 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_703 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_709 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_721 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_724 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_734 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_740 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_746 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_752 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_758 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_764 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_776 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_793 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_806 ();
 sky130_fd_sc_hd__decap_8 FILLER_177_819 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_827 ();
 sky130_fd_sc_hd__decap_3 FILLER_177_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_414 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_438 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_456 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_463 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_495 ();
 sky130_fd_sc_hd__decap_8 FILLER_178_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_512 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_518 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_178_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_178_570 ();
 sky130_fd_sc_hd__decap_3 FILLER_178_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_589 ();
 sky130_fd_sc_hd__decap_3 FILLER_178_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_606 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_632 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_649 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_653 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_660 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_672 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_684 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_705 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_717 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_742 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_748 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_763 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_772 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_778 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_784 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_790 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_796 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_802 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_808 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_824 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_828 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_838 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_409 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_412 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_426 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_430 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_179_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_467 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_486 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_495 ();
 sky130_fd_sc_hd__decap_3 FILLER_179_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_515 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_521 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_581 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_587 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_591 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_606 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_641 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_670 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_744 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_756 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_768 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_771 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_783 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_789 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_792 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_798 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_804 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_823 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_827 ();
 sky130_fd_sc_hd__decap_3 FILLER_179_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_413 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_180_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_484 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_490 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_496 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_514 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_542 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_548 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_560 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_564 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_567 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_619 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_633 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_639 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_649 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_661 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_681 ();
 sky130_fd_sc_hd__decap_8 FILLER_180_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_695 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_180_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_717 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_722 ();
 sky130_fd_sc_hd__decap_8 FILLER_180_734 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_742 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_746 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_752 ();
 sky130_fd_sc_hd__decap_8 FILLER_180_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_765 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_768 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_788 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_794 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_802 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_808 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_817 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_821 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_826 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_836 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_447 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_464 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_484 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_490 ();
 sky130_fd_sc_hd__decap_8 FILLER_181_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_521 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_525 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_528 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_532 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_535 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_547 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_577 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_588 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_597 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_603 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_615 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_181_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_639 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_651 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_181_669 ();
 sky130_fd_sc_hd__decap_8 FILLER_181_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_681 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_692 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_698 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_704 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_710 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_716 ();
 sky130_fd_sc_hd__decap_8 FILLER_181_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_737 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_740 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_744 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_747 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_753 ();
 sky130_fd_sc_hd__decap_8 FILLER_181_759 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_767 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_770 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_792 ();
 sky130_fd_sc_hd__decap_8 FILLER_181_798 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_806 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_809 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_815 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_821 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_825 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_828 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_459 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_463 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_466 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_470 ();
 sky130_fd_sc_hd__decap_3 FILLER_182_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_499 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_508 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_514 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_520 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_542 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_548 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_554 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_560 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_566 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_572 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_576 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_579 ();
 sky130_fd_sc_hd__decap_3 FILLER_182_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_593 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_605 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_655 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_661 ();
 sky130_fd_sc_hd__decap_8 FILLER_182_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_675 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_678 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_685 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_710 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_716 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_722 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_728 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_734 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_740 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_746 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_761 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_767 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_773 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_784 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_790 ();
 sky130_fd_sc_hd__decap_8 FILLER_182_796 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_804 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_808 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_818 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_183_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_183_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_515 ();
 sky130_fd_sc_hd__decap_8 FILLER_183_526 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_534 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_570 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_576 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_582 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_588 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_594 ();
 sky130_fd_sc_hd__decap_8 FILLER_183_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_614 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_628 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_634 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_638 ();
 sky130_fd_sc_hd__decap_8 FILLER_183_641 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_677 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_683 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_686 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_693 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_738 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_749 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_761 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_767 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_773 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_777 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_782 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_791 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_808 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_814 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_827 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_833 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_445 ();
 sky130_fd_sc_hd__decap_8 FILLER_184_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_523 ();
 sky130_fd_sc_hd__decap_3 FILLER_184_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_553 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_562 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_566 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_593 ();
 sky130_fd_sc_hd__decap_3 FILLER_184_605 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_610 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_622 ();
 sky130_fd_sc_hd__decap_8 FILLER_184_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_669 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_683 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_687 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_690 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_719 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_725 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_762 ();
 sky130_fd_sc_hd__decap_8 FILLER_184_768 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_778 ();
 sky130_fd_sc_hd__decap_8 FILLER_184_786 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_810 ();
 sky130_fd_sc_hd__decap_3 FILLER_184_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_184_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_833 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_838 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_185_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_469 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_472 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_481 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_487 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_509 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_521 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_532 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_538 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_558 ();
 sky130_fd_sc_hd__decap_3 FILLER_185_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_577 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_583 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_595 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_606 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_627 ();
 sky130_fd_sc_hd__decap_3 FILLER_185_639 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_644 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_656 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_684 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_690 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_696 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_702 ();
 sky130_fd_sc_hd__decap_8 FILLER_185_708 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_716 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_719 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_751 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_762 ();
 sky130_fd_sc_hd__decap_8 FILLER_185_771 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_779 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_782 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_791 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_794 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_814 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_834 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_186_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_463 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_481 ();
 sky130_fd_sc_hd__decap_8 FILLER_186_487 ();
 sky130_fd_sc_hd__decap_3 FILLER_186_495 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_500 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_504 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_507 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_540 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_554 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_568 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_593 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_622 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_628 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_634 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_649 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_661 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_683 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_689 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_186_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_721 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_725 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_731 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_737 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_743 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_757 ();
 sky130_fd_sc_hd__decap_3 FILLER_186_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_774 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_780 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_786 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_792 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_798 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_804 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_810 ();
 sky130_fd_sc_hd__decap_3 FILLER_186_813 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_836 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_447 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_463 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_469 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_503 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_519 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_530 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_536 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_542 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_548 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_583 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_594 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_614 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_640 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_652 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_670 ();
 sky130_fd_sc_hd__decap_8 FILLER_187_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_681 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_685 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_691 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_703 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_734 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_740 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_744 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_753 ();
 sky130_fd_sc_hd__decap_8 FILLER_187_759 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_767 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_770 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_789 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_795 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_798 ();
 sky130_fd_sc_hd__decap_8 FILLER_187_808 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_816 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_820 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_839 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_462 ();
 sky130_fd_sc_hd__decap_8 FILLER_188_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_519 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_549 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_555 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_566 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_577 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_587 ();
 sky130_fd_sc_hd__decap_3 FILLER_188_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_611 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_643 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_649 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_675 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_687 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_719 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_725 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_737 ();
 sky130_fd_sc_hd__decap_8 FILLER_188_745 ();
 sky130_fd_sc_hd__decap_3 FILLER_188_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_768 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_788 ();
 sky130_fd_sc_hd__decap_8 FILLER_188_794 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_804 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_810 ();
 sky130_fd_sc_hd__decap_3 FILLER_188_813 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_818 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_489 ();
 sky130_fd_sc_hd__decap_8 FILLER_189_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_523 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_529 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_535 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_553 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_580 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_586 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_592 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_598 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_604 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_610 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_626 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_632 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_638 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_647 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_659 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_671 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_679 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_682 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_689 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_189_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_741 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_753 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_756 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_762 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_770 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_776 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_789 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_801 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_805 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_811 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_818 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_499 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_521 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_190_541 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_551 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_557 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_563 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_575 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_593 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_599 ();
 sky130_fd_sc_hd__decap_8 FILLER_190_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_626 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_632 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_649 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_655 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_667 ();
 sky130_fd_sc_hd__decap_3 FILLER_190_679 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_684 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_688 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_691 ();
 sky130_fd_sc_hd__decap_3 FILLER_190_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_705 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_711 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_719 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_730 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_736 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_742 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_766 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_772 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_791 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_795 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_798 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_804 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_810 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_820 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_824 ();
 sky130_fd_sc_hd__decap_8 FILLER_190_828 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_191_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_480 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_486 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_492 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_496 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_509 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_516 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_522 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_528 ();
 sky130_fd_sc_hd__decap_8 FILLER_191_538 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_546 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_191_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_579 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_585 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_591 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_597 ();
 sky130_fd_sc_hd__decap_3 FILLER_191_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_614 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_640 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_652 ();
 sky130_fd_sc_hd__decap_8 FILLER_191_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_682 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_689 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_695 ();
 sky130_fd_sc_hd__decap_8 FILLER_191_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_709 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_191_753 ();
 sky130_fd_sc_hd__decap_8 FILLER_191_758 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_766 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_770 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_778 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_796 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_809 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_815 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_827 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_833 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_192_481 ();
 sky130_fd_sc_hd__decap_8 FILLER_192_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_192_514 ();
 sky130_fd_sc_hd__decap_3 FILLER_192_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_192_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_567 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_607 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_630 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_642 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_668 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_672 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_680 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_686 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_711 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_717 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_732 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_739 ();
 sky130_fd_sc_hd__decap_8 FILLER_192_745 ();
 sky130_fd_sc_hd__decap_3 FILLER_192_753 ();
 sky130_fd_sc_hd__decap_8 FILLER_192_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_765 ();
 sky130_fd_sc_hd__decap_8 FILLER_192_774 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_782 ();
 sky130_fd_sc_hd__decap_8 FILLER_192_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_793 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_818 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_824 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_479 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_482 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_516 ();
 sky130_fd_sc_hd__decap_8 FILLER_193_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_535 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_551 ();
 sky130_fd_sc_hd__decap_3 FILLER_193_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_577 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_581 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_587 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_593 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_615 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_623 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_647 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_659 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_663 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_670 ();
 sky130_fd_sc_hd__decap_3 FILLER_193_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_683 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_689 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_707 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_719 ();
 sky130_fd_sc_hd__decap_3 FILLER_193_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_733 ();
 sky130_fd_sc_hd__decap_8 FILLER_193_742 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_750 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_763 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_769 ();
 sky130_fd_sc_hd__decap_3 FILLER_193_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_789 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_795 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_801 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_811 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_817 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_821 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_824 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_491 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_500 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_506 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_512 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_520 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_551 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_557 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_563 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_575 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_593 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_605 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_194_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_194_637 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_642 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_649 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_662 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_669 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_676 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_688 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_725 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_732 ();
 sky130_fd_sc_hd__decap_8 FILLER_194_738 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_746 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_761 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_765 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_811 ();
 sky130_fd_sc_hd__decap_8 FILLER_194_813 ();
 sky130_fd_sc_hd__decap_3 FILLER_194_821 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_826 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_195_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_471 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_491 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_529 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_535 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_541 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_547 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_195_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_573 ();
 sky130_fd_sc_hd__decap_8 FILLER_195_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_591 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_594 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_606 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_627 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_648 ();
 sky130_fd_sc_hd__decap_8 FILLER_195_660 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_677 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_683 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_705 ();
 sky130_fd_sc_hd__decap_8 FILLER_195_711 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_724 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_738 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_744 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_750 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_756 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_762 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_768 ();
 sky130_fd_sc_hd__decap_8 FILLER_195_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_797 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_809 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_196_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_464 ();
 sky130_fd_sc_hd__decap_3 FILLER_196_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_495 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_514 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_523 ();
 sky130_fd_sc_hd__decap_3 FILLER_196_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_541 ();
 sky130_fd_sc_hd__decap_8 FILLER_196_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_555 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_571 ();
 sky130_fd_sc_hd__decap_8 FILLER_196_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_196_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_196_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_671 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_691 ();
 sky130_fd_sc_hd__decap_3 FILLER_196_697 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_707 ();
 sky130_fd_sc_hd__decap_8 FILLER_196_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_745 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_196_761 ();
 sky130_fd_sc_hd__decap_3 FILLER_196_769 ();
 sky130_fd_sc_hd__decap_8 FILLER_196_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_787 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_790 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_796 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_830 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_197_461 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_466 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_492 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_498 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_547 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_579 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_604 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_633 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_639 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_197_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_697 ();
 sky130_fd_sc_hd__decap_8 FILLER_197_709 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_717 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_197_733 ();
 sky130_fd_sc_hd__decap_3 FILLER_197_741 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_746 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_758 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_764 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_783 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_791 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_801 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_807 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_815 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_822 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_198_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_494 ();
 sky130_fd_sc_hd__decap_8 FILLER_198_506 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_514 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_518 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_522 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_549 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_567 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_573 ();
 sky130_fd_sc_hd__decap_8 FILLER_198_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_593 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_599 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_611 ();
 sky130_fd_sc_hd__decap_3 FILLER_198_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_663 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_735 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_198_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_768 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_774 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_782 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_795 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_808 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_813 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_817 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_823 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_826 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_832 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_836 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_476 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_482 ();
 sky130_fd_sc_hd__decap_8 FILLER_199_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_502 ();
 sky130_fd_sc_hd__decap_8 FILLER_199_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_513 ();
 sky130_fd_sc_hd__decap_8 FILLER_199_516 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_524 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_527 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_547 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_570 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_576 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_585 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_591 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_641 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_644 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_648 ();
 sky130_fd_sc_hd__decap_3 FILLER_199_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_677 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_689 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_199_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_741 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_745 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_748 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_759 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_765 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_771 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_199_789 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_797 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_801 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_821 ();
 sky130_fd_sc_hd__decap_8 FILLER_199_827 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_445 ();
 sky130_fd_sc_hd__decap_8 FILLER_200_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_484 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_490 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_502 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_506 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_514 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_537 ();
 sky130_fd_sc_hd__decap_8 FILLER_200_543 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_551 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_557 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_563 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_596 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_610 ();
 sky130_fd_sc_hd__decap_8 FILLER_200_616 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_628 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_642 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_668 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_674 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_686 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_698 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_701 ();
 sky130_fd_sc_hd__decap_3 FILLER_200_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_718 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_730 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_742 ();
 sky130_fd_sc_hd__decap_3 FILLER_200_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_766 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_772 ();
 sky130_fd_sc_hd__decap_8 FILLER_200_778 ();
 sky130_fd_sc_hd__decap_3 FILLER_200_786 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_791 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_797 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_817 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_447 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_472 ();
 sky130_fd_sc_hd__decap_8 FILLER_201_478 ();
 sky130_fd_sc_hd__decap_8 FILLER_201_488 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_498 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_521 ();
 sky130_fd_sc_hd__decap_8 FILLER_201_538 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_565 ();
 sky130_fd_sc_hd__decap_8 FILLER_201_571 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_579 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_595 ();
 sky130_fd_sc_hd__decap_8 FILLER_201_608 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_638 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_644 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_648 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_652 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_678 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_684 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_696 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_702 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_712 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_718 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_724 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_741 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_755 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_761 ();
 sky130_fd_sc_hd__decap_8 FILLER_201_767 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_775 ();
 sky130_fd_sc_hd__decap_3 FILLER_201_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_789 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_802 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_808 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_812 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_815 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_828 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_457 ();
 sky130_fd_sc_hd__decap_3 FILLER_202_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_487 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_491 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_497 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_503 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_523 ();
 sky130_fd_sc_hd__decap_3 FILLER_202_529 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_540 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_560 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_566 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_609 ();
 sky130_fd_sc_hd__decap_8 FILLER_202_619 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_649 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_653 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_656 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_669 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_675 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_685 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_691 ();
 sky130_fd_sc_hd__decap_3 FILLER_202_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_706 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_719 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_731 ();
 sky130_fd_sc_hd__decap_3 FILLER_202_743 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_761 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_767 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_773 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_790 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_796 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_806 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_817 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_821 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_826 ();
 sky130_fd_sc_hd__decap_3 FILLER_202_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_203_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_203_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_203_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_203_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_203_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_203_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_203_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_203_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_461 ();
 sky130_fd_sc_hd__decap_6 FILLER_203_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_473 ();
 sky130_fd_sc_hd__decap_6 FILLER_203_482 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_515 ();
 sky130_fd_sc_hd__decap_6 FILLER_203_521 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_527 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_550 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_203_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_574 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_580 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_586 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_598 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_602 ();
 sky130_fd_sc_hd__decap_6 FILLER_203_610 ();
 sky130_fd_sc_hd__decap_6 FILLER_203_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_628 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_648 ();
 sky130_fd_sc_hd__decap_6 FILLER_203_654 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_660 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_663 ();
 sky130_fd_sc_hd__decap_3 FILLER_203_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_684 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_695 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_702 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_708 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_717 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_741 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_753 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_759 ();
 sky130_fd_sc_hd__decap_8 FILLER_203_765 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_773 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_789 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_795 ();
 sky130_fd_sc_hd__decap_8 FILLER_203_801 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_809 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_812 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_818 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_204_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_204_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_204_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_204_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_204_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_204_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_204_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_481 ();
 sky130_fd_sc_hd__decap_6 FILLER_204_498 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_504 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_512 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_519 ();
 sky130_fd_sc_hd__decap_6 FILLER_204_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_551 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_557 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_563 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_613 ();
 sky130_fd_sc_hd__decap_3 FILLER_204_625 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_204_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_667 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_711 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_723 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_735 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_741 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_747 ();
 sky130_fd_sc_hd__decap_3 FILLER_204_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_204_761 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_767 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_770 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_794 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_800 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_820 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_827 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_467 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_495 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_205_518 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_538 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_544 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_548 ();
 sky130_fd_sc_hd__decap_3 FILLER_205_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_568 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_574 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_580 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_592 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_604 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_678 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_686 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_692 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_695 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_702 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_708 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_714 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_720 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_724 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_738 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_744 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_750 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_756 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_760 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_763 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_769 ();
 sky130_fd_sc_hd__decap_3 FILLER_205_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_789 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_795 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_799 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_809 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_812 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_818 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_824 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_445 ();
 sky130_fd_sc_hd__decap_3 FILLER_206_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_510 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_516 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_520 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_206_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_545 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_562 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_568 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_577 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_593 ();
 sky130_fd_sc_hd__decap_8 FILLER_206_599 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_611 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_623 ();
 sky130_fd_sc_hd__decap_8 FILLER_206_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_701 ();
 sky130_fd_sc_hd__decap_3 FILLER_206_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_732 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_741 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_747 ();
 sky130_fd_sc_hd__decap_3 FILLER_206_753 ();
 sky130_fd_sc_hd__decap_3 FILLER_206_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_762 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_774 ();
 sky130_fd_sc_hd__decap_8 FILLER_206_786 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_810 ();
 sky130_fd_sc_hd__decap_3 FILLER_206_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_818 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_824 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_469 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_527 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_539 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_542 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_571 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_577 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_207_625 ();
 sky130_fd_sc_hd__decap_3 FILLER_207_633 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_638 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_650 ();
 sky130_fd_sc_hd__decap_8 FILLER_207_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_670 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_207_733 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_741 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_749 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_756 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_762 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_770 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_776 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_794 ();
 sky130_fd_sc_hd__decap_8 FILLER_207_800 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_808 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_811 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_818 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_824 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_489 ();
 sky130_fd_sc_hd__decap_8 FILLER_208_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_512 ();
 sky130_fd_sc_hd__decap_8 FILLER_208_518 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_526 ();
 sky130_fd_sc_hd__decap_3 FILLER_208_529 ();
 sky130_fd_sc_hd__decap_8 FILLER_208_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_544 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_552 ();
 sky130_fd_sc_hd__decap_3 FILLER_208_564 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_614 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_634 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_640 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_665 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_677 ();
 sky130_fd_sc_hd__decap_8 FILLER_208_689 ();
 sky130_fd_sc_hd__decap_3 FILLER_208_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_713 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_725 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_731 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_734 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_761 ();
 sky130_fd_sc_hd__decap_3 FILLER_208_773 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_778 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_784 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_790 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_796 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_804 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_831 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_835 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_209_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_522 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_526 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_529 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_545 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_559 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_570 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_584 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_590 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_635 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_641 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_648 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_683 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_689 ();
 sky130_fd_sc_hd__decap_8 FILLER_209_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_709 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_712 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_718 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_724 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_733 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_737 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_740 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_744 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_750 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_762 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_209_789 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_797 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_800 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_807 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_827 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_834 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_493 ();
 sky130_fd_sc_hd__decap_8 FILLER_210_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_507 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_522 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_528 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_542 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_550 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_556 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_566 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_572 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_576 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_579 ();
 sky130_fd_sc_hd__decap_3 FILLER_210_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_605 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_609 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_626 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_663 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_676 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_689 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_699 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_720 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_734 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_740 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_746 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_752 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_761 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_772 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_778 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_784 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_788 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_791 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_797 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_803 ();
 sky130_fd_sc_hd__decap_3 FILLER_210_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_813 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_831 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_211_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_211_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_211_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_211_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_211_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_211_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_211_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_211_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_472 ();
 sky130_fd_sc_hd__decap_8 FILLER_211_478 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_486 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_495 ();
 sky130_fd_sc_hd__decap_3 FILLER_211_501 ();
 sky130_fd_sc_hd__decap_6 FILLER_211_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_527 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_538 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_542 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_211_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_575 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_583 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_211_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_629 ();
 sky130_fd_sc_hd__decap_8 FILLER_211_641 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_658 ();
 sky130_fd_sc_hd__decap_6 FILLER_211_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_697 ();
 sky130_fd_sc_hd__decap_8 FILLER_211_710 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_718 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_724 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_738 ();
 sky130_fd_sc_hd__decap_8 FILLER_211_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_774 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_780 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_789 ();
 sky130_fd_sc_hd__decap_8 FILLER_211_795 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_803 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_807 ();
 sky130_fd_sc_hd__decap_6 FILLER_211_827 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_833 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_212_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_212_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_212_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_212_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_212_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_212_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_212_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_445 ();
 sky130_fd_sc_hd__decap_3 FILLER_212_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_212_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_212_497 ();
 sky130_fd_sc_hd__decap_6 FILLER_212_511 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_212_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_212_530 ();
 sky130_fd_sc_hd__decap_4 FILLER_212_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_212_543 ();
 sky130_fd_sc_hd__decap_6 FILLER_212_556 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_562 ();
 sky130_fd_sc_hd__decap_4 FILLER_212_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_587 ();
 sky130_fd_sc_hd__decap_8 FILLER_212_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_607 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_619 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_212_660 ();
 sky130_fd_sc_hd__decap_8 FILLER_212_666 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_674 ();
 sky130_fd_sc_hd__decap_4 FILLER_212_686 ();
 sky130_fd_sc_hd__decap_6 FILLER_212_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_212_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_212_706 ();
 sky130_fd_sc_hd__decap_4 FILLER_212_728 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_732 ();
 sky130_fd_sc_hd__decap_6 FILLER_212_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_212_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_212_761 ();
 sky130_fd_sc_hd__decap_8 FILLER_212_773 ();
 sky130_fd_sc_hd__decap_4 FILLER_212_789 ();
 sky130_fd_sc_hd__decap_6 FILLER_212_795 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_801 ();
 sky130_fd_sc_hd__decap_4 FILLER_212_804 ();
 sky130_fd_sc_hd__fill_2 FILLER_212_810 ();
 sky130_fd_sc_hd__decap_4 FILLER_212_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_212_820 ();
 sky130_fd_sc_hd__fill_2 FILLER_212_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_213_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_213_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_213_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_213_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_213_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_213_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_213_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_213_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_213_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_469 ();
 sky130_fd_sc_hd__decap_4 FILLER_213_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_213_479 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_213_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_213_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_213_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_213_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_213_514 ();
 sky130_fd_sc_hd__decap_4 FILLER_213_520 ();
 sky130_fd_sc_hd__decap_4 FILLER_213_526 ();
 sky130_fd_sc_hd__decap_6 FILLER_213_532 ();
 sky130_fd_sc_hd__decap_6 FILLER_213_540 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_546 ();
 sky130_fd_sc_hd__decap_6 FILLER_213_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_213_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_213_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_213_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_579 ();
 sky130_fd_sc_hd__decap_4 FILLER_213_584 ();
 sky130_fd_sc_hd__decap_8 FILLER_213_590 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_598 ();
 sky130_fd_sc_hd__decap_8 FILLER_213_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_213_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_213_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_213_684 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_690 ();
 sky130_fd_sc_hd__decap_4 FILLER_213_694 ();
 sky130_fd_sc_hd__decap_4 FILLER_213_714 ();
 sky130_fd_sc_hd__decap_6 FILLER_213_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_213_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_213_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_213_742 ();
 sky130_fd_sc_hd__decap_4 FILLER_213_749 ();
 sky130_fd_sc_hd__decap_8 FILLER_213_755 ();
 sky130_fd_sc_hd__decap_8 FILLER_213_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_213_778 ();
 sky130_fd_sc_hd__fill_2 FILLER_213_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_213_792 ();
 sky130_fd_sc_hd__decap_4 FILLER_213_810 ();
 sky130_fd_sc_hd__decap_4 FILLER_213_816 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_820 ();
 sky130_fd_sc_hd__decap_4 FILLER_213_823 ();
 sky130_fd_sc_hd__decap_4 FILLER_213_836 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_214_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_214_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_214_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_214_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_214_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_214_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_214_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_214_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_214_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_481 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_493 ();
 sky130_fd_sc_hd__decap_8 FILLER_214_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_214_516 ();
 sky130_fd_sc_hd__fill_2 FILLER_214_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_214_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_214_537 ();
 sky130_fd_sc_hd__decap_8 FILLER_214_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_553 ();
 sky130_fd_sc_hd__decap_4 FILLER_214_564 ();
 sky130_fd_sc_hd__decap_6 FILLER_214_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_214_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_214_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_214_593 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_214_610 ();
 sky130_fd_sc_hd__decap_4 FILLER_214_616 ();
 sky130_fd_sc_hd__decap_4 FILLER_214_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_214_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_669 ();
 sky130_fd_sc_hd__decap_3 FILLER_214_681 ();
 sky130_fd_sc_hd__decap_8 FILLER_214_686 ();
 sky130_fd_sc_hd__fill_2 FILLER_214_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_214_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_214_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_214_705 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_709 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_712 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_724 ();
 sky130_fd_sc_hd__fill_2 FILLER_214_736 ();
 sky130_fd_sc_hd__decap_4 FILLER_214_740 ();
 sky130_fd_sc_hd__decap_8 FILLER_214_746 ();
 sky130_fd_sc_hd__fill_2 FILLER_214_754 ();
 sky130_fd_sc_hd__decap_6 FILLER_214_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_763 ();
 sky130_fd_sc_hd__decap_4 FILLER_214_766 ();
 sky130_fd_sc_hd__decap_4 FILLER_214_778 ();
 sky130_fd_sc_hd__decap_4 FILLER_214_798 ();
 sky130_fd_sc_hd__decap_4 FILLER_214_804 ();
 sky130_fd_sc_hd__fill_2 FILLER_214_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_214_813 ();
 sky130_fd_sc_hd__decap_6 FILLER_214_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_214_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_214_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_214_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_215_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_215_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_215_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_215_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_215_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_215_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_215_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_215_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_215_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_215_469 ();
 sky130_fd_sc_hd__decap_4 FILLER_215_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_479 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_215_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_215_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_215_519 ();
 sky130_fd_sc_hd__decap_4 FILLER_215_532 ();
 sky130_fd_sc_hd__decap_4 FILLER_215_542 ();
 sky130_fd_sc_hd__decap_4 FILLER_215_550 ();
 sky130_fd_sc_hd__decap_4 FILLER_215_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_215_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_215_569 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_575 ();
 sky130_fd_sc_hd__decap_4 FILLER_215_583 ();
 sky130_fd_sc_hd__decap_6 FILLER_215_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_595 ();
 sky130_fd_sc_hd__decap_4 FILLER_215_604 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_608 ();
 sky130_fd_sc_hd__decap_4 FILLER_215_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_615 ();
 sky130_fd_sc_hd__decap_6 FILLER_215_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_215_631 ();
 sky130_fd_sc_hd__decap_4 FILLER_215_637 ();
 sky130_fd_sc_hd__decap_4 FILLER_215_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_649 ();
 sky130_fd_sc_hd__decap_8 FILLER_215_661 ();
 sky130_fd_sc_hd__decap_3 FILLER_215_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_215_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_215_684 ();
 sky130_fd_sc_hd__decap_4 FILLER_215_690 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_696 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_708 ();
 sky130_fd_sc_hd__decap_8 FILLER_215_720 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_741 ();
 sky130_fd_sc_hd__decap_6 FILLER_215_753 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_759 ();
 sky130_fd_sc_hd__decap_4 FILLER_215_762 ();
 sky130_fd_sc_hd__fill_2 FILLER_215_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_215_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_215_789 ();
 sky130_fd_sc_hd__decap_4 FILLER_215_799 ();
 sky130_fd_sc_hd__decap_4 FILLER_215_812 ();
 sky130_fd_sc_hd__decap_8 FILLER_215_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_833 ();
 sky130_fd_sc_hd__fill_2 FILLER_215_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_216_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_216_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_216_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_216_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_216_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_216_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_216_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_445 ();
 sky130_fd_sc_hd__decap_6 FILLER_216_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_216_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_216_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_216_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_216_495 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_216_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_216_521 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_527 ();
 sky130_fd_sc_hd__fill_2 FILLER_216_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_216_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_216_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_216_543 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_216_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_216_566 ();
 sky130_fd_sc_hd__decap_6 FILLER_216_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_216_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_216_593 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_216_609 ();
 sky130_fd_sc_hd__decap_6 FILLER_216_615 ();
 sky130_fd_sc_hd__decap_6 FILLER_216_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_216_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_216_653 ();
 sky130_fd_sc_hd__decap_4 FILLER_216_659 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_663 ();
 sky130_fd_sc_hd__decap_4 FILLER_216_680 ();
 sky130_fd_sc_hd__decap_4 FILLER_216_687 ();
 sky130_fd_sc_hd__decap_6 FILLER_216_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_216_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_705 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_216_733 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_216_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_755 ();
 sky130_fd_sc_hd__decap_8 FILLER_216_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_765 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_768 ();
 sky130_fd_sc_hd__fill_2 FILLER_216_780 ();
 sky130_fd_sc_hd__decap_4 FILLER_216_784 ();
 sky130_fd_sc_hd__decap_4 FILLER_216_790 ();
 sky130_fd_sc_hd__fill_2 FILLER_216_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_216_813 ();
 sky130_fd_sc_hd__decap_6 FILLER_216_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_216_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_829 ();
 sky130_fd_sc_hd__decap_4 FILLER_216_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_216_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_217_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_217_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_217_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_217_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_217_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_217_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_217_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_217_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_217_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_453 ();
 sky130_fd_sc_hd__decap_6 FILLER_217_470 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_492 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_217_517 ();
 sky130_fd_sc_hd__decap_8 FILLER_217_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_217_536 ();
 sky130_fd_sc_hd__decap_4 FILLER_217_542 ();
 sky130_fd_sc_hd__decap_4 FILLER_217_548 ();
 sky130_fd_sc_hd__decap_6 FILLER_217_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_217_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_217_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_217_575 ();
 sky130_fd_sc_hd__decap_4 FILLER_217_588 ();
 sky130_fd_sc_hd__decap_6 FILLER_217_594 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_217_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_217_614 ();
 sky130_fd_sc_hd__decap_4 FILLER_217_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_217_624 ();
 sky130_fd_sc_hd__decap_4 FILLER_217_630 ();
 sky130_fd_sc_hd__decap_4 FILLER_217_638 ();
 sky130_fd_sc_hd__decap_4 FILLER_217_659 ();
 sky130_fd_sc_hd__decap_6 FILLER_217_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_217_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_217_682 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_686 ();
 sky130_fd_sc_hd__decap_4 FILLER_217_692 ();
 sky130_fd_sc_hd__decap_4 FILLER_217_698 ();
 sky130_fd_sc_hd__decap_4 FILLER_217_704 ();
 sky130_fd_sc_hd__decap_4 FILLER_217_710 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_716 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_217_741 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_745 ();
 sky130_fd_sc_hd__decap_4 FILLER_217_762 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_768 ();
 sky130_fd_sc_hd__decap_4 FILLER_217_780 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_785 ();
 sky130_fd_sc_hd__decap_3 FILLER_217_797 ();
 sky130_fd_sc_hd__decap_4 FILLER_217_803 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_807 ();
 sky130_fd_sc_hd__decap_4 FILLER_217_810 ();
 sky130_fd_sc_hd__decap_4 FILLER_217_816 ();
 sky130_fd_sc_hd__decap_6 FILLER_217_822 ();
 sky130_fd_sc_hd__decap_4 FILLER_217_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_217_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_218_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_218_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_218_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_218_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_218_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_218_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_218_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_445 ();
 sky130_fd_sc_hd__decap_8 FILLER_218_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_218_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_218_474 ();
 sky130_fd_sc_hd__decap_3 FILLER_218_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_218_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_218_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_495 ();
 sky130_fd_sc_hd__decap_4 FILLER_218_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_218_521 ();
 sky130_fd_sc_hd__decap_4 FILLER_218_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_531 ();
 sky130_fd_sc_hd__decap_6 FILLER_218_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_539 ();
 sky130_fd_sc_hd__decap_4 FILLER_218_548 ();
 sky130_fd_sc_hd__decap_4 FILLER_218_557 ();
 sky130_fd_sc_hd__decap_4 FILLER_218_563 ();
 sky130_fd_sc_hd__decap_8 FILLER_218_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_218_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_218_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_218_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_218_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_218_605 ();
 sky130_fd_sc_hd__decap_4 FILLER_218_611 ();
 sky130_fd_sc_hd__decap_6 FILLER_218_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_623 ();
 sky130_fd_sc_hd__decap_6 FILLER_218_626 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_632 ();
 sky130_fd_sc_hd__decap_4 FILLER_218_635 ();
 sky130_fd_sc_hd__fill_2 FILLER_218_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_218_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_218_655 ();
 sky130_fd_sc_hd__decap_4 FILLER_218_661 ();
 sky130_fd_sc_hd__decap_4 FILLER_218_674 ();
 sky130_fd_sc_hd__decap_8 FILLER_218_680 ();
 sky130_fd_sc_hd__decap_4 FILLER_218_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_218_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_218_706 ();
 sky130_fd_sc_hd__decap_4 FILLER_218_712 ();
 sky130_fd_sc_hd__decap_4 FILLER_218_718 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_724 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_736 ();
 sky130_fd_sc_hd__decap_8 FILLER_218_748 ();
 sky130_fd_sc_hd__fill_2 FILLER_218_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_218_767 ();
 sky130_fd_sc_hd__decap_4 FILLER_218_773 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_779 ();
 sky130_fd_sc_hd__decap_8 FILLER_218_791 ();
 sky130_fd_sc_hd__decap_3 FILLER_218_799 ();
 sky130_fd_sc_hd__decap_4 FILLER_218_804 ();
 sky130_fd_sc_hd__fill_2 FILLER_218_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_218_813 ();
 sky130_fd_sc_hd__decap_6 FILLER_218_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_218_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_218_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_219_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_219_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_219_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_219_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_219_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_219_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_219_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_219_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_219_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_467 ();
 sky130_fd_sc_hd__decap_4 FILLER_219_470 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_476 ();
 sky130_fd_sc_hd__decap_8 FILLER_219_488 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_496 ();
 sky130_fd_sc_hd__decap_4 FILLER_219_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_219_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_219_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_219_521 ();
 sky130_fd_sc_hd__decap_6 FILLER_219_527 ();
 sky130_fd_sc_hd__decap_4 FILLER_219_535 ();
 sky130_fd_sc_hd__decap_6 FILLER_219_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_219_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_219_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_219_583 ();
 sky130_fd_sc_hd__decap_6 FILLER_219_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_219_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_219_621 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_219_630 ();
 sky130_fd_sc_hd__decap_4 FILLER_219_642 ();
 sky130_fd_sc_hd__decap_8 FILLER_219_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_219_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_219_677 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_681 ();
 sky130_fd_sc_hd__decap_4 FILLER_219_699 ();
 sky130_fd_sc_hd__decap_4 FILLER_219_711 ();
 sky130_fd_sc_hd__decap_4 FILLER_219_717 ();
 sky130_fd_sc_hd__decap_4 FILLER_219_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_219_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_219_733 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_767 ();
 sky130_fd_sc_hd__decap_4 FILLER_219_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_785 ();
 sky130_fd_sc_hd__decap_3 FILLER_219_797 ();
 sky130_fd_sc_hd__decap_4 FILLER_219_802 ();
 sky130_fd_sc_hd__decap_4 FILLER_219_812 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_816 ();
 sky130_fd_sc_hd__decap_4 FILLER_219_820 ();
 sky130_fd_sc_hd__decap_6 FILLER_219_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_839 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_220_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_220_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_220_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_220_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_220_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_220_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_220_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_220_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_220_497 ();
 sky130_fd_sc_hd__decap_4 FILLER_220_512 ();
 sky130_fd_sc_hd__decap_4 FILLER_220_518 ();
 sky130_fd_sc_hd__decap_4 FILLER_220_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_220_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_220_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_220_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_220_562 ();
 sky130_fd_sc_hd__decap_4 FILLER_220_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_220_578 ();
 sky130_fd_sc_hd__decap_4 FILLER_220_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_220_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_220_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_220_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_220_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_220_633 ();
 sky130_fd_sc_hd__decap_4 FILLER_220_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_220_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_220_650 ();
 sky130_fd_sc_hd__decap_4 FILLER_220_656 ();
 sky130_fd_sc_hd__decap_4 FILLER_220_662 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_666 ();
 sky130_fd_sc_hd__decap_4 FILLER_220_674 ();
 sky130_fd_sc_hd__decap_8 FILLER_220_680 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_688 ();
 sky130_fd_sc_hd__decap_4 FILLER_220_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_220_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_220_705 ();
 sky130_fd_sc_hd__decap_8 FILLER_220_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_725 ();
 sky130_fd_sc_hd__decap_4 FILLER_220_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_220_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_220_748 ();
 sky130_fd_sc_hd__fill_2 FILLER_220_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_220_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_762 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_774 ();
 sky130_fd_sc_hd__decap_8 FILLER_220_786 ();
 sky130_fd_sc_hd__decap_4 FILLER_220_796 ();
 sky130_fd_sc_hd__decap_4 FILLER_220_802 ();
 sky130_fd_sc_hd__decap_4 FILLER_220_808 ();
 sky130_fd_sc_hd__decap_4 FILLER_220_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_220_820 ();
 sky130_fd_sc_hd__fill_2 FILLER_220_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_221_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_221_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_221_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_221_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_221_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_221_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_221_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_221_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_221_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_221_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_221_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_221_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_221_521 ();
 sky130_fd_sc_hd__decap_4 FILLER_221_534 ();
 sky130_fd_sc_hd__decap_4 FILLER_221_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_221_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_221_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_221_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_221_578 ();
 sky130_fd_sc_hd__decap_4 FILLER_221_584 ();
 sky130_fd_sc_hd__decap_4 FILLER_221_590 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_594 ();
 sky130_fd_sc_hd__decap_4 FILLER_221_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_221_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_221_641 ();
 sky130_fd_sc_hd__decap_4 FILLER_221_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_221_651 ();
 sky130_fd_sc_hd__decap_4 FILLER_221_657 ();
 sky130_fd_sc_hd__decap_8 FILLER_221_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_671 ();
 sky130_fd_sc_hd__decap_6 FILLER_221_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_679 ();
 sky130_fd_sc_hd__decap_6 FILLER_221_682 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_688 ();
 sky130_fd_sc_hd__decap_4 FILLER_221_693 ();
 sky130_fd_sc_hd__decap_4 FILLER_221_700 ();
 sky130_fd_sc_hd__decap_4 FILLER_221_706 ();
 sky130_fd_sc_hd__fill_2 FILLER_221_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_221_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_221_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_221_752 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_758 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_770 ();
 sky130_fd_sc_hd__fill_2 FILLER_221_782 ();
 sky130_fd_sc_hd__decap_3 FILLER_221_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_221_790 ();
 sky130_fd_sc_hd__decap_4 FILLER_221_802 ();
 sky130_fd_sc_hd__decap_6 FILLER_221_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_221_822 ();
 sky130_fd_sc_hd__decap_4 FILLER_221_829 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_833 ();
 sky130_fd_sc_hd__fill_2 FILLER_221_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_222_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_222_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_222_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_222_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_222_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_222_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_222_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_445 ();
 sky130_fd_sc_hd__decap_6 FILLER_222_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_222_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_222_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_222_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_222_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_222_495 ();
 sky130_fd_sc_hd__decap_8 FILLER_222_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_222_509 ();
 sky130_fd_sc_hd__decap_6 FILLER_222_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_222_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_222_530 ();
 sky130_fd_sc_hd__decap_3 FILLER_222_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_222_538 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_546 ();
 sky130_fd_sc_hd__decap_4 FILLER_222_554 ();
 sky130_fd_sc_hd__decap_4 FILLER_222_563 ();
 sky130_fd_sc_hd__decap_4 FILLER_222_570 ();
 sky130_fd_sc_hd__decap_4 FILLER_222_576 ();
 sky130_fd_sc_hd__decap_6 FILLER_222_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_222_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_222_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_222_606 ();
 sky130_fd_sc_hd__decap_4 FILLER_222_612 ();
 sky130_fd_sc_hd__decap_4 FILLER_222_624 ();
 sky130_fd_sc_hd__decap_4 FILLER_222_630 ();
 sky130_fd_sc_hd__decap_8 FILLER_222_636 ();
 sky130_fd_sc_hd__decap_4 FILLER_222_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_649 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_652 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_664 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_676 ();
 sky130_fd_sc_hd__decap_4 FILLER_222_688 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_692 ();
 sky130_fd_sc_hd__decap_4 FILLER_222_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_222_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_222_705 ();
 sky130_fd_sc_hd__decap_8 FILLER_222_712 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_720 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_724 ();
 sky130_fd_sc_hd__decap_3 FILLER_222_736 ();
 sky130_fd_sc_hd__decap_4 FILLER_222_741 ();
 sky130_fd_sc_hd__decap_4 FILLER_222_747 ();
 sky130_fd_sc_hd__decap_3 FILLER_222_753 ();
 sky130_fd_sc_hd__decap_8 FILLER_222_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_765 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_768 ();
 sky130_fd_sc_hd__fill_2 FILLER_222_780 ();
 sky130_fd_sc_hd__decap_4 FILLER_222_784 ();
 sky130_fd_sc_hd__decap_4 FILLER_222_790 ();
 sky130_fd_sc_hd__fill_2 FILLER_222_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_222_813 ();
 sky130_fd_sc_hd__decap_6 FILLER_222_817 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_823 ();
 sky130_fd_sc_hd__fill_2 FILLER_222_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_223_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_223_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_223_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_223_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_223_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_223_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_223_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_223_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_223_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_223_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_479 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_223_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_523 ();
 sky130_fd_sc_hd__decap_8 FILLER_223_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_223_534 ();
 sky130_fd_sc_hd__decap_4 FILLER_223_538 ();
 sky130_fd_sc_hd__decap_4 FILLER_223_549 ();
 sky130_fd_sc_hd__decap_4 FILLER_223_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_223_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_223_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_223_575 ();
 sky130_fd_sc_hd__decap_4 FILLER_223_581 ();
 sky130_fd_sc_hd__decap_4 FILLER_223_587 ();
 sky130_fd_sc_hd__decap_4 FILLER_223_593 ();
 sky130_fd_sc_hd__decap_8 FILLER_223_599 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_607 ();
 sky130_fd_sc_hd__decap_6 FILLER_223_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_223_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_223_635 ();
 sky130_fd_sc_hd__decap_4 FILLER_223_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_647 ();
 sky130_fd_sc_hd__decap_8 FILLER_223_659 ();
 sky130_fd_sc_hd__decap_3 FILLER_223_669 ();
 sky130_fd_sc_hd__decap_8 FILLER_223_673 ();
 sky130_fd_sc_hd__decap_3 FILLER_223_681 ();
 sky130_fd_sc_hd__decap_4 FILLER_223_686 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_707 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_710 ();
 sky130_fd_sc_hd__decap_6 FILLER_223_722 ();
 sky130_fd_sc_hd__decap_8 FILLER_223_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_737 ();
 sky130_fd_sc_hd__decap_8 FILLER_223_746 ();
 sky130_fd_sc_hd__decap_4 FILLER_223_761 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_765 ();
 sky130_fd_sc_hd__fill_2 FILLER_223_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_223_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_223_795 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_803 ();
 sky130_fd_sc_hd__decap_4 FILLER_223_812 ();
 sky130_fd_sc_hd__decap_4 FILLER_223_818 ();
 sky130_fd_sc_hd__decap_4 FILLER_223_824 ();
 sky130_fd_sc_hd__decap_4 FILLER_223_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_223_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_224_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_224_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_224_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_224_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_224_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_224_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_224_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_445 ();
 sky130_fd_sc_hd__decap_8 FILLER_224_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_224_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_224_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_224_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_481 ();
 sky130_fd_sc_hd__decap_8 FILLER_224_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_224_521 ();
 sky130_fd_sc_hd__decap_4 FILLER_224_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_531 ();
 sky130_fd_sc_hd__decap_6 FILLER_224_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_539 ();
 sky130_fd_sc_hd__decap_4 FILLER_224_542 ();
 sky130_fd_sc_hd__decap_4 FILLER_224_548 ();
 sky130_fd_sc_hd__decap_4 FILLER_224_554 ();
 sky130_fd_sc_hd__decap_8 FILLER_224_560 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_568 ();
 sky130_fd_sc_hd__decap_4 FILLER_224_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_224_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_224_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_224_593 ();
 sky130_fd_sc_hd__decap_8 FILLER_224_599 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_607 ();
 sky130_fd_sc_hd__decap_6 FILLER_224_610 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_616 ();
 sky130_fd_sc_hd__decap_4 FILLER_224_620 ();
 sky130_fd_sc_hd__decap_8 FILLER_224_626 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_634 ();
 sky130_fd_sc_hd__decap_6 FILLER_224_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_224_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_224_649 ();
 sky130_fd_sc_hd__decap_8 FILLER_224_655 ();
 sky130_fd_sc_hd__decap_4 FILLER_224_665 ();
 sky130_fd_sc_hd__decap_4 FILLER_224_678 ();
 sky130_fd_sc_hd__decap_4 FILLER_224_684 ();
 sky130_fd_sc_hd__decap_8 FILLER_224_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_224_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_224_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_711 ();
 sky130_fd_sc_hd__decap_8 FILLER_224_723 ();
 sky130_fd_sc_hd__decap_4 FILLER_224_747 ();
 sky130_fd_sc_hd__decap_3 FILLER_224_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_224_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_224_764 ();
 sky130_fd_sc_hd__decap_4 FILLER_224_784 ();
 sky130_fd_sc_hd__decap_4 FILLER_224_795 ();
 sky130_fd_sc_hd__decap_6 FILLER_224_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_224_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_224_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_224_823 ();
 sky130_fd_sc_hd__decap_4 FILLER_224_830 ();
 sky130_fd_sc_hd__decap_4 FILLER_224_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_225_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_225_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_225_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_225_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_225_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_225_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_225_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_225_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_461 ();
 sky130_fd_sc_hd__decap_6 FILLER_225_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_479 ();
 sky130_fd_sc_hd__decap_4 FILLER_225_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_225_494 ();
 sky130_fd_sc_hd__decap_4 FILLER_225_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_225_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_225_509 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_225_518 ();
 sky130_fd_sc_hd__decap_4 FILLER_225_538 ();
 sky130_fd_sc_hd__decap_4 FILLER_225_544 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_548 ();
 sky130_fd_sc_hd__decap_4 FILLER_225_551 ();
 sky130_fd_sc_hd__decap_3 FILLER_225_557 ();
 sky130_fd_sc_hd__decap_6 FILLER_225_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_567 ();
 sky130_fd_sc_hd__decap_4 FILLER_225_575 ();
 sky130_fd_sc_hd__decap_6 FILLER_225_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_225_606 ();
 sky130_fd_sc_hd__decap_4 FILLER_225_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_225_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_225_621 ();
 sky130_fd_sc_hd__decap_8 FILLER_225_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_225_643 ();
 sky130_fd_sc_hd__decap_6 FILLER_225_649 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_655 ();
 sky130_fd_sc_hd__decap_6 FILLER_225_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_225_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_225_678 ();
 sky130_fd_sc_hd__decap_4 FILLER_225_698 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_702 ();
 sky130_fd_sc_hd__decap_4 FILLER_225_709 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_715 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_225_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_225_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_225_742 ();
 sky130_fd_sc_hd__decap_4 FILLER_225_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_753 ();
 sky130_fd_sc_hd__decap_4 FILLER_225_758 ();
 sky130_fd_sc_hd__decap_4 FILLER_225_766 ();
 sky130_fd_sc_hd__decap_8 FILLER_225_773 ();
 sky130_fd_sc_hd__decap_3 FILLER_225_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_225_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_225_804 ();
 sky130_fd_sc_hd__decap_4 FILLER_225_810 ();
 sky130_fd_sc_hd__decap_4 FILLER_225_816 ();
 sky130_fd_sc_hd__decap_6 FILLER_225_822 ();
 sky130_fd_sc_hd__decap_4 FILLER_225_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_225_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_226_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_226_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_226_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_226_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_226_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_226_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_226_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_226_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_226_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_226_495 ();
 sky130_fd_sc_hd__decap_4 FILLER_226_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_226_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_226_521 ();
 sky130_fd_sc_hd__decap_4 FILLER_226_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_226_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_226_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_541 ();
 sky130_fd_sc_hd__decap_8 FILLER_226_544 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_552 ();
 sky130_fd_sc_hd__decap_4 FILLER_226_555 ();
 sky130_fd_sc_hd__decap_4 FILLER_226_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_226_567 ();
 sky130_fd_sc_hd__decap_4 FILLER_226_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_226_579 ();
 sky130_fd_sc_hd__decap_3 FILLER_226_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_226_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_226_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_226_599 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_605 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_226_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_226_635 ();
 sky130_fd_sc_hd__decap_3 FILLER_226_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_226_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_226_666 ();
 sky130_fd_sc_hd__decap_4 FILLER_226_686 ();
 sky130_fd_sc_hd__decap_8 FILLER_226_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_226_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_226_719 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_725 ();
 sky130_fd_sc_hd__decap_4 FILLER_226_737 ();
 sky130_fd_sc_hd__decap_4 FILLER_226_743 ();
 sky130_fd_sc_hd__decap_6 FILLER_226_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_226_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_226_788 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_794 ();
 sky130_fd_sc_hd__decap_6 FILLER_226_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_803 ();
 sky130_fd_sc_hd__decap_6 FILLER_226_806 ();
 sky130_fd_sc_hd__decap_3 FILLER_226_813 ();
 sky130_fd_sc_hd__decap_6 FILLER_226_823 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_829 ();
 sky130_fd_sc_hd__decap_4 FILLER_226_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_226_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_227_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_227_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_227_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_227_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_227_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_227_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_227_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_227_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_227_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_227_480 ();
 sky130_fd_sc_hd__decap_8 FILLER_227_486 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_227_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_227_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_227_516 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_522 ();
 sky130_fd_sc_hd__decap_4 FILLER_227_539 ();
 sky130_fd_sc_hd__decap_4 FILLER_227_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_227_551 ();
 sky130_fd_sc_hd__decap_3 FILLER_227_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_227_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_227_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_227_582 ();
 sky130_fd_sc_hd__decap_4 FILLER_227_594 ();
 sky130_fd_sc_hd__decap_4 FILLER_227_600 ();
 sky130_fd_sc_hd__decap_8 FILLER_227_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_227_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_227_629 ();
 sky130_fd_sc_hd__decap_8 FILLER_227_638 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_646 ();
 sky130_fd_sc_hd__decap_4 FILLER_227_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_227_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_227_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_227_684 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_690 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_702 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_227_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_227_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_797 ();
 sky130_fd_sc_hd__decap_6 FILLER_227_809 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_815 ();
 sky130_fd_sc_hd__decap_4 FILLER_227_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_227_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_228_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_228_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_228_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_228_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_228_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_228_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_228_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_228_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_228_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_481 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_484 ();
 sky130_fd_sc_hd__decap_3 FILLER_228_496 ();
 sky130_fd_sc_hd__decap_6 FILLER_228_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_228_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_228_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_228_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_228_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_228_550 ();
 sky130_fd_sc_hd__decap_6 FILLER_228_556 ();
 sky130_fd_sc_hd__decap_4 FILLER_228_578 ();
 sky130_fd_sc_hd__decap_4 FILLER_228_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_228_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_228_599 ();
 sky130_fd_sc_hd__decap_8 FILLER_228_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_228_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_228_623 ();
 sky130_fd_sc_hd__decap_4 FILLER_228_629 ();
 sky130_fd_sc_hd__decap_8 FILLER_228_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_643 ();
 sky130_fd_sc_hd__decap_6 FILLER_228_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_651 ();
 sky130_fd_sc_hd__decap_8 FILLER_228_655 ();
 sky130_fd_sc_hd__decap_4 FILLER_228_683 ();
 sky130_fd_sc_hd__decap_8 FILLER_228_689 ();
 sky130_fd_sc_hd__decap_3 FILLER_228_697 ();
 sky130_fd_sc_hd__decap_8 FILLER_228_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_228_709 ();
 sky130_fd_sc_hd__decap_4 FILLER_228_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_228_722 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_726 ();
 sky130_fd_sc_hd__decap_8 FILLER_228_729 ();
 sky130_fd_sc_hd__decap_3 FILLER_228_737 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_742 ();
 sky130_fd_sc_hd__fill_2 FILLER_228_754 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_228_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_811 ();
 sky130_fd_sc_hd__decap_4 FILLER_228_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_228_819 ();
 sky130_fd_sc_hd__decap_4 FILLER_228_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_829 ();
 sky130_fd_sc_hd__decap_4 FILLER_228_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_228_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_229_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_229_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_229_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_229_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_229_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_229_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_229_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_229_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_229_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_229_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_229_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_229_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_229_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_229_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_229_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_229_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_485 ();
 sky130_fd_sc_hd__decap_3 FILLER_229_497 ();
 sky130_fd_sc_hd__fill_2 FILLER_229_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_229_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_229_515 ();
 sky130_fd_sc_hd__fill_1 FILLER_229_521 ();
 sky130_fd_sc_hd__decap_8 FILLER_229_532 ();
 sky130_fd_sc_hd__fill_1 FILLER_229_540 ();
 sky130_fd_sc_hd__decap_3 FILLER_229_557 ();
 sky130_fd_sc_hd__decap_4 FILLER_229_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_229_568 ();
 sky130_fd_sc_hd__decap_4 FILLER_229_574 ();
 sky130_fd_sc_hd__fill_1 FILLER_229_578 ();
 sky130_fd_sc_hd__decap_4 FILLER_229_585 ();
 sky130_fd_sc_hd__decap_4 FILLER_229_592 ();
 sky130_fd_sc_hd__decap_4 FILLER_229_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_229_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_229_635 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_641 ();
 sky130_fd_sc_hd__decap_8 FILLER_229_653 ();
 sky130_fd_sc_hd__decap_3 FILLER_229_661 ();
 sky130_fd_sc_hd__decap_6 FILLER_229_666 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_685 ();
 sky130_fd_sc_hd__decap_4 FILLER_229_697 ();
 sky130_fd_sc_hd__fill_1 FILLER_229_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_229_704 ();
 sky130_fd_sc_hd__decap_4 FILLER_229_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_229_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_229_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_229_733 ();
 sky130_fd_sc_hd__fill_1 FILLER_229_741 ();
 sky130_fd_sc_hd__decap_8 FILLER_229_746 ();
 sky130_fd_sc_hd__fill_1 FILLER_229_754 ();
 sky130_fd_sc_hd__decap_4 FILLER_229_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_229_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_229_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_229_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_229_801 ();
 sky130_fd_sc_hd__decap_4 FILLER_229_804 ();
 sky130_fd_sc_hd__decap_4 FILLER_229_810 ();
 sky130_fd_sc_hd__decap_4 FILLER_229_816 ();
 sky130_fd_sc_hd__decap_4 FILLER_229_822 ();
 sky130_fd_sc_hd__decap_6 FILLER_229_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_229_839 ();
 sky130_fd_sc_hd__fill_1 FILLER_229_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_230_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_230_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_230_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_230_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_230_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_230_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_230_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_230_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_489 ();
 sky130_fd_sc_hd__decap_6 FILLER_230_501 ();
 sky130_fd_sc_hd__decap_6 FILLER_230_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_230_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_230_523 ();
 sky130_fd_sc_hd__decap_3 FILLER_230_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_230_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_230_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_230_563 ();
 sky130_fd_sc_hd__decap_4 FILLER_230_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_230_575 ();
 sky130_fd_sc_hd__decap_6 FILLER_230_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_230_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_230_593 ();
 sky130_fd_sc_hd__decap_8 FILLER_230_599 ();
 sky130_fd_sc_hd__decap_3 FILLER_230_607 ();
 sky130_fd_sc_hd__decap_4 FILLER_230_612 ();
 sky130_fd_sc_hd__decap_4 FILLER_230_619 ();
 sky130_fd_sc_hd__decap_4 FILLER_230_625 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_230_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_699 ();
 sky130_fd_sc_hd__decap_3 FILLER_230_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_230_706 ();
 sky130_fd_sc_hd__decap_4 FILLER_230_726 ();
 sky130_fd_sc_hd__decap_6 FILLER_230_736 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_742 ();
 sky130_fd_sc_hd__decap_6 FILLER_230_745 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_751 ();
 sky130_fd_sc_hd__fill_2 FILLER_230_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_230_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_230_787 ();
 sky130_fd_sc_hd__decap_4 FILLER_230_792 ();
 sky130_fd_sc_hd__decap_6 FILLER_230_798 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_804 ();
 sky130_fd_sc_hd__decap_4 FILLER_230_808 ();
 sky130_fd_sc_hd__decap_4 FILLER_230_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_230_819 ();
 sky130_fd_sc_hd__decap_4 FILLER_230_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_230_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_231_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_231_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_231_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_231_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_231_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_231_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_231_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_231_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_231_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_231_472 ();
 sky130_fd_sc_hd__decap_4 FILLER_231_478 ();
 sky130_fd_sc_hd__decap_6 FILLER_231_484 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_490 ();
 sky130_fd_sc_hd__decap_8 FILLER_231_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_231_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_231_529 ();
 sky130_fd_sc_hd__decap_6 FILLER_231_534 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_540 ();
 sky130_fd_sc_hd__decap_4 FILLER_231_546 ();
 sky130_fd_sc_hd__decap_4 FILLER_231_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_231_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_231_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_231_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_231_571 ();
 sky130_fd_sc_hd__decap_8 FILLER_231_577 ();
 sky130_fd_sc_hd__decap_4 FILLER_231_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_593 ();
 sky130_fd_sc_hd__decap_8 FILLER_231_605 ();
 sky130_fd_sc_hd__decap_3 FILLER_231_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_231_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_649 ();
 sky130_fd_sc_hd__decap_8 FILLER_231_661 ();
 sky130_fd_sc_hd__decap_3 FILLER_231_669 ();
 sky130_fd_sc_hd__decap_4 FILLER_231_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_231_680 ();
 sky130_fd_sc_hd__decap_4 FILLER_231_693 ();
 sky130_fd_sc_hd__decap_4 FILLER_231_699 ();
 sky130_fd_sc_hd__decap_6 FILLER_231_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_231_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_231_719 ();
 sky130_fd_sc_hd__fill_2 FILLER_231_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_231_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_231_741 ();
 sky130_fd_sc_hd__decap_4 FILLER_231_749 ();
 sky130_fd_sc_hd__decap_4 FILLER_231_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_231_764 ();
 sky130_fd_sc_hd__fill_2 FILLER_231_772 ();
 sky130_fd_sc_hd__decap_4 FILLER_231_780 ();
 sky130_fd_sc_hd__fill_2 FILLER_231_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_231_794 ();
 sky130_fd_sc_hd__decap_4 FILLER_231_800 ();
 sky130_fd_sc_hd__decap_8 FILLER_231_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_821 ();
 sky130_fd_sc_hd__fill_2 FILLER_231_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_232_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_232_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_232_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_232_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_232_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_232_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_232_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_445 ();
 sky130_fd_sc_hd__decap_3 FILLER_232_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_232_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_232_474 ();
 sky130_fd_sc_hd__decap_6 FILLER_232_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_232_491 ();
 sky130_fd_sc_hd__decap_4 FILLER_232_497 ();
 sky130_fd_sc_hd__decap_4 FILLER_232_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_507 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_510 ();
 sky130_fd_sc_hd__decap_8 FILLER_232_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_232_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_232_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_232_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_232_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_232_549 ();
 sky130_fd_sc_hd__decap_8 FILLER_232_555 ();
 sky130_fd_sc_hd__fill_2 FILLER_232_563 ();
 sky130_fd_sc_hd__decap_4 FILLER_232_567 ();
 sky130_fd_sc_hd__decap_4 FILLER_232_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_232_579 ();
 sky130_fd_sc_hd__decap_3 FILLER_232_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_232_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_593 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_605 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_232_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_232_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_232_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_232_649 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_658 ();
 sky130_fd_sc_hd__decap_4 FILLER_232_670 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_674 ();
 sky130_fd_sc_hd__decap_4 FILLER_232_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_232_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_232_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_232_711 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_717 ();
 sky130_fd_sc_hd__decap_4 FILLER_232_723 ();
 sky130_fd_sc_hd__decap_4 FILLER_232_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_232_738 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_744 ();
 sky130_fd_sc_hd__decap_6 FILLER_232_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_763 ();
 sky130_fd_sc_hd__decap_4 FILLER_232_766 ();
 sky130_fd_sc_hd__decap_4 FILLER_232_772 ();
 sky130_fd_sc_hd__decap_6 FILLER_232_784 ();
 sky130_fd_sc_hd__decap_4 FILLER_232_798 ();
 sky130_fd_sc_hd__fill_2 FILLER_232_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_232_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_232_820 ();
 sky130_fd_sc_hd__decap_4 FILLER_232_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_232_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_233_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_233_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_233_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_233_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_233_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_233_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_233_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_233_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_233_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_233_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_233_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_233_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_233_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_233_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_233_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_233_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_233_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_233_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_233_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_233_495 ();
 sky130_fd_sc_hd__decap_3 FILLER_233_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_233_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_233_509 ();
 sky130_fd_sc_hd__decap_6 FILLER_233_515 ();
 sky130_fd_sc_hd__fill_1 FILLER_233_521 ();
 sky130_fd_sc_hd__decap_4 FILLER_233_530 ();
 sky130_fd_sc_hd__decap_4 FILLER_233_536 ();
 sky130_fd_sc_hd__decap_4 FILLER_233_542 ();
 sky130_fd_sc_hd__decap_4 FILLER_233_548 ();
 sky130_fd_sc_hd__decap_6 FILLER_233_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_233_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_233_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_233_576 ();
 sky130_fd_sc_hd__decap_4 FILLER_233_588 ();
 sky130_fd_sc_hd__decap_4 FILLER_233_594 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_233_612 ();
 sky130_fd_sc_hd__decap_6 FILLER_233_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_233_623 ();
 sky130_fd_sc_hd__decap_4 FILLER_233_644 ();
 sky130_fd_sc_hd__decap_4 FILLER_233_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_233_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_233_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_233_677 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_684 ();
 sky130_fd_sc_hd__decap_4 FILLER_233_696 ();
 sky130_fd_sc_hd__fill_1 FILLER_233_700 ();
 sky130_fd_sc_hd__decap_4 FILLER_233_707 ();
 sky130_fd_sc_hd__decap_4 FILLER_233_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_233_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_233_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_733 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_745 ();
 sky130_fd_sc_hd__decap_6 FILLER_233_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_233_763 ();
 sky130_fd_sc_hd__decap_6 FILLER_233_770 ();
 sky130_fd_sc_hd__fill_1 FILLER_233_776 ();
 sky130_fd_sc_hd__fill_2 FILLER_233_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_233_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_233_807 ();
 sky130_fd_sc_hd__decap_4 FILLER_233_815 ();
 sky130_fd_sc_hd__decap_4 FILLER_233_822 ();
 sky130_fd_sc_hd__decap_4 FILLER_233_829 ();
 sky130_fd_sc_hd__fill_1 FILLER_233_833 ();
 sky130_fd_sc_hd__fill_2 FILLER_233_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_233_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_234_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_234_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_234_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_234_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_234_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_234_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_234_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_457 ();
 sky130_fd_sc_hd__decap_3 FILLER_234_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_234_474 ();
 sky130_fd_sc_hd__decap_6 FILLER_234_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_234_486 ();
 sky130_fd_sc_hd__decap_4 FILLER_234_492 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_496 ();
 sky130_fd_sc_hd__decap_4 FILLER_234_504 ();
 sky130_fd_sc_hd__decap_6 FILLER_234_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_234_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_234_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_234_543 ();
 sky130_fd_sc_hd__decap_8 FILLER_234_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_557 ();
 sky130_fd_sc_hd__decap_4 FILLER_234_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_234_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_234_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_234_607 ();
 sky130_fd_sc_hd__decap_4 FILLER_234_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_234_619 ();
 sky130_fd_sc_hd__decap_6 FILLER_234_625 ();
 sky130_fd_sc_hd__decap_4 FILLER_234_634 ();
 sky130_fd_sc_hd__decap_4 FILLER_234_640 ();
 sky130_fd_sc_hd__decap_3 FILLER_234_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_234_665 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_671 ();
 sky130_fd_sc_hd__decap_8 FILLER_234_685 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_693 ();
 sky130_fd_sc_hd__decap_4 FILLER_234_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_234_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_234_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_234_712 ();
 sky130_fd_sc_hd__decap_4 FILLER_234_718 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_724 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_736 ();
 sky130_fd_sc_hd__decap_4 FILLER_234_748 ();
 sky130_fd_sc_hd__fill_2 FILLER_234_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_234_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_234_764 ();
 sky130_fd_sc_hd__fill_2 FILLER_234_772 ();
 sky130_fd_sc_hd__decap_4 FILLER_234_776 ();
 sky130_fd_sc_hd__decap_4 FILLER_234_783 ();
 sky130_fd_sc_hd__decap_4 FILLER_234_794 ();
 sky130_fd_sc_hd__decap_6 FILLER_234_806 ();
 sky130_fd_sc_hd__fill_2 FILLER_234_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_234_817 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_825 ();
 sky130_fd_sc_hd__decap_8 FILLER_234_828 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_836 ();
 sky130_fd_sc_hd__fill_2 FILLER_234_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_235_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_235_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_235_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_235_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_235_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_235_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_235_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_235_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_235_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_235_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_235_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_235_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_235_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_235_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_235_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_235_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_235_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_235_469 ();
 sky130_fd_sc_hd__decap_4 FILLER_235_491 ();
 sky130_fd_sc_hd__decap_6 FILLER_235_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_235_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_235_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_235_514 ();
 sky130_fd_sc_hd__fill_1 FILLER_235_520 ();
 sky130_fd_sc_hd__decap_6 FILLER_235_526 ();
 sky130_fd_sc_hd__fill_1 FILLER_235_532 ();
 sky130_fd_sc_hd__decap_4 FILLER_235_540 ();
 sky130_fd_sc_hd__decap_4 FILLER_235_546 ();
 sky130_fd_sc_hd__decap_4 FILLER_235_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_235_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_235_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_235_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_235_573 ();
 sky130_fd_sc_hd__decap_6 FILLER_235_583 ();
 sky130_fd_sc_hd__decap_4 FILLER_235_596 ();
 sky130_fd_sc_hd__decap_8 FILLER_235_602 ();
 sky130_fd_sc_hd__fill_1 FILLER_235_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_235_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_235_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_235_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_235_633 ();
 sky130_fd_sc_hd__decap_4 FILLER_235_639 ();
 sky130_fd_sc_hd__decap_4 FILLER_235_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_235_651 ();
 sky130_fd_sc_hd__decap_4 FILLER_235_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_235_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_235_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_235_677 ();
 sky130_fd_sc_hd__decap_6 FILLER_235_694 ();
 sky130_fd_sc_hd__fill_1 FILLER_235_700 ();
 sky130_fd_sc_hd__decap_4 FILLER_235_717 ();
 sky130_fd_sc_hd__decap_4 FILLER_235_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_235_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_765 ();
 sky130_fd_sc_hd__decap_3 FILLER_235_777 ();
 sky130_fd_sc_hd__fill_2 FILLER_235_782 ();
 sky130_fd_sc_hd__decap_4 FILLER_235_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_235_794 ();
 sky130_fd_sc_hd__decap_4 FILLER_235_800 ();
 sky130_fd_sc_hd__decap_4 FILLER_235_806 ();
 sky130_fd_sc_hd__decap_4 FILLER_235_812 ();
 sky130_fd_sc_hd__decap_4 FILLER_235_818 ();
 sky130_fd_sc_hd__decap_4 FILLER_235_824 ();
 sky130_fd_sc_hd__decap_4 FILLER_235_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_235_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_235_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_236_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_236_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_236_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_236_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_236_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_236_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_236_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_236_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_236_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_493 ();
 sky130_fd_sc_hd__decap_6 FILLER_236_511 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_517 ();
 sky130_fd_sc_hd__decap_6 FILLER_236_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_236_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_236_544 ();
 sky130_fd_sc_hd__decap_6 FILLER_236_550 ();
 sky130_fd_sc_hd__decap_4 FILLER_236_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_236_577 ();
 sky130_fd_sc_hd__decap_4 FILLER_236_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_236_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_236_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_236_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_236_605 ();
 sky130_fd_sc_hd__decap_4 FILLER_236_625 ();
 sky130_fd_sc_hd__decap_8 FILLER_236_631 ();
 sky130_fd_sc_hd__decap_3 FILLER_236_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_236_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_236_649 ();
 sky130_fd_sc_hd__decap_8 FILLER_236_655 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_663 ();
 sky130_fd_sc_hd__decap_4 FILLER_236_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_236_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_236_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_705 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_719 ();
 sky130_fd_sc_hd__decap_3 FILLER_236_731 ();
 sky130_fd_sc_hd__decap_4 FILLER_236_736 ();
 sky130_fd_sc_hd__decap_4 FILLER_236_745 ();
 sky130_fd_sc_hd__decap_4 FILLER_236_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_236_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_761 ();
 sky130_fd_sc_hd__decap_8 FILLER_236_773 ();
 sky130_fd_sc_hd__fill_2 FILLER_236_781 ();
 sky130_fd_sc_hd__decap_4 FILLER_236_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_236_791 ();
 sky130_fd_sc_hd__decap_4 FILLER_236_797 ();
 sky130_fd_sc_hd__decap_4 FILLER_236_803 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_807 ();
 sky130_fd_sc_hd__fill_2 FILLER_236_810 ();
 sky130_fd_sc_hd__decap_6 FILLER_236_813 ();
 sky130_fd_sc_hd__decap_6 FILLER_236_821 ();
 sky130_fd_sc_hd__decap_4 FILLER_236_830 ();
 sky130_fd_sc_hd__decap_4 FILLER_236_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_237_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_237_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_237_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_237_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_237_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_237_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_237_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_237_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_237_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_503 ();
 sky130_fd_sc_hd__decap_3 FILLER_237_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_237_510 ();
 sky130_fd_sc_hd__decap_8 FILLER_237_516 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_524 ();
 sky130_fd_sc_hd__decap_4 FILLER_237_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_237_539 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_237_546 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_237_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_237_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_237_565 ();
 sky130_fd_sc_hd__decap_8 FILLER_237_571 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_579 ();
 sky130_fd_sc_hd__decap_4 FILLER_237_588 ();
 sky130_fd_sc_hd__decap_4 FILLER_237_594 ();
 sky130_fd_sc_hd__decap_4 FILLER_237_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_237_606 ();
 sky130_fd_sc_hd__decap_4 FILLER_237_612 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_237_648 ();
 sky130_fd_sc_hd__decap_6 FILLER_237_654 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_660 ();
 sky130_fd_sc_hd__fill_2 FILLER_237_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_237_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_237_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_237_685 ();
 sky130_fd_sc_hd__decap_4 FILLER_237_689 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_237_725 ();
 sky130_fd_sc_hd__decap_6 FILLER_237_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_237_751 ();
 sky130_fd_sc_hd__decap_4 FILLER_237_758 ();
 sky130_fd_sc_hd__decap_4 FILLER_237_766 ();
 sky130_fd_sc_hd__decap_4 FILLER_237_772 ();
 sky130_fd_sc_hd__decap_6 FILLER_237_778 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_237_797 ();
 sky130_fd_sc_hd__decap_4 FILLER_237_805 ();
 sky130_fd_sc_hd__decap_4 FILLER_237_811 ();
 sky130_fd_sc_hd__decap_4 FILLER_237_817 ();
 sky130_fd_sc_hd__decap_6 FILLER_237_828 ();
 sky130_fd_sc_hd__fill_2 FILLER_237_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_238_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_238_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_238_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_238_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_238_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_238_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_238_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_445 ();
 sky130_fd_sc_hd__decap_6 FILLER_238_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_238_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_238_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_238_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_238_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_238_494 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_500 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_512 ();
 sky130_fd_sc_hd__decap_4 FILLER_238_515 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_519 ();
 sky130_fd_sc_hd__decap_4 FILLER_238_522 ();
 sky130_fd_sc_hd__decap_4 FILLER_238_528 ();
 sky130_fd_sc_hd__decap_4 FILLER_238_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_238_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_238_555 ();
 sky130_fd_sc_hd__decap_4 FILLER_238_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_238_567 ();
 sky130_fd_sc_hd__decap_4 FILLER_238_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_238_579 ();
 sky130_fd_sc_hd__decap_3 FILLER_238_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_238_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_238_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_238_603 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_609 ();
 sky130_fd_sc_hd__decap_8 FILLER_238_621 ();
 sky130_fd_sc_hd__decap_6 FILLER_238_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_238_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_238_653 ();
 sky130_fd_sc_hd__decap_8 FILLER_238_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_681 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_685 ();
 sky130_fd_sc_hd__decap_3 FILLER_238_697 ();
 sky130_fd_sc_hd__decap_8 FILLER_238_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_238_709 ();
 sky130_fd_sc_hd__decap_4 FILLER_238_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_238_722 ();
 sky130_fd_sc_hd__decap_8 FILLER_238_728 ();
 sky130_fd_sc_hd__decap_4 FILLER_238_742 ();
 sky130_fd_sc_hd__decap_6 FILLER_238_750 ();
 sky130_fd_sc_hd__decap_4 FILLER_238_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_761 ();
 sky130_fd_sc_hd__decap_4 FILLER_238_771 ();
 sky130_fd_sc_hd__decap_8 FILLER_238_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_238_790 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_794 ();
 sky130_fd_sc_hd__decap_4 FILLER_238_797 ();
 sky130_fd_sc_hd__fill_2 FILLER_238_810 ();
 sky130_fd_sc_hd__decap_4 FILLER_238_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_238_819 ();
 sky130_fd_sc_hd__decap_3 FILLER_238_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_239_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_239_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_239_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_239_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_239_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_239_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_239_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_239_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_239_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_239_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_239_480 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_484 ();
 sky130_fd_sc_hd__decap_4 FILLER_239_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_239_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_503 ();
 sky130_fd_sc_hd__decap_6 FILLER_239_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_239_525 ();
 sky130_fd_sc_hd__decap_4 FILLER_239_536 ();
 sky130_fd_sc_hd__decap_4 FILLER_239_542 ();
 sky130_fd_sc_hd__decap_4 FILLER_239_548 ();
 sky130_fd_sc_hd__decap_6 FILLER_239_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_239_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_239_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_239_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_239_577 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_581 ();
 sky130_fd_sc_hd__decap_4 FILLER_239_590 ();
 sky130_fd_sc_hd__decap_6 FILLER_239_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_239_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_239_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_239_632 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_636 ();
 sky130_fd_sc_hd__decap_4 FILLER_239_639 ();
 sky130_fd_sc_hd__decap_4 FILLER_239_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_239_651 ();
 sky130_fd_sc_hd__decap_4 FILLER_239_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_661 ();
 sky130_fd_sc_hd__decap_6 FILLER_239_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_239_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_677 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_689 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_239_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_239_724 ();
 sky130_fd_sc_hd__fill_2 FILLER_239_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_239_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_751 ();
 sky130_fd_sc_hd__decap_8 FILLER_239_758 ();
 sky130_fd_sc_hd__fill_2 FILLER_239_782 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_239_797 ();
 sky130_fd_sc_hd__decap_4 FILLER_239_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_811 ();
 sky130_fd_sc_hd__decap_4 FILLER_239_814 ();
 sky130_fd_sc_hd__fill_2 FILLER_239_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_240_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_240_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_240_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_240_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_240_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_240_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_240_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_445 ();
 sky130_fd_sc_hd__decap_8 FILLER_240_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_240_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_240_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_240_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_240_497 ();
 sky130_fd_sc_hd__decap_4 FILLER_240_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_240_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_240_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_240_521 ();
 sky130_fd_sc_hd__decap_4 FILLER_240_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_240_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_240_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_240_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_240_549 ();
 sky130_fd_sc_hd__decap_4 FILLER_240_555 ();
 sky130_fd_sc_hd__decap_4 FILLER_240_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_579 ();
 sky130_fd_sc_hd__decap_6 FILLER_240_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_240_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_240_594 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_600 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_612 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_624 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_636 ();
 sky130_fd_sc_hd__decap_4 FILLER_240_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_240_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_240_649 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_655 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_667 ();
 sky130_fd_sc_hd__decap_4 FILLER_240_679 ();
 sky130_fd_sc_hd__decap_4 FILLER_240_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_240_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_240_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_240_705 ();
 sky130_fd_sc_hd__decap_6 FILLER_240_712 ();
 sky130_fd_sc_hd__decap_4 FILLER_240_720 ();
 sky130_fd_sc_hd__decap_4 FILLER_240_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_240_733 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_737 ();
 sky130_fd_sc_hd__decap_8 FILLER_240_742 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_750 ();
 sky130_fd_sc_hd__fill_2 FILLER_240_754 ();
 sky130_fd_sc_hd__decap_3 FILLER_240_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_240_765 ();
 sky130_fd_sc_hd__decap_4 FILLER_240_774 ();
 sky130_fd_sc_hd__decap_4 FILLER_240_782 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_790 ();
 sky130_fd_sc_hd__decap_3 FILLER_240_802 ();
 sky130_fd_sc_hd__fill_2 FILLER_240_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_240_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_240_818 ();
 sky130_fd_sc_hd__decap_4 FILLER_240_829 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_833 ();
 sky130_fd_sc_hd__decap_4 FILLER_240_838 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_241_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_241_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_241_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_241_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_241_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_241_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_241_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_241_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_241_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_241_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_241_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_241_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_241_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_241_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_241_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_241_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_241_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_241_467 ();
 sky130_fd_sc_hd__decap_4 FILLER_241_470 ();
 sky130_fd_sc_hd__decap_4 FILLER_241_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_241_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_241_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_241_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_241_517 ();
 sky130_fd_sc_hd__decap_6 FILLER_241_523 ();
 sky130_fd_sc_hd__decap_4 FILLER_241_535 ();
 sky130_fd_sc_hd__decap_4 FILLER_241_541 ();
 sky130_fd_sc_hd__decap_8 FILLER_241_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_241_555 ();
 sky130_fd_sc_hd__fill_2 FILLER_241_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_241_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_241_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_241_577 ();
 sky130_fd_sc_hd__decap_6 FILLER_241_583 ();
 sky130_fd_sc_hd__decap_4 FILLER_241_591 ();
 sky130_fd_sc_hd__decap_4 FILLER_241_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_241_603 ();
 sky130_fd_sc_hd__decap_6 FILLER_241_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_241_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_241_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_621 ();
 sky130_fd_sc_hd__fill_1 FILLER_241_633 ();
 sky130_fd_sc_hd__decap_4 FILLER_241_642 ();
 sky130_fd_sc_hd__decap_4 FILLER_241_663 ();
 sky130_fd_sc_hd__decap_3 FILLER_241_669 ();
 sky130_fd_sc_hd__decap_8 FILLER_241_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_241_700 ();
 sky130_fd_sc_hd__decap_4 FILLER_241_720 ();
 sky130_fd_sc_hd__fill_2 FILLER_241_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_241_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_241_737 ();
 sky130_fd_sc_hd__decap_4 FILLER_241_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_241_761 ();
 sky130_fd_sc_hd__decap_4 FILLER_241_768 ();
 sky130_fd_sc_hd__decap_6 FILLER_241_778 ();
 sky130_fd_sc_hd__fill_2 FILLER_241_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_241_789 ();
 sky130_fd_sc_hd__decap_3 FILLER_241_797 ();
 sky130_fd_sc_hd__decap_4 FILLER_241_802 ();
 sky130_fd_sc_hd__decap_8 FILLER_241_814 ();
 sky130_fd_sc_hd__fill_2 FILLER_241_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_241_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_242_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_242_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_242_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_242_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_242_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_242_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_242_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_242_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_242_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_242_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_242_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_242_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_242_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_242_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_242_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_457 ();
 sky130_fd_sc_hd__decap_3 FILLER_242_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_242_474 ();
 sky130_fd_sc_hd__decap_6 FILLER_242_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_242_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_242_492 ();
 sky130_fd_sc_hd__fill_1 FILLER_242_496 ();
 sky130_fd_sc_hd__decap_4 FILLER_242_499 ();
 sky130_fd_sc_hd__decap_4 FILLER_242_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_242_523 ();
 sky130_fd_sc_hd__decap_3 FILLER_242_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_242_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_242_551 ();
 sky130_fd_sc_hd__decap_4 FILLER_242_554 ();
 sky130_fd_sc_hd__decap_4 FILLER_242_572 ();
 sky130_fd_sc_hd__decap_6 FILLER_242_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_242_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_242_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_242_593 ();
 sky130_fd_sc_hd__decap_8 FILLER_242_599 ();
 sky130_fd_sc_hd__fill_1 FILLER_242_607 ();
 sky130_fd_sc_hd__decap_4 FILLER_242_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_242_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_242_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_242_649 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_655 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_667 ();
 sky130_fd_sc_hd__decap_6 FILLER_242_679 ();
 sky130_fd_sc_hd__fill_1 FILLER_242_685 ();
 sky130_fd_sc_hd__decap_8 FILLER_242_689 ();
 sky130_fd_sc_hd__decap_3 FILLER_242_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_242_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_705 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_717 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_242_753 ();
 sky130_fd_sc_hd__decap_4 FILLER_242_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_242_761 ();
 sky130_fd_sc_hd__decap_4 FILLER_242_765 ();
 sky130_fd_sc_hd__decap_8 FILLER_242_771 ();
 sky130_fd_sc_hd__decap_3 FILLER_242_779 ();
 sky130_fd_sc_hd__decap_4 FILLER_242_784 ();
 sky130_fd_sc_hd__decap_4 FILLER_242_797 ();
 sky130_fd_sc_hd__decap_3 FILLER_242_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_242_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_242_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_242_823 ();
 sky130_fd_sc_hd__fill_1 FILLER_242_827 ();
 sky130_fd_sc_hd__decap_4 FILLER_242_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_242_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_243_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_243_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_243_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_243_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_243_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_243_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_243_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_243_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_243_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_243_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_243_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_243_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_243_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_243_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_243_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_243_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_461 ();
 sky130_fd_sc_hd__decap_6 FILLER_243_473 ();
 sky130_fd_sc_hd__decap_8 FILLER_243_481 ();
 sky130_fd_sc_hd__decap_3 FILLER_243_489 ();
 sky130_fd_sc_hd__decap_8 FILLER_243_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_243_502 ();
 sky130_fd_sc_hd__decap_8 FILLER_243_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_243_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_243_518 ();
 sky130_fd_sc_hd__fill_1 FILLER_243_522 ();
 sky130_fd_sc_hd__decap_4 FILLER_243_525 ();
 sky130_fd_sc_hd__decap_8 FILLER_243_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_243_539 ();
 sky130_fd_sc_hd__decap_4 FILLER_243_542 ();
 sky130_fd_sc_hd__decap_8 FILLER_243_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_243_558 ();
 sky130_fd_sc_hd__decap_6 FILLER_243_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_243_575 ();
 sky130_fd_sc_hd__decap_4 FILLER_243_586 ();
 sky130_fd_sc_hd__decap_4 FILLER_243_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_243_603 ();
 sky130_fd_sc_hd__fill_1 FILLER_243_609 ();
 sky130_fd_sc_hd__decap_3 FILLER_243_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_243_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_243_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_243_633 ();
 sky130_fd_sc_hd__decap_6 FILLER_243_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_243_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_243_648 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_654 ();
 sky130_fd_sc_hd__decap_6 FILLER_243_666 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_243_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_243_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_765 ();
 sky130_fd_sc_hd__fill_2 FILLER_243_777 ();
 sky130_fd_sc_hd__decap_3 FILLER_243_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_243_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_243_791 ();
 sky130_fd_sc_hd__fill_1 FILLER_243_797 ();
 sky130_fd_sc_hd__decap_4 FILLER_243_806 ();
 sky130_fd_sc_hd__decap_6 FILLER_243_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_243_819 ();
 sky130_fd_sc_hd__decap_4 FILLER_243_822 ();
 sky130_fd_sc_hd__decap_6 FILLER_243_828 ();
 sky130_fd_sc_hd__fill_2 FILLER_243_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_243_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_244_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_244_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_244_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_244_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_244_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_244_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_244_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_244_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_244_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_244_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_244_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_244_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_244_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_244_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_244_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_244_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_244_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_489 ();
 sky130_fd_sc_hd__decap_8 FILLER_244_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_244_516 ();
 sky130_fd_sc_hd__decap_6 FILLER_244_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_244_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_244_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_244_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_244_543 ();
 sky130_fd_sc_hd__decap_8 FILLER_244_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_244_557 ();
 sky130_fd_sc_hd__decap_4 FILLER_244_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_244_576 ();
 sky130_fd_sc_hd__decap_6 FILLER_244_582 ();
 sky130_fd_sc_hd__decap_3 FILLER_244_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_244_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_244_605 ();
 sky130_fd_sc_hd__decap_4 FILLER_244_611 ();
 sky130_fd_sc_hd__decap_4 FILLER_244_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_244_623 ();
 sky130_fd_sc_hd__decap_4 FILLER_244_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_244_635 ();
 sky130_fd_sc_hd__decap_3 FILLER_244_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_244_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_244_649 ();
 sky130_fd_sc_hd__decap_4 FILLER_244_655 ();
 sky130_fd_sc_hd__decap_8 FILLER_244_661 ();
 sky130_fd_sc_hd__decap_4 FILLER_244_675 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_244_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_244_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_244_725 ();
 sky130_fd_sc_hd__decap_8 FILLER_244_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_244_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_244_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_244_769 ();
 sky130_fd_sc_hd__fill_1 FILLER_244_773 ();
 sky130_fd_sc_hd__decap_4 FILLER_244_777 ();
 sky130_fd_sc_hd__decap_4 FILLER_244_790 ();
 sky130_fd_sc_hd__decap_6 FILLER_244_799 ();
 sky130_fd_sc_hd__fill_1 FILLER_244_805 ();
 sky130_fd_sc_hd__decap_4 FILLER_244_808 ();
 sky130_fd_sc_hd__decap_4 FILLER_244_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_244_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_244_820 ();
 sky130_fd_sc_hd__decap_4 FILLER_244_826 ();
 sky130_fd_sc_hd__decap_4 FILLER_244_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_244_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_245_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_245_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_245_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_245_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_245_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_245_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_245_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_245_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_245_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_245_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_245_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_245_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_245_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_245_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_245_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_245_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_245_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_245_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_245_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_245_509 ();
 sky130_fd_sc_hd__decap_8 FILLER_245_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_245_527 ();
 sky130_fd_sc_hd__decap_6 FILLER_245_536 ();
 sky130_fd_sc_hd__decap_4 FILLER_245_550 ();
 sky130_fd_sc_hd__decap_4 FILLER_245_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_245_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_245_565 ();
 sky130_fd_sc_hd__decap_6 FILLER_245_574 ();
 sky130_fd_sc_hd__decap_6 FILLER_245_587 ();
 sky130_fd_sc_hd__decap_4 FILLER_245_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_245_605 ();
 sky130_fd_sc_hd__decap_4 FILLER_245_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_245_615 ();
 sky130_fd_sc_hd__decap_6 FILLER_245_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_245_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_245_635 ();
 sky130_fd_sc_hd__decap_4 FILLER_245_644 ();
 sky130_fd_sc_hd__decap_6 FILLER_245_650 ();
 sky130_fd_sc_hd__decap_4 FILLER_245_659 ();
 sky130_fd_sc_hd__decap_6 FILLER_245_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_245_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_245_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_245_677 ();
 sky130_fd_sc_hd__fill_1 FILLER_245_681 ();
 sky130_fd_sc_hd__decap_4 FILLER_245_684 ();
 sky130_fd_sc_hd__decap_8 FILLER_245_690 ();
 sky130_fd_sc_hd__decap_8 FILLER_245_700 ();
 sky130_fd_sc_hd__fill_1 FILLER_245_708 ();
 sky130_fd_sc_hd__decap_4 FILLER_245_712 ();
 sky130_fd_sc_hd__decap_3 FILLER_245_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_245_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_245_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_245_748 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_754 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_766 ();
 sky130_fd_sc_hd__decap_6 FILLER_245_778 ();
 sky130_fd_sc_hd__decap_4 FILLER_245_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_245_789 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_793 ();
 sky130_fd_sc_hd__decap_4 FILLER_245_805 ();
 sky130_fd_sc_hd__decap_4 FILLER_245_811 ();
 sky130_fd_sc_hd__decap_4 FILLER_245_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_245_823 ();
 sky130_fd_sc_hd__fill_1 FILLER_245_827 ();
 sky130_fd_sc_hd__decap_4 FILLER_245_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_245_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_245_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_246_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_246_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_246_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_246_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_246_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_246_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_246_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_246_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_246_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_246_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_246_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_246_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_246_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_246_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_246_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_246_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_246_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_246_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_246_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_246_516 ();
 sky130_fd_sc_hd__fill_2 FILLER_246_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_246_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_246_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_246_551 ();
 sky130_fd_sc_hd__decap_4 FILLER_246_557 ();
 sky130_fd_sc_hd__decap_4 FILLER_246_563 ();
 sky130_fd_sc_hd__decap_4 FILLER_246_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_246_575 ();
 sky130_fd_sc_hd__decap_6 FILLER_246_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_246_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_246_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_246_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_246_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_246_605 ();
 sky130_fd_sc_hd__decap_4 FILLER_246_611 ();
 sky130_fd_sc_hd__decap_8 FILLER_246_621 ();
 sky130_fd_sc_hd__fill_1 FILLER_246_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_246_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_246_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_246_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_246_650 ();
 sky130_fd_sc_hd__fill_1 FILLER_246_658 ();
 sky130_fd_sc_hd__decap_4 FILLER_246_668 ();
 sky130_fd_sc_hd__fill_1 FILLER_246_672 ();
 sky130_fd_sc_hd__decap_6 FILLER_246_682 ();
 sky130_fd_sc_hd__fill_1 FILLER_246_688 ();
 sky130_fd_sc_hd__fill_2 FILLER_246_698 ();
 sky130_fd_sc_hd__decap_3 FILLER_246_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_246_720 ();
 sky130_fd_sc_hd__decap_6 FILLER_246_727 ();
 sky130_fd_sc_hd__decap_6 FILLER_246_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_246_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_246_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_761 ();
 sky130_fd_sc_hd__decap_4 FILLER_246_773 ();
 sky130_fd_sc_hd__fill_1 FILLER_246_777 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_246_797 ();
 sky130_fd_sc_hd__decap_4 FILLER_246_803 ();
 sky130_fd_sc_hd__fill_2 FILLER_246_810 ();
 sky130_fd_sc_hd__decap_6 FILLER_246_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_246_826 ();
 sky130_fd_sc_hd__fill_2 FILLER_246_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_247_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_247_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_247_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_247_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_247_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_247_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_247_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_247_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_247_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_247_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_247_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_247_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_247_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_247_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_247_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_247_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_247_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_247_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_247_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_247_487 ();
 sky130_fd_sc_hd__decap_8 FILLER_247_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_247_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_247_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_247_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_247_512 ();
 sky130_fd_sc_hd__decap_4 FILLER_247_524 ();
 sky130_fd_sc_hd__fill_1 FILLER_247_528 ();
 sky130_fd_sc_hd__decap_4 FILLER_247_538 ();
 sky130_fd_sc_hd__decap_4 FILLER_247_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_247_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_247_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_247_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_247_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_247_577 ();
 sky130_fd_sc_hd__decap_4 FILLER_247_583 ();
 sky130_fd_sc_hd__decap_8 FILLER_247_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_247_603 ();
 sky130_fd_sc_hd__decap_6 FILLER_247_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_247_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_247_621 ();
 sky130_fd_sc_hd__fill_1 FILLER_247_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_247_647 ();
 sky130_fd_sc_hd__decap_4 FILLER_247_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_247_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_247_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_247_700 ();
 sky130_fd_sc_hd__decap_4 FILLER_247_706 ();
 sky130_fd_sc_hd__fill_1 FILLER_247_710 ();
 sky130_fd_sc_hd__decap_4 FILLER_247_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_247_720 ();
 sky130_fd_sc_hd__fill_2 FILLER_247_726 ();
 sky130_fd_sc_hd__decap_6 FILLER_247_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_247_735 ();
 sky130_fd_sc_hd__decap_4 FILLER_247_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_247_746 ();
 sky130_fd_sc_hd__decap_6 FILLER_247_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_247_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_247_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_247_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_247_801 ();
 sky130_fd_sc_hd__decap_6 FILLER_247_805 ();
 sky130_fd_sc_hd__decap_4 FILLER_247_818 ();
 sky130_fd_sc_hd__fill_2 FILLER_247_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_247_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_248_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_248_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_248_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_248_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_248_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_248_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_248_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_248_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_248_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_248_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_248_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_248_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_248_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_248_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_248_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_248_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_248_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_248_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_248_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_248_507 ();
 sky130_fd_sc_hd__decap_6 FILLER_248_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_248_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_248_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_248_540 ();
 sky130_fd_sc_hd__decap_4 FILLER_248_554 ();
 sky130_fd_sc_hd__decap_4 FILLER_248_564 ();
 sky130_fd_sc_hd__decap_4 FILLER_248_574 ();
 sky130_fd_sc_hd__decap_4 FILLER_248_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_248_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_248_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_248_605 ();
 sky130_fd_sc_hd__decap_4 FILLER_248_614 ();
 sky130_fd_sc_hd__decap_8 FILLER_248_620 ();
 sky130_fd_sc_hd__decap_4 FILLER_248_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_248_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_248_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_248_666 ();
 sky130_fd_sc_hd__fill_1 FILLER_248_674 ();
 sky130_fd_sc_hd__decap_4 FILLER_248_684 ();
 sky130_fd_sc_hd__decap_4 FILLER_248_691 ();
 sky130_fd_sc_hd__decap_3 FILLER_248_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_725 ();
 sky130_fd_sc_hd__decap_4 FILLER_248_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_248_743 ();
 sky130_fd_sc_hd__fill_1 FILLER_248_749 ();
 sky130_fd_sc_hd__decap_3 FILLER_248_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_248_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_248_768 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_774 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_786 ();
 sky130_fd_sc_hd__decap_3 FILLER_248_798 ();
 sky130_fd_sc_hd__decap_4 FILLER_248_803 ();
 sky130_fd_sc_hd__decap_3 FILLER_248_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_248_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_248_817 ();
 sky130_fd_sc_hd__fill_1 FILLER_248_821 ();
 sky130_fd_sc_hd__decap_4 FILLER_248_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_248_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_248_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_249_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_249_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_249_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_249_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_249_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_249_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_249_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_249_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_249_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_249_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_249_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_249_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_249_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_249_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_249_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_249_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_249_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_249_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_249_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_249_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_249_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_249_521 ();
 sky130_fd_sc_hd__decap_4 FILLER_249_527 ();
 sky130_fd_sc_hd__decap_4 FILLER_249_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_249_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_249_546 ();
 sky130_fd_sc_hd__decap_4 FILLER_249_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_249_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_249_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_249_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_249_576 ();
 sky130_fd_sc_hd__decap_4 FILLER_249_582 ();
 sky130_fd_sc_hd__decap_4 FILLER_249_588 ();
 sky130_fd_sc_hd__decap_4 FILLER_249_594 ();
 sky130_fd_sc_hd__fill_2 FILLER_249_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_249_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_249_621 ();
 sky130_fd_sc_hd__decap_8 FILLER_249_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_249_638 ();
 sky130_fd_sc_hd__decap_4 FILLER_249_644 ();
 sky130_fd_sc_hd__decap_4 FILLER_249_650 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_656 ();
 sky130_fd_sc_hd__fill_2 FILLER_249_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_249_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_249_691 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_249_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_249_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_249_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_735 ();
 sky130_fd_sc_hd__fill_1 FILLER_249_747 ();
 sky130_fd_sc_hd__decap_4 FILLER_249_750 ();
 sky130_fd_sc_hd__fill_1 FILLER_249_754 ();
 sky130_fd_sc_hd__decap_4 FILLER_249_758 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_764 ();
 sky130_fd_sc_hd__fill_1 FILLER_249_776 ();
 sky130_fd_sc_hd__decap_4 FILLER_249_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_249_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_785 ();
 sky130_fd_sc_hd__decap_3 FILLER_249_797 ();
 sky130_fd_sc_hd__decap_4 FILLER_249_806 ();
 sky130_fd_sc_hd__decap_4 FILLER_249_812 ();
 sky130_fd_sc_hd__fill_1 FILLER_249_816 ();
 sky130_fd_sc_hd__decap_6 FILLER_249_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_249_839 ();
 sky130_fd_sc_hd__fill_1 FILLER_249_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_250_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_250_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_250_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_250_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_250_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_250_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_250_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_250_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_250_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_250_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_250_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_250_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_250_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_250_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_250_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_250_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_250_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_250_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_250_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_250_494 ();
 sky130_fd_sc_hd__decap_4 FILLER_250_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_506 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_250_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_250_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_250_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_250_543 ();
 sky130_fd_sc_hd__decap_6 FILLER_250_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_250_555 ();
 sky130_fd_sc_hd__decap_4 FILLER_250_558 ();
 sky130_fd_sc_hd__decap_8 FILLER_250_570 ();
 sky130_fd_sc_hd__fill_2 FILLER_250_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_250_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_250_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_250_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_250_605 ();
 sky130_fd_sc_hd__decap_4 FILLER_250_611 ();
 sky130_fd_sc_hd__decap_4 FILLER_250_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_623 ();
 sky130_fd_sc_hd__fill_1 FILLER_250_635 ();
 sky130_fd_sc_hd__decap_6 FILLER_250_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_250_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_250_649 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_655 ();
 sky130_fd_sc_hd__decap_6 FILLER_250_667 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_676 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_688 ();
 sky130_fd_sc_hd__decap_4 FILLER_250_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_250_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_250_711 ();
 sky130_fd_sc_hd__fill_1 FILLER_250_715 ();
 sky130_fd_sc_hd__decap_4 FILLER_250_718 ();
 sky130_fd_sc_hd__fill_1 FILLER_250_722 ();
 sky130_fd_sc_hd__decap_4 FILLER_250_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_250_735 ();
 sky130_fd_sc_hd__decap_8 FILLER_250_741 ();
 sky130_fd_sc_hd__fill_2 FILLER_250_749 ();
 sky130_fd_sc_hd__fill_2 FILLER_250_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_250_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_250_775 ();
 sky130_fd_sc_hd__decap_4 FILLER_250_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_250_795 ();
 sky130_fd_sc_hd__decap_6 FILLER_250_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_250_811 ();
 sky130_fd_sc_hd__decap_4 FILLER_250_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_250_819 ();
 sky130_fd_sc_hd__decap_4 FILLER_250_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_250_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_250_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_251_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_251_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_251_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_251_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_251_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_251_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_251_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_251_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_251_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_251_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_251_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_251_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_251_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_251_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_251_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_251_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_251_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_251_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_251_495 ();
 sky130_fd_sc_hd__decap_3 FILLER_251_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_529 ();
 sky130_fd_sc_hd__decap_4 FILLER_251_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_251_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_251_548 ();
 sky130_fd_sc_hd__decap_6 FILLER_251_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_251_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_251_579 ();
 sky130_fd_sc_hd__decap_4 FILLER_251_599 ();
 sky130_fd_sc_hd__decap_6 FILLER_251_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_251_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_251_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_251_633 ();
 sky130_fd_sc_hd__fill_1 FILLER_251_637 ();
 sky130_fd_sc_hd__decap_4 FILLER_251_640 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_646 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_251_670 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_685 ();
 sky130_fd_sc_hd__decap_3 FILLER_251_697 ();
 sky130_fd_sc_hd__decap_4 FILLER_251_706 ();
 sky130_fd_sc_hd__decap_4 FILLER_251_716 ();
 sky130_fd_sc_hd__decap_6 FILLER_251_722 ();
 sky130_fd_sc_hd__decap_6 FILLER_251_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_737 ();
 sky130_fd_sc_hd__decap_8 FILLER_251_749 ();
 sky130_fd_sc_hd__decap_8 FILLER_251_759 ();
 sky130_fd_sc_hd__decap_8 FILLER_251_773 ();
 sky130_fd_sc_hd__decap_3 FILLER_251_781 ();
 sky130_fd_sc_hd__decap_8 FILLER_251_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_251_793 ();
 sky130_fd_sc_hd__decap_8 FILLER_251_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_807 ();
 sky130_fd_sc_hd__decap_8 FILLER_251_819 ();
 sky130_fd_sc_hd__decap_4 FILLER_251_829 ();
 sky130_fd_sc_hd__fill_1 FILLER_251_833 ();
 sky130_fd_sc_hd__fill_2 FILLER_251_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_251_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_252_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_252_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_252_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_252_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_252_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_252_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_252_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_252_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_252_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_252_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_252_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_252_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_252_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_252_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_252_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_252_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_252_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_252_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_252_492 ();
 sky130_fd_sc_hd__decap_4 FILLER_252_512 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_252_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_252_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_252_549 ();
 sky130_fd_sc_hd__decap_8 FILLER_252_552 ();
 sky130_fd_sc_hd__fill_1 FILLER_252_560 ();
 sky130_fd_sc_hd__decap_6 FILLER_252_564 ();
 sky130_fd_sc_hd__fill_1 FILLER_252_570 ();
 sky130_fd_sc_hd__decap_4 FILLER_252_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_252_579 ();
 sky130_fd_sc_hd__decap_3 FILLER_252_585 ();
 sky130_fd_sc_hd__decap_6 FILLER_252_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_252_595 ();
 sky130_fd_sc_hd__decap_4 FILLER_252_602 ();
 sky130_fd_sc_hd__decap_4 FILLER_252_608 ();
 sky130_fd_sc_hd__decap_6 FILLER_252_614 ();
 sky130_fd_sc_hd__decap_4 FILLER_252_622 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_628 ();
 sky130_fd_sc_hd__decap_4 FILLER_252_640 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_252_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_252_665 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_670 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_682 ();
 sky130_fd_sc_hd__decap_6 FILLER_252_694 ();
 sky130_fd_sc_hd__decap_4 FILLER_252_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_252_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_252_708 ();
 sky130_fd_sc_hd__decap_4 FILLER_252_714 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_720 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_732 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_744 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_252_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_252_776 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_782 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_794 ();
 sky130_fd_sc_hd__decap_6 FILLER_252_806 ();
 sky130_fd_sc_hd__decap_4 FILLER_252_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_252_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_252_820 ();
 sky130_fd_sc_hd__decap_4 FILLER_252_826 ();
 sky130_fd_sc_hd__decap_4 FILLER_252_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_252_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_253_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_253_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_253_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_253_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_253_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_253_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_253_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_253_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_253_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_253_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_253_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_253_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_253_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_253_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_253_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_253_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_473 ();
 sky130_fd_sc_hd__decap_8 FILLER_253_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_253_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_253_502 ();
 sky130_fd_sc_hd__decap_6 FILLER_253_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_253_514 ();
 sky130_fd_sc_hd__decap_4 FILLER_253_520 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_538 ();
 sky130_fd_sc_hd__decap_8 FILLER_253_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_253_558 ();
 sky130_fd_sc_hd__decap_3 FILLER_253_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_253_566 ();
 sky130_fd_sc_hd__decap_4 FILLER_253_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_253_578 ();
 sky130_fd_sc_hd__decap_4 FILLER_253_584 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_590 ();
 sky130_fd_sc_hd__decap_4 FILLER_253_604 ();
 sky130_fd_sc_hd__decap_6 FILLER_253_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_253_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_253_622 ();
 sky130_fd_sc_hd__decap_4 FILLER_253_628 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_634 ();
 sky130_fd_sc_hd__decap_4 FILLER_253_646 ();
 sky130_fd_sc_hd__decap_4 FILLER_253_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_253_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_253_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_253_700 ();
 sky130_fd_sc_hd__decap_4 FILLER_253_706 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_712 ();
 sky130_fd_sc_hd__decap_4 FILLER_253_724 ();
 sky130_fd_sc_hd__fill_2 FILLER_253_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_733 ();
 sky130_fd_sc_hd__decap_3 FILLER_253_745 ();
 sky130_fd_sc_hd__decap_4 FILLER_253_750 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_756 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_768 ();
 sky130_fd_sc_hd__decap_4 FILLER_253_780 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_797 ();
 sky130_fd_sc_hd__decap_4 FILLER_253_809 ();
 sky130_fd_sc_hd__decap_6 FILLER_253_816 ();
 sky130_fd_sc_hd__decap_4 FILLER_253_824 ();
 sky130_fd_sc_hd__decap_4 FILLER_253_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_253_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_253_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_254_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_254_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_254_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_254_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_254_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_254_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_254_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_254_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_254_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_254_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_254_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_254_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_254_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_254_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_254_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_254_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_254_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_254_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_254_496 ();
 sky130_fd_sc_hd__decap_4 FILLER_254_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_254_508 ();
 sky130_fd_sc_hd__decap_4 FILLER_254_520 ();
 sky130_fd_sc_hd__decap_6 FILLER_254_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_254_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_254_553 ();
 sky130_fd_sc_hd__decap_4 FILLER_254_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_564 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_576 ();
 sky130_fd_sc_hd__decap_8 FILLER_254_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_254_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_254_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_254_608 ();
 sky130_fd_sc_hd__decap_4 FILLER_254_620 ();
 sky130_fd_sc_hd__decap_4 FILLER_254_632 ();
 sky130_fd_sc_hd__decap_6 FILLER_254_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_254_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_254_666 ();
 sky130_fd_sc_hd__decap_4 FILLER_254_679 ();
 sky130_fd_sc_hd__decap_4 FILLER_254_685 ();
 sky130_fd_sc_hd__decap_4 FILLER_254_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_254_695 ();
 sky130_fd_sc_hd__fill_2 FILLER_254_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_254_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_254_722 ();
 sky130_fd_sc_hd__decap_4 FILLER_254_734 ();
 sky130_fd_sc_hd__fill_1 FILLER_254_738 ();
 sky130_fd_sc_hd__decap_4 FILLER_254_746 ();
 sky130_fd_sc_hd__decap_4 FILLER_254_752 ();
 sky130_fd_sc_hd__fill_2 FILLER_254_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_761 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_773 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_254_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_254_803 ();
 sky130_fd_sc_hd__decap_6 FILLER_254_806 ();
 sky130_fd_sc_hd__decap_3 FILLER_254_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_254_818 ();
 sky130_fd_sc_hd__decap_4 FILLER_254_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_254_838 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_255_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_255_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_255_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_255_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_255_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_255_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_255_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_255_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_255_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_255_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_255_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_255_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_255_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_255_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_255_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_255_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_255_497 ();
 sky130_fd_sc_hd__decap_4 FILLER_255_500 ();
 sky130_fd_sc_hd__decap_4 FILLER_255_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_255_525 ();
 sky130_fd_sc_hd__decap_4 FILLER_255_531 ();
 sky130_fd_sc_hd__decap_8 FILLER_255_537 ();
 sky130_fd_sc_hd__decap_3 FILLER_255_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_255_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_255_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_255_566 ();
 sky130_fd_sc_hd__decap_4 FILLER_255_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_255_578 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_584 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_596 ();
 sky130_fd_sc_hd__fill_2 FILLER_255_608 ();
 sky130_fd_sc_hd__decap_4 FILLER_255_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_255_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_255_635 ();
 sky130_fd_sc_hd__decap_4 FILLER_255_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_647 ();
 sky130_fd_sc_hd__decap_6 FILLER_255_659 ();
 sky130_fd_sc_hd__fill_1 FILLER_255_665 ();
 sky130_fd_sc_hd__decap_3 FILLER_255_669 ();
 sky130_fd_sc_hd__decap_8 FILLER_255_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_255_681 ();
 sky130_fd_sc_hd__decap_8 FILLER_255_702 ();
 sky130_fd_sc_hd__decap_4 FILLER_255_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_255_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_255_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_255_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_255_750 ();
 sky130_fd_sc_hd__decap_4 FILLER_255_759 ();
 sky130_fd_sc_hd__decap_4 FILLER_255_765 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_771 ();
 sky130_fd_sc_hd__fill_1 FILLER_255_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_255_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_255_791 ();
 sky130_fd_sc_hd__fill_1 FILLER_255_799 ();
 sky130_fd_sc_hd__decap_4 FILLER_255_806 ();
 sky130_fd_sc_hd__decap_8 FILLER_255_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_255_821 ();
 sky130_fd_sc_hd__fill_2 FILLER_255_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_255_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_256_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_256_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_256_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_256_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_256_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_256_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_256_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_256_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_256_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_256_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_256_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_256_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_256_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_256_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_256_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_256_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_256_475 ();
 sky130_fd_sc_hd__decap_6 FILLER_256_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_256_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_256_492 ();
 sky130_fd_sc_hd__decap_4 FILLER_256_498 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_504 ();
 sky130_fd_sc_hd__fill_1 FILLER_256_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_256_519 ();
 sky130_fd_sc_hd__decap_6 FILLER_256_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_256_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_256_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_256_545 ();
 sky130_fd_sc_hd__decap_6 FILLER_256_562 ();
 sky130_fd_sc_hd__decap_4 FILLER_256_576 ();
 sky130_fd_sc_hd__decap_6 FILLER_256_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_256_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_256_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_256_599 ();
 sky130_fd_sc_hd__decap_6 FILLER_256_605 ();
 sky130_fd_sc_hd__decap_4 FILLER_256_627 ();
 sky130_fd_sc_hd__decap_8 FILLER_256_633 ();
 sky130_fd_sc_hd__decap_3 FILLER_256_641 ();
 sky130_fd_sc_hd__decap_8 FILLER_256_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_256_653 ();
 sky130_fd_sc_hd__decap_4 FILLER_256_657 ();
 sky130_fd_sc_hd__decap_8 FILLER_256_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_256_685 ();
 sky130_fd_sc_hd__decap_8 FILLER_256_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_256_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_256_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_256_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_256_716 ();
 sky130_fd_sc_hd__decap_4 FILLER_256_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_256_741 ();
 sky130_fd_sc_hd__decap_4 FILLER_256_752 ();
 sky130_fd_sc_hd__fill_2 FILLER_256_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_256_761 ();
 sky130_fd_sc_hd__fill_1 FILLER_256_767 ();
 sky130_fd_sc_hd__decap_4 FILLER_256_772 ();
 sky130_fd_sc_hd__decap_4 FILLER_256_784 ();
 sky130_fd_sc_hd__decap_4 FILLER_256_790 ();
 sky130_fd_sc_hd__fill_1 FILLER_256_794 ();
 sky130_fd_sc_hd__decap_4 FILLER_256_804 ();
 sky130_fd_sc_hd__fill_2 FILLER_256_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_256_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_256_822 ();
 sky130_fd_sc_hd__fill_1 FILLER_256_826 ();
 sky130_fd_sc_hd__decap_6 FILLER_256_836 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_257_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_257_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_257_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_257_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_257_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_257_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_257_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_257_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_257_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_257_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_257_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_257_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_257_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_257_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_257_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_257_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_461 ();
 sky130_fd_sc_hd__decap_6 FILLER_257_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_257_479 ();
 sky130_fd_sc_hd__decap_4 FILLER_257_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_257_502 ();
 sky130_fd_sc_hd__decap_8 FILLER_257_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_257_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_257_522 ();
 sky130_fd_sc_hd__decap_8 FILLER_257_542 ();
 sky130_fd_sc_hd__decap_6 FILLER_257_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_257_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_257_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_257_565 ();
 sky130_fd_sc_hd__decap_6 FILLER_257_585 ();
 sky130_fd_sc_hd__decap_4 FILLER_257_599 ();
 sky130_fd_sc_hd__decap_8 FILLER_257_605 ();
 sky130_fd_sc_hd__decap_3 FILLER_257_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_257_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_257_625 ();
 sky130_fd_sc_hd__decap_4 FILLER_257_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_257_633 ();
 sky130_fd_sc_hd__decap_4 FILLER_257_653 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_659 ();
 sky130_fd_sc_hd__fill_1 FILLER_257_671 ();
 sky130_fd_sc_hd__decap_8 FILLER_257_673 ();
 sky130_fd_sc_hd__decap_3 FILLER_257_681 ();
 sky130_fd_sc_hd__decap_4 FILLER_257_686 ();
 sky130_fd_sc_hd__decap_4 FILLER_257_699 ();
 sky130_fd_sc_hd__decap_8 FILLER_257_705 ();
 sky130_fd_sc_hd__fill_1 FILLER_257_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_257_716 ();
 sky130_fd_sc_hd__decap_3 FILLER_257_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_257_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_257_738 ();
 sky130_fd_sc_hd__decap_4 FILLER_257_749 ();
 sky130_fd_sc_hd__decap_4 FILLER_257_762 ();
 sky130_fd_sc_hd__decap_4 FILLER_257_768 ();
 sky130_fd_sc_hd__fill_1 FILLER_257_772 ();
 sky130_fd_sc_hd__fill_2 FILLER_257_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_257_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_257_790 ();
 sky130_fd_sc_hd__decap_4 FILLER_257_804 ();
 sky130_fd_sc_hd__decap_4 FILLER_257_816 ();
 sky130_fd_sc_hd__decap_6 FILLER_257_828 ();
 sky130_fd_sc_hd__fill_2 FILLER_257_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_257_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_258_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_258_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_258_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_258_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_258_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_258_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_258_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_258_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_258_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_258_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_258_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_258_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_258_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_258_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_258_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_258_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_258_475 ();
 sky130_fd_sc_hd__decap_6 FILLER_258_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_258_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_258_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_258_493 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_499 ();
 sky130_fd_sc_hd__decap_8 FILLER_258_511 ();
 sky130_fd_sc_hd__decap_3 FILLER_258_519 ();
 sky130_fd_sc_hd__decap_4 FILLER_258_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_258_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_258_545 ();
 sky130_fd_sc_hd__decap_8 FILLER_258_555 ();
 sky130_fd_sc_hd__decap_3 FILLER_258_563 ();
 sky130_fd_sc_hd__decap_4 FILLER_258_568 ();
 sky130_fd_sc_hd__decap_8 FILLER_258_574 ();
 sky130_fd_sc_hd__fill_1 FILLER_258_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_258_586 ();
 sky130_fd_sc_hd__decap_4 FILLER_258_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_258_609 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_627 ();
 sky130_fd_sc_hd__fill_2 FILLER_258_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_258_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_258_656 ();
 sky130_fd_sc_hd__decap_6 FILLER_258_662 ();
 sky130_fd_sc_hd__decap_4 FILLER_258_674 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_680 ();
 sky130_fd_sc_hd__decap_8 FILLER_258_692 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_701 ();
 sky130_fd_sc_hd__decap_3 FILLER_258_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_258_718 ();
 sky130_fd_sc_hd__decap_4 FILLER_258_729 ();
 sky130_fd_sc_hd__decap_3 FILLER_258_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_258_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_258_768 ();
 sky130_fd_sc_hd__fill_1 FILLER_258_776 ();
 sky130_fd_sc_hd__decap_4 FILLER_258_784 ();
 sky130_fd_sc_hd__decap_4 FILLER_258_796 ();
 sky130_fd_sc_hd__decap_6 FILLER_258_806 ();
 sky130_fd_sc_hd__fill_2 FILLER_258_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_258_819 ();
 sky130_fd_sc_hd__decap_4 FILLER_258_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_258_829 ();
 sky130_fd_sc_hd__decap_4 FILLER_258_833 ();
 sky130_fd_sc_hd__fill_2 FILLER_258_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_259_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_259_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_259_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_259_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_259_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_259_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_259_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_259_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_259_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_259_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_259_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_259_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_259_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_259_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_259_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_259_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_259_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_259_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_259_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_509 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_521 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_259_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_259_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_259_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_259_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_259_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_259_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_259_576 ();
 sky130_fd_sc_hd__decap_4 FILLER_259_583 ();
 sky130_fd_sc_hd__decap_4 FILLER_259_603 ();
 sky130_fd_sc_hd__decap_6 FILLER_259_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_259_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_259_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_259_650 ();
 sky130_fd_sc_hd__decap_4 FILLER_259_656 ();
 sky130_fd_sc_hd__decap_8 FILLER_259_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_259_670 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_259_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_259_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_259_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_259_733 ();
 sky130_fd_sc_hd__fill_1 FILLER_259_737 ();
 sky130_fd_sc_hd__decap_4 FILLER_259_740 ();
 sky130_fd_sc_hd__decap_4 FILLER_259_746 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_766 ();
 sky130_fd_sc_hd__fill_2 FILLER_259_778 ();
 sky130_fd_sc_hd__fill_2 FILLER_259_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_259_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_259_789 ();
 sky130_fd_sc_hd__decap_4 FILLER_259_795 ();
 sky130_fd_sc_hd__decap_4 FILLER_259_805 ();
 sky130_fd_sc_hd__decap_4 FILLER_259_815 ();
 sky130_fd_sc_hd__decap_6 FILLER_259_821 ();
 sky130_fd_sc_hd__fill_1 FILLER_259_827 ();
 sky130_fd_sc_hd__fill_2 FILLER_259_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_259_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_260_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_260_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_260_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_260_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_260_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_260_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_260_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_260_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_260_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_260_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_260_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_260_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_260_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_260_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_260_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_260_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_260_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_260_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_260_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_260_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_260_494 ();
 sky130_fd_sc_hd__decap_4 FILLER_260_500 ();
 sky130_fd_sc_hd__decap_4 FILLER_260_506 ();
 sky130_fd_sc_hd__decap_4 FILLER_260_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_260_519 ();
 sky130_fd_sc_hd__decap_6 FILLER_260_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_260_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_260_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_260_549 ();
 sky130_fd_sc_hd__decap_6 FILLER_260_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_260_559 ();
 sky130_fd_sc_hd__decap_4 FILLER_260_563 ();
 sky130_fd_sc_hd__decap_4 FILLER_260_569 ();
 sky130_fd_sc_hd__decap_8 FILLER_260_575 ();
 sky130_fd_sc_hd__decap_3 FILLER_260_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_260_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_260_599 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_605 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_260_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_260_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_260_650 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_658 ();
 sky130_fd_sc_hd__fill_1 FILLER_260_670 ();
 sky130_fd_sc_hd__decap_6 FILLER_260_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_260_681 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_260_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_737 ();
 sky130_fd_sc_hd__fill_2 FILLER_260_749 ();
 sky130_fd_sc_hd__fill_2 FILLER_260_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_260_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_761 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_773 ();
 sky130_fd_sc_hd__fill_1 FILLER_260_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_260_788 ();
 sky130_fd_sc_hd__decap_8 FILLER_260_798 ();
 sky130_fd_sc_hd__decap_4 FILLER_260_808 ();
 sky130_fd_sc_hd__decap_4 FILLER_260_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_260_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_260_820 ();
 sky130_fd_sc_hd__decap_4 FILLER_260_826 ();
 sky130_fd_sc_hd__fill_2 FILLER_260_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_261_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_261_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_261_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_261_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_261_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_261_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_261_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_261_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_261_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_261_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_261_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_261_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_261_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_261_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_261_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_261_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_261_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_261_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_261_486 ();
 sky130_fd_sc_hd__decap_6 FILLER_261_498 ();
 sky130_fd_sc_hd__decap_6 FILLER_261_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_261_511 ();
 sky130_fd_sc_hd__decap_6 FILLER_261_520 ();
 sky130_fd_sc_hd__fill_1 FILLER_261_526 ();
 sky130_fd_sc_hd__decap_4 FILLER_261_530 ();
 sky130_fd_sc_hd__decap_4 FILLER_261_536 ();
 sky130_fd_sc_hd__decap_6 FILLER_261_542 ();
 sky130_fd_sc_hd__fill_1 FILLER_261_548 ();
 sky130_fd_sc_hd__decap_3 FILLER_261_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_261_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_261_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_261_577 ();
 sky130_fd_sc_hd__decap_4 FILLER_261_583 ();
 sky130_fd_sc_hd__decap_4 FILLER_261_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_595 ();
 sky130_fd_sc_hd__decap_8 FILLER_261_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_261_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_261_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_261_637 ();
 sky130_fd_sc_hd__decap_4 FILLER_261_656 ();
 sky130_fd_sc_hd__decap_3 FILLER_261_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_261_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_261_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_261_687 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_693 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_705 ();
 sky130_fd_sc_hd__decap_6 FILLER_261_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_261_723 ();
 sky130_fd_sc_hd__fill_2 FILLER_261_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_261_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_733 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_745 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_769 ();
 sky130_fd_sc_hd__decap_3 FILLER_261_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_261_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_261_803 ();
 sky130_fd_sc_hd__decap_4 FILLER_261_806 ();
 sky130_fd_sc_hd__decap_4 FILLER_261_812 ();
 sky130_fd_sc_hd__decap_4 FILLER_261_818 ();
 sky130_fd_sc_hd__decap_4 FILLER_261_824 ();
 sky130_fd_sc_hd__decap_4 FILLER_261_831 ();
 sky130_fd_sc_hd__fill_2 FILLER_261_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_261_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_262_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_262_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_262_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_262_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_262_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_262_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_262_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_262_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_262_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_262_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_262_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_262_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_262_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_262_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_262_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_262_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_262_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_262_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_262_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_262_504 ();
 sky130_fd_sc_hd__decap_4 FILLER_262_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_262_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_262_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_262_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_262_563 ();
 sky130_fd_sc_hd__decap_4 FILLER_262_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_262_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_262_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_593 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_605 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_262_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_262_669 ();
 sky130_fd_sc_hd__decap_4 FILLER_262_679 ();
 sky130_fd_sc_hd__decap_6 FILLER_262_686 ();
 sky130_fd_sc_hd__decap_4 FILLER_262_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_262_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_262_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_262_712 ();
 sky130_fd_sc_hd__decap_4 FILLER_262_718 ();
 sky130_fd_sc_hd__decap_8 FILLER_262_724 ();
 sky130_fd_sc_hd__decap_4 FILLER_262_738 ();
 sky130_fd_sc_hd__decap_4 FILLER_262_744 ();
 sky130_fd_sc_hd__decap_6 FILLER_262_750 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_262_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_262_773 ();
 sky130_fd_sc_hd__fill_1 FILLER_262_777 ();
 sky130_fd_sc_hd__decap_8 FILLER_262_798 ();
 sky130_fd_sc_hd__fill_2 FILLER_262_806 ();
 sky130_fd_sc_hd__fill_2 FILLER_262_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_262_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_262_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_262_823 ();
 sky130_fd_sc_hd__decap_6 FILLER_262_836 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_263_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_263_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_263_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_263_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_263_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_263_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_263_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_263_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_263_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_263_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_263_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_263_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_263_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_263_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_263_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_263_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_263_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_263_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_263_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_509 ();
 sky130_fd_sc_hd__fill_1 FILLER_263_521 ();
 sky130_fd_sc_hd__decap_4 FILLER_263_524 ();
 sky130_fd_sc_hd__decap_4 FILLER_263_544 ();
 sky130_fd_sc_hd__decap_8 FILLER_263_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_263_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_263_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_263_565 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_571 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_583 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_595 ();
 sky130_fd_sc_hd__decap_8 FILLER_263_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_263_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_641 ();
 sky130_fd_sc_hd__decap_8 FILLER_263_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_263_661 ();
 sky130_fd_sc_hd__decap_6 FILLER_263_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_263_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_263_691 ();
 sky130_fd_sc_hd__decap_4 FILLER_263_711 ();
 sky130_fd_sc_hd__decap_4 FILLER_263_724 ();
 sky130_fd_sc_hd__decap_6 FILLER_263_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_263_735 ();
 sky130_fd_sc_hd__decap_4 FILLER_263_744 ();
 sky130_fd_sc_hd__decap_4 FILLER_263_752 ();
 sky130_fd_sc_hd__decap_4 FILLER_263_758 ();
 sky130_fd_sc_hd__decap_8 FILLER_263_764 ();
 sky130_fd_sc_hd__fill_1 FILLER_263_772 ();
 sky130_fd_sc_hd__fill_2 FILLER_263_782 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_797 ();
 sky130_fd_sc_hd__decap_3 FILLER_263_809 ();
 sky130_fd_sc_hd__decap_4 FILLER_263_814 ();
 sky130_fd_sc_hd__decap_4 FILLER_263_827 ();
 sky130_fd_sc_hd__decap_6 FILLER_263_834 ();
 sky130_fd_sc_hd__fill_1 FILLER_263_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_264_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_264_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_264_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_264_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_264_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_264_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_264_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_264_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_264_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_264_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_264_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_264_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_264_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_264_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_264_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_264_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_264_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_264_525 ();
 sky130_fd_sc_hd__decap_4 FILLER_264_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_264_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_264_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_264_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_593 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_605 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_264_641 ();
 sky130_fd_sc_hd__decap_4 FILLER_264_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_264_651 ();
 sky130_fd_sc_hd__decap_8 FILLER_264_674 ();
 sky130_fd_sc_hd__decap_4 FILLER_264_691 ();
 sky130_fd_sc_hd__decap_3 FILLER_264_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_264_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_264_722 ();
 sky130_fd_sc_hd__decap_4 FILLER_264_731 ();
 sky130_fd_sc_hd__decap_4 FILLER_264_737 ();
 sky130_fd_sc_hd__decap_4 FILLER_264_743 ();
 sky130_fd_sc_hd__fill_1 FILLER_264_747 ();
 sky130_fd_sc_hd__fill_2 FILLER_264_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_264_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_264_765 ();
 sky130_fd_sc_hd__fill_1 FILLER_264_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_264_773 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_786 ();
 sky130_fd_sc_hd__decap_3 FILLER_264_798 ();
 sky130_fd_sc_hd__fill_2 FILLER_264_810 ();
 sky130_fd_sc_hd__decap_4 FILLER_264_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_264_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_264_820 ();
 sky130_fd_sc_hd__fill_2 FILLER_264_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_265_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_265_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_265_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_265_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_265_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_265_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_265_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_265_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_265_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_265_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_265_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_265_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_265_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_265_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_265_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_265_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_265_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_265_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_265_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_265_527 ();
 sky130_fd_sc_hd__decap_4 FILLER_265_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_265_540 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_265_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_265_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_265_565 ();
 sky130_fd_sc_hd__decap_6 FILLER_265_568 ();
 sky130_fd_sc_hd__decap_4 FILLER_265_576 ();
 sky130_fd_sc_hd__decap_4 FILLER_265_582 ();
 sky130_fd_sc_hd__decap_4 FILLER_265_594 ();
 sky130_fd_sc_hd__decap_4 FILLER_265_600 ();
 sky130_fd_sc_hd__decap_8 FILLER_265_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_265_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_265_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_265_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_265_685 ();
 sky130_fd_sc_hd__decap_4 FILLER_265_693 ();
 sky130_fd_sc_hd__decap_4 FILLER_265_699 ();
 sky130_fd_sc_hd__decap_4 FILLER_265_706 ();
 sky130_fd_sc_hd__fill_2 FILLER_265_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_265_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_265_734 ();
 sky130_fd_sc_hd__fill_2 FILLER_265_742 ();
 sky130_fd_sc_hd__decap_4 FILLER_265_746 ();
 sky130_fd_sc_hd__decap_4 FILLER_265_754 ();
 sky130_fd_sc_hd__decap_6 FILLER_265_760 ();
 sky130_fd_sc_hd__fill_2 FILLER_265_782 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_265_797 ();
 sky130_fd_sc_hd__decap_4 FILLER_265_800 ();
 sky130_fd_sc_hd__decap_4 FILLER_265_808 ();
 sky130_fd_sc_hd__fill_1 FILLER_265_812 ();
 sky130_fd_sc_hd__decap_4 FILLER_265_829 ();
 sky130_fd_sc_hd__decap_4 FILLER_265_836 ();
 sky130_fd_sc_hd__fill_1 FILLER_265_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_266_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_266_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_266_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_266_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_266_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_266_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_266_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_266_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_266_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_266_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_266_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_266_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_266_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_266_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_266_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_266_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_266_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_266_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_266_497 ();
 sky130_fd_sc_hd__decap_4 FILLER_266_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_266_508 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_514 ();
 sky130_fd_sc_hd__decap_6 FILLER_266_526 ();
 sky130_fd_sc_hd__decap_4 FILLER_266_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_266_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_266_546 ();
 sky130_fd_sc_hd__decap_4 FILLER_266_552 ();
 sky130_fd_sc_hd__decap_6 FILLER_266_558 ();
 sky130_fd_sc_hd__fill_1 FILLER_266_564 ();
 sky130_fd_sc_hd__decap_4 FILLER_266_567 ();
 sky130_fd_sc_hd__decap_8 FILLER_266_574 ();
 sky130_fd_sc_hd__fill_1 FILLER_266_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_266_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_266_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_266_607 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_266_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_266_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_266_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_266_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_266_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_266_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_266_732 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_738 ();
 sky130_fd_sc_hd__decap_6 FILLER_266_750 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_781 ();
 sky130_fd_sc_hd__decap_6 FILLER_266_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_266_799 ();
 sky130_fd_sc_hd__decap_4 FILLER_266_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_266_811 ();
 sky130_fd_sc_hd__decap_8 FILLER_266_813 ();
 sky130_fd_sc_hd__decap_6 FILLER_266_830 ();
 sky130_fd_sc_hd__fill_1 FILLER_266_836 ();
 sky130_fd_sc_hd__fill_2 FILLER_266_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_267_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_267_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_267_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_267_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_267_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_267_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_267_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_267_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_267_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_267_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_267_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_267_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_267_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_267_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_267_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_267_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_267_497 ();
 sky130_fd_sc_hd__decap_4 FILLER_267_500 ();
 sky130_fd_sc_hd__decap_4 FILLER_267_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_267_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_267_518 ();
 sky130_fd_sc_hd__decap_4 FILLER_267_524 ();
 sky130_fd_sc_hd__decap_8 FILLER_267_530 ();
 sky130_fd_sc_hd__decap_6 FILLER_267_554 ();
 sky130_fd_sc_hd__decap_6 FILLER_267_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_267_567 ();
 sky130_fd_sc_hd__decap_4 FILLER_267_576 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_596 ();
 sky130_fd_sc_hd__decap_8 FILLER_267_608 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_641 ();
 sky130_fd_sc_hd__fill_1 FILLER_267_653 ();
 sky130_fd_sc_hd__decap_8 FILLER_267_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_267_665 ();
 sky130_fd_sc_hd__fill_2 FILLER_267_670 ();
 sky130_fd_sc_hd__decap_6 FILLER_267_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_681 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_693 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_705 ();
 sky130_fd_sc_hd__decap_8 FILLER_267_717 ();
 sky130_fd_sc_hd__decap_3 FILLER_267_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_267_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_267_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_809 ();
 sky130_fd_sc_hd__fill_1 FILLER_267_821 ();
 sky130_fd_sc_hd__decap_4 FILLER_267_824 ();
 sky130_fd_sc_hd__decap_4 FILLER_267_831 ();
 sky130_fd_sc_hd__fill_2 FILLER_267_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_267_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_268_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_268_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_268_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_268_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_268_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_268_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_268_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_268_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_268_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_268_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_268_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_268_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_268_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_268_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_268_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_268_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_268_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_268_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_268_498 ();
 sky130_fd_sc_hd__fill_1 FILLER_268_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_268_506 ();
 sky130_fd_sc_hd__decap_6 FILLER_268_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_268_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_268_537 ();
 sky130_fd_sc_hd__decap_8 FILLER_268_543 ();
 sky130_fd_sc_hd__decap_3 FILLER_268_551 ();
 sky130_fd_sc_hd__decap_4 FILLER_268_556 ();
 sky130_fd_sc_hd__decap_4 FILLER_268_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_268_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_625 ();
 sky130_fd_sc_hd__decap_3 FILLER_268_637 ();
 sky130_fd_sc_hd__fill_2 FILLER_268_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_268_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_268_666 ();
 sky130_fd_sc_hd__decap_4 FILLER_268_679 ();
 sky130_fd_sc_hd__decap_4 FILLER_268_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_268_698 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_725 ();
 sky130_fd_sc_hd__decap_6 FILLER_268_737 ();
 sky130_fd_sc_hd__decap_8 FILLER_268_745 ();
 sky130_fd_sc_hd__decap_3 FILLER_268_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_268_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_765 ();
 sky130_fd_sc_hd__decap_8 FILLER_268_786 ();
 sky130_fd_sc_hd__fill_2 FILLER_268_794 ();
 sky130_fd_sc_hd__decap_4 FILLER_268_798 ();
 sky130_fd_sc_hd__decap_4 FILLER_268_808 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_268_827 ();
 sky130_fd_sc_hd__decap_4 FILLER_268_833 ();
 sky130_fd_sc_hd__fill_2 FILLER_268_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_269_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_269_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_269_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_269_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_269_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_269_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_269_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_269_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_269_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_269_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_269_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_269_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_269_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_269_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_269_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_269_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_269_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_269_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_269_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_269_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_269_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_269_519 ();
 sky130_fd_sc_hd__decap_4 FILLER_269_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_269_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_269_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_269_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_269_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_269_572 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_580 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_592 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_604 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_269_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_269_671 ();
 sky130_fd_sc_hd__decap_3 FILLER_269_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_269_679 ();
 sky130_fd_sc_hd__fill_1 FILLER_269_683 ();
 sky130_fd_sc_hd__decap_4 FILLER_269_686 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_710 ();
 sky130_fd_sc_hd__decap_6 FILLER_269_722 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_269_741 ();
 sky130_fd_sc_hd__decap_4 FILLER_269_745 ();
 sky130_fd_sc_hd__decap_4 FILLER_269_758 ();
 sky130_fd_sc_hd__decap_8 FILLER_269_764 ();
 sky130_fd_sc_hd__fill_1 FILLER_269_772 ();
 sky130_fd_sc_hd__fill_2 FILLER_269_782 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_269_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_269_801 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_811 ();
 sky130_fd_sc_hd__decap_6 FILLER_269_823 ();
 sky130_fd_sc_hd__decap_4 FILLER_269_831 ();
 sky130_fd_sc_hd__fill_2 FILLER_269_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_269_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_270_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_270_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_270_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_270_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_270_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_270_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_270_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_270_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_270_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_270_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_270_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_270_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_270_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_270_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_270_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_270_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_270_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_270_492 ();
 sky130_fd_sc_hd__decap_4 FILLER_270_498 ();
 sky130_fd_sc_hd__decap_6 FILLER_270_504 ();
 sky130_fd_sc_hd__decap_4 FILLER_270_518 ();
 sky130_fd_sc_hd__decap_4 FILLER_270_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_270_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_270_547 ();
 sky130_fd_sc_hd__fill_2 FILLER_270_555 ();
 sky130_fd_sc_hd__decap_4 FILLER_270_559 ();
 sky130_fd_sc_hd__decap_4 FILLER_270_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_270_571 ();
 sky130_fd_sc_hd__decap_8 FILLER_270_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_270_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_270_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_270_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_270_669 ();
 sky130_fd_sc_hd__decap_4 FILLER_270_687 ();
 sky130_fd_sc_hd__decap_6 FILLER_270_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_270_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_270_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_270_717 ();
 sky130_fd_sc_hd__decap_4 FILLER_270_730 ();
 sky130_fd_sc_hd__decap_8 FILLER_270_736 ();
 sky130_fd_sc_hd__fill_1 FILLER_270_744 ();
 sky130_fd_sc_hd__fill_2 FILLER_270_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_270_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_270_765 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_776 ();
 sky130_fd_sc_hd__decap_6 FILLER_270_788 ();
 sky130_fd_sc_hd__fill_2 FILLER_270_810 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_270_827 ();
 sky130_fd_sc_hd__decap_4 FILLER_270_833 ();
 sky130_fd_sc_hd__fill_2 FILLER_270_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_271_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_271_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_271_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_271_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_271_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_271_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_271_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_271_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_271_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_271_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_271_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_271_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_271_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_271_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_271_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_271_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_473 ();
 sky130_fd_sc_hd__decap_8 FILLER_271_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_271_493 ();
 sky130_fd_sc_hd__decap_8 FILLER_271_496 ();
 sky130_fd_sc_hd__decap_4 FILLER_271_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_271_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_531 ();
 sky130_fd_sc_hd__decap_8 FILLER_271_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_271_553 ();
 sky130_fd_sc_hd__decap_3 FILLER_271_557 ();
 sky130_fd_sc_hd__decap_3 FILLER_271_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_271_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_271_571 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_588 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_271_612 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_271_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_271_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_271_697 ();
 sky130_fd_sc_hd__decap_6 FILLER_271_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_271_707 ();
 sky130_fd_sc_hd__decap_4 FILLER_271_717 ();
 sky130_fd_sc_hd__decap_4 FILLER_271_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_271_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_271_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_271_734 ();
 sky130_fd_sc_hd__fill_1 FILLER_271_742 ();
 sky130_fd_sc_hd__decap_6 FILLER_271_759 ();
 sky130_fd_sc_hd__fill_1 FILLER_271_765 ();
 sky130_fd_sc_hd__fill_2 FILLER_271_782 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_785 ();
 sky130_fd_sc_hd__decap_3 FILLER_271_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_803 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_815 ();
 sky130_fd_sc_hd__fill_1 FILLER_271_827 ();
 sky130_fd_sc_hd__decap_3 FILLER_271_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_271_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_272_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_272_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_272_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_272_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_272_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_272_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_272_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_272_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_272_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_272_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_272_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_272_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_272_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_272_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_272_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_272_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_272_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_513 ();
 sky130_fd_sc_hd__decap_3 FILLER_272_525 ();
 sky130_fd_sc_hd__fill_2 FILLER_272_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_272_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_272_543 ();
 sky130_fd_sc_hd__fill_1 FILLER_272_551 ();
 sky130_fd_sc_hd__decap_4 FILLER_272_568 ();
 sky130_fd_sc_hd__decap_4 FILLER_272_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_272_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_272_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_593 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_605 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_272_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_669 ();
 sky130_fd_sc_hd__decap_8 FILLER_272_681 ();
 sky130_fd_sc_hd__fill_1 FILLER_272_689 ();
 sky130_fd_sc_hd__decap_6 FILLER_272_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_272_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_272_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_272_712 ();
 sky130_fd_sc_hd__fill_1 FILLER_272_716 ();
 sky130_fd_sc_hd__decap_4 FILLER_272_720 ();
 sky130_fd_sc_hd__decap_4 FILLER_272_743 ();
 sky130_fd_sc_hd__decap_6 FILLER_272_750 ();
 sky130_fd_sc_hd__fill_2 FILLER_272_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_761 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_773 ();
 sky130_fd_sc_hd__fill_2 FILLER_272_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_789 ();
 sky130_fd_sc_hd__decap_8 FILLER_272_801 ();
 sky130_fd_sc_hd__decap_3 FILLER_272_809 ();
 sky130_fd_sc_hd__decap_4 FILLER_272_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_272_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_272_820 ();
 sky130_fd_sc_hd__decap_4 FILLER_272_833 ();
 sky130_fd_sc_hd__fill_2 FILLER_272_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_273_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_273_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_273_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_273_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_273_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_273_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_273_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_273_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_273_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_273_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_273_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_273_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_273_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_273_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_273_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_273_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_273_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_273_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_273_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_273_510 ();
 sky130_fd_sc_hd__decap_4 FILLER_273_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_273_522 ();
 sky130_fd_sc_hd__decap_4 FILLER_273_529 ();
 sky130_fd_sc_hd__decap_6 FILLER_273_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_273_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_273_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_273_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_273_577 ();
 sky130_fd_sc_hd__decap_4 FILLER_273_583 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_273_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_273_641 ();
 sky130_fd_sc_hd__fill_1 FILLER_273_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_648 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_660 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_273_704 ();
 sky130_fd_sc_hd__decap_4 FILLER_273_724 ();
 sky130_fd_sc_hd__fill_2 FILLER_273_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_273_740 ();
 sky130_fd_sc_hd__decap_4 FILLER_273_749 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_767 ();
 sky130_fd_sc_hd__decap_4 FILLER_273_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_273_783 ();
 sky130_fd_sc_hd__decap_4 FILLER_273_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_798 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_273_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_273_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_274_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_274_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_274_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_274_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_274_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_274_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_274_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_274_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_274_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_274_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_274_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_274_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_274_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_274_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_274_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_274_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_274_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_489 ();
 sky130_fd_sc_hd__decap_6 FILLER_274_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_274_507 ();
 sky130_fd_sc_hd__decap_4 FILLER_274_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_274_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_274_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_274_527 ();
 sky130_fd_sc_hd__fill_2 FILLER_274_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_274_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_537 ();
 sky130_fd_sc_hd__decap_3 FILLER_274_549 ();
 sky130_fd_sc_hd__decap_4 FILLER_274_554 ();
 sky130_fd_sc_hd__decap_8 FILLER_274_560 ();
 sky130_fd_sc_hd__decap_4 FILLER_274_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_274_577 ();
 sky130_fd_sc_hd__decap_4 FILLER_274_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_274_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_274_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_274_643 ();
 sky130_fd_sc_hd__decap_3 FILLER_274_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_274_667 ();
 sky130_fd_sc_hd__decap_4 FILLER_274_674 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_680 ();
 sky130_fd_sc_hd__decap_8 FILLER_274_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_274_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_274_706 ();
 sky130_fd_sc_hd__fill_1 FILLER_274_714 ();
 sky130_fd_sc_hd__decap_6 FILLER_274_731 ();
 sky130_fd_sc_hd__fill_1 FILLER_274_737 ();
 sky130_fd_sc_hd__fill_2 FILLER_274_754 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_274_781 ();
 sky130_fd_sc_hd__decap_4 FILLER_274_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_274_798 ();
 sky130_fd_sc_hd__fill_1 FILLER_274_804 ();
 sky130_fd_sc_hd__decap_4 FILLER_274_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_274_811 ();
 sky130_fd_sc_hd__decap_6 FILLER_274_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_274_819 ();
 sky130_fd_sc_hd__decap_4 FILLER_274_822 ();
 sky130_fd_sc_hd__decap_8 FILLER_274_829 ();
 sky130_fd_sc_hd__fill_2 FILLER_274_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_275_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_275_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_275_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_275_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_275_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_275_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_275_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_275_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_275_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_275_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_275_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_275_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_275_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_275_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_275_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_275_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_275_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_275_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_275_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_275_559 ();
 sky130_fd_sc_hd__decap_4 FILLER_275_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_275_565 ();
 sky130_fd_sc_hd__decap_8 FILLER_275_568 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_592 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_604 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_641 ();
 sky130_fd_sc_hd__fill_1 FILLER_275_653 ();
 sky130_fd_sc_hd__decap_4 FILLER_275_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_275_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_275_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_275_684 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_275_702 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_706 ();
 sky130_fd_sc_hd__decap_6 FILLER_275_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_275_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_275_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_275_733 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_739 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_751 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_763 ();
 sky130_fd_sc_hd__decap_4 FILLER_275_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_275_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_275_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_275_803 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_811 ();
 sky130_fd_sc_hd__decap_4 FILLER_275_823 ();
 sky130_fd_sc_hd__fill_1 FILLER_275_827 ();
 sky130_fd_sc_hd__fill_2 FILLER_275_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_275_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_276_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_276_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_276_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_276_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_276_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_276_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_276_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_276_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_276_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_276_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_276_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_276_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_276_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_276_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_276_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_276_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_276_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_501 ();
 sky130_fd_sc_hd__decap_8 FILLER_276_513 ();
 sky130_fd_sc_hd__decap_8 FILLER_276_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_276_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_545 ();
 sky130_fd_sc_hd__decap_8 FILLER_276_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_276_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_276_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_276_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_276_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_276_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_593 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_605 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_276_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_276_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_276_677 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_683 ();
 sky130_fd_sc_hd__decap_4 FILLER_276_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_276_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_276_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_276_755 ();
 sky130_fd_sc_hd__decap_4 FILLER_276_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_276_761 ();
 sky130_fd_sc_hd__decap_4 FILLER_276_764 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_774 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_786 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_798 ();
 sky130_fd_sc_hd__fill_2 FILLER_276_810 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_813 ();
 sky130_fd_sc_hd__decap_6 FILLER_276_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_276_833 ();
 sky130_fd_sc_hd__fill_2 FILLER_276_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_277_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_277_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_277_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_277_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_277_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_277_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_277_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_277_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_277_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_277_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_277_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_277_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_277_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_277_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_277_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_277_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_277_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_277_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_277_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_277_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_277_523 ();
 sky130_fd_sc_hd__decap_4 FILLER_277_529 ();
 sky130_fd_sc_hd__decap_4 FILLER_277_535 ();
 sky130_fd_sc_hd__decap_6 FILLER_277_541 ();
 sky130_fd_sc_hd__decap_4 FILLER_277_549 ();
 sky130_fd_sc_hd__decap_4 FILLER_277_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_277_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_277_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_277_576 ();
 sky130_fd_sc_hd__fill_1 FILLER_277_580 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_583 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_595 ();
 sky130_fd_sc_hd__decap_8 FILLER_277_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_277_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_277_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_277_671 ();
 sky130_fd_sc_hd__decap_4 FILLER_277_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_679 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_691 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_703 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_715 ();
 sky130_fd_sc_hd__fill_1 FILLER_277_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_753 ();
 sky130_fd_sc_hd__decap_4 FILLER_277_765 ();
 sky130_fd_sc_hd__decap_8 FILLER_277_776 ();
 sky130_fd_sc_hd__fill_2 FILLER_277_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_277_807 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_818 ();
 sky130_fd_sc_hd__decap_6 FILLER_277_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_277_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_277_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_278_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_278_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_278_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_278_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_278_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_278_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_278_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_278_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_278_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_278_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_278_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_278_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_278_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_278_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_278_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_278_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_278_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_278_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_278_497 ();
 sky130_fd_sc_hd__decap_4 FILLER_278_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_278_514 ();
 sky130_fd_sc_hd__decap_6 FILLER_278_520 ();
 sky130_fd_sc_hd__fill_1 FILLER_278_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_278_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_278_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_278_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_278_549 ();
 sky130_fd_sc_hd__decap_4 FILLER_278_555 ();
 sky130_fd_sc_hd__decap_4 FILLER_278_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_278_567 ();
 sky130_fd_sc_hd__decap_8 FILLER_278_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_278_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_278_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_278_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_278_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_278_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_737 ();
 sky130_fd_sc_hd__decap_3 FILLER_278_749 ();
 sky130_fd_sc_hd__fill_2 FILLER_278_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_278_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_278_779 ();
 sky130_fd_sc_hd__decap_8 FILLER_278_789 ();
 sky130_fd_sc_hd__decap_3 FILLER_278_797 ();
 sky130_fd_sc_hd__decap_8 FILLER_278_802 ();
 sky130_fd_sc_hd__fill_2 FILLER_278_810 ();
 sky130_fd_sc_hd__decap_8 FILLER_278_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_278_821 ();
 sky130_fd_sc_hd__decap_4 FILLER_278_824 ();
 sky130_fd_sc_hd__fill_2 FILLER_278_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_279_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_279_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_279_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_279_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_279_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_279_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_279_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_279_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_279_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_279_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_279_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_279_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_279_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_279_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_279_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_279_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_279_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_279_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_279_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_279_525 ();
 sky130_fd_sc_hd__decap_4 FILLER_279_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_279_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_279_550 ();
 sky130_fd_sc_hd__decap_4 FILLER_279_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_279_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_279_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_279_577 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_583 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_595 ();
 sky130_fd_sc_hd__decap_8 FILLER_279_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_279_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_279_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_279_671 ();
 sky130_fd_sc_hd__decap_3 FILLER_279_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_678 ();
 sky130_fd_sc_hd__decap_8 FILLER_279_690 ();
 sky130_fd_sc_hd__decap_8 FILLER_279_701 ();
 sky130_fd_sc_hd__decap_3 FILLER_279_709 ();
 sky130_fd_sc_hd__decap_4 FILLER_279_714 ();
 sky130_fd_sc_hd__decap_4 FILLER_279_720 ();
 sky130_fd_sc_hd__fill_2 FILLER_279_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_279_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_279_740 ();
 sky130_fd_sc_hd__decap_8 FILLER_279_746 ();
 sky130_fd_sc_hd__decap_3 FILLER_279_754 ();
 sky130_fd_sc_hd__decap_4 FILLER_279_759 ();
 sky130_fd_sc_hd__decap_4 FILLER_279_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_279_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_279_783 ();
 sky130_fd_sc_hd__decap_4 FILLER_279_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_279_795 ();
 sky130_fd_sc_hd__fill_1 FILLER_279_801 ();
 sky130_fd_sc_hd__decap_6 FILLER_279_808 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_826 ();
 sky130_fd_sc_hd__fill_2 FILLER_279_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_279_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_280_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_280_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_280_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_280_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_280_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_280_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_280_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_280_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_280_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_280_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_280_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_280_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_280_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_280_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_280_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_280_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_280_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_280_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_280_520 ();
 sky130_fd_sc_hd__fill_1 FILLER_280_524 ();
 sky130_fd_sc_hd__decap_4 FILLER_280_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_280_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_280_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_280_551 ();
 sky130_fd_sc_hd__decap_4 FILLER_280_571 ();
 sky130_fd_sc_hd__decap_8 FILLER_280_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_280_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_280_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_280_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_280_669 ();
 sky130_fd_sc_hd__decap_4 FILLER_280_674 ();
 sky130_fd_sc_hd__decap_4 FILLER_280_687 ();
 sky130_fd_sc_hd__decap_6 FILLER_280_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_280_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_280_712 ();
 sky130_fd_sc_hd__decap_4 FILLER_280_721 ();
 sky130_fd_sc_hd__decap_4 FILLER_280_734 ();
 sky130_fd_sc_hd__decap_4 FILLER_280_741 ();
 sky130_fd_sc_hd__decap_4 FILLER_280_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_280_751 ();
 sky130_fd_sc_hd__fill_2 FILLER_280_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_280_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_280_768 ();
 sky130_fd_sc_hd__decap_4 FILLER_280_774 ();
 sky130_fd_sc_hd__fill_1 FILLER_280_778 ();
 sky130_fd_sc_hd__decap_4 FILLER_280_788 ();
 sky130_fd_sc_hd__decap_6 FILLER_280_794 ();
 sky130_fd_sc_hd__decap_3 FILLER_280_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_280_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_280_831 ();
 sky130_fd_sc_hd__decap_4 FILLER_280_838 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_281_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_281_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_281_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_281_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_281_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_281_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_281_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_281_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_281_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_281_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_281_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_281_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_281_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_281_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_281_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_281_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_281_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_281_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_281_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_522 ();
 sky130_fd_sc_hd__fill_1 FILLER_281_534 ();
 sky130_fd_sc_hd__decap_4 FILLER_281_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_281_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_281_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_281_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_281_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_281_671 ();
 sky130_fd_sc_hd__decap_4 FILLER_281_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_281_693 ();
 sky130_fd_sc_hd__decap_4 FILLER_281_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_281_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_281_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_281_747 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_758 ();
 sky130_fd_sc_hd__decap_3 FILLER_281_770 ();
 sky130_fd_sc_hd__fill_2 FILLER_281_782 ();
 sky130_fd_sc_hd__decap_8 FILLER_281_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_281_793 ();
 sky130_fd_sc_hd__decap_4 FILLER_281_810 ();
 sky130_fd_sc_hd__decap_4 FILLER_281_817 ();
 sky130_fd_sc_hd__fill_1 FILLER_281_821 ();
 sky130_fd_sc_hd__fill_2 FILLER_281_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_281_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_282_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_282_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_282_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_282_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_282_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_282_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_282_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_282_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_282_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_282_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_282_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_282_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_282_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_282_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_282_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_282_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_282_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_282_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_282_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_282_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_282_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_282_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_282_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_282_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_282_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_282_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_282_684 ();
 sky130_fd_sc_hd__decap_3 FILLER_282_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_282_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_282_705 ();
 sky130_fd_sc_hd__decap_6 FILLER_282_728 ();
 sky130_fd_sc_hd__fill_1 FILLER_282_734 ();
 sky130_fd_sc_hd__fill_2 FILLER_282_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_282_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_282_775 ();
 sky130_fd_sc_hd__decap_4 FILLER_282_795 ();
 sky130_fd_sc_hd__decap_8 FILLER_282_802 ();
 sky130_fd_sc_hd__fill_2 FILLER_282_810 ();
 sky130_fd_sc_hd__decap_4 FILLER_282_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_282_826 ();
 sky130_fd_sc_hd__fill_1 FILLER_282_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_282_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_283_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_283_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_283_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_283_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_283_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_283_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_283_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_283_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_283_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_283_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_283_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_283_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_283_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_283_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_283_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_283_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_283_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_283_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_283_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_283_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_283_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_283_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_283_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_283_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_283_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_283_678 ();
 sky130_fd_sc_hd__decap_6 FILLER_283_686 ();
 sky130_fd_sc_hd__fill_1 FILLER_283_692 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_283_707 ();
 sky130_fd_sc_hd__decap_4 FILLER_283_711 ();
 sky130_fd_sc_hd__decap_4 FILLER_283_717 ();
 sky130_fd_sc_hd__decap_4 FILLER_283_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_283_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_283_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_733 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_745 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_283_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_283_778 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_283_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_283_839 ();
 sky130_fd_sc_hd__fill_1 FILLER_283_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_284_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_284_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_284_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_284_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_284_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_284_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_284_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_284_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_284_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_284_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_284_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_284_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_284_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_284_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_284_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_284_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_284_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_284_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_284_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_284_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_284_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_284_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_284_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_284_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_284_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_284_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_284_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_284_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_284_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_284_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_284_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_285_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_285_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_285_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_285_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_285_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_285_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_285_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_285_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_285_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_285_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_285_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_285_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_285_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_285_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_285_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_285_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_285_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_285_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_285_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_285_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_285_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_285_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_285_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_285_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_685 ();
 sky130_fd_sc_hd__decap_3 FILLER_285_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_285_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_285_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_769 ();
 sky130_fd_sc_hd__decap_3 FILLER_285_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_797 ();
 sky130_fd_sc_hd__decap_3 FILLER_285_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_825 ();
 sky130_fd_sc_hd__decap_3 FILLER_285_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_285_841 ();
 assign o_mem_addr_high[7] = net212;
endmodule

