magic
tech sky130A
magscale 1 2
timestamp 1672446661
<< nwell >>
rect 1066 106885 108874 107451
rect 1066 105797 108874 106363
rect 1066 104709 108874 105275
rect 1066 103621 108874 104187
rect 1066 102533 108874 103099
rect 1066 101445 108874 102011
rect 1066 100357 108874 100923
rect 1066 99269 108874 99835
rect 1066 98181 108874 98747
rect 1066 97093 108874 97659
rect 1066 96005 108874 96571
rect 1066 94917 108874 95483
rect 1066 93829 108874 94395
rect 1066 92741 108874 93307
rect 1066 91653 108874 92219
rect 1066 90565 108874 91131
rect 1066 89477 108874 90043
rect 1066 88389 108874 88955
rect 1066 87301 108874 87867
rect 1066 86213 108874 86779
rect 1066 85125 108874 85691
rect 1066 84037 108874 84603
rect 1066 82949 108874 83515
rect 1066 81861 108874 82427
rect 1066 80773 108874 81339
rect 1066 79685 108874 80251
rect 1066 78597 108874 79163
rect 1066 77509 108874 78075
rect 1066 76421 108874 76987
rect 1066 75333 108874 75899
rect 1066 74245 108874 74811
rect 1066 73157 108874 73723
rect 1066 72069 108874 72635
rect 1066 70981 108874 71547
rect 1066 69893 108874 70459
rect 1066 68805 108874 69371
rect 1066 67717 108874 68283
rect 1066 66629 108874 67195
rect 1066 65541 108874 66107
rect 1066 64453 108874 65019
rect 1066 63365 108874 63931
rect 1066 62277 108874 62843
rect 1066 61189 108874 61755
rect 1066 60101 108874 60667
rect 1066 59013 108874 59579
rect 1066 57925 108874 58491
rect 1066 56837 108874 57403
rect 1066 55749 108874 56315
rect 1066 54661 108874 55227
rect 1066 53573 108874 54139
rect 1066 52485 108874 53051
rect 1066 51397 108874 51963
rect 1066 50309 108874 50875
rect 1066 49221 108874 49787
rect 1066 48133 108874 48699
rect 1066 47045 108874 47611
rect 1066 45957 108874 46523
rect 1066 44869 108874 45435
rect 1066 43781 108874 44347
rect 1066 42693 108874 43259
rect 1066 41605 108874 42171
rect 1066 40517 108874 41083
rect 1066 39429 108874 39995
rect 1066 38341 108874 38907
rect 1066 37253 108874 37819
rect 1066 36165 108874 36731
rect 1066 35077 108874 35643
rect 1066 33989 108874 34555
rect 1066 32901 108874 33467
rect 1066 31813 108874 32379
rect 1066 30725 108874 31291
rect 1066 29637 108874 30203
rect 1066 28549 108874 29115
rect 1066 27461 108874 28027
rect 1066 26373 108874 26939
rect 1066 25285 108874 25851
rect 1066 24197 108874 24763
rect 1066 23109 108874 23675
rect 1066 22021 108874 22587
rect 1066 20933 108874 21499
rect 1066 19845 108874 20411
rect 1066 18757 108874 19323
rect 1066 17669 108874 18235
rect 1066 16581 108874 17147
rect 1066 15493 108874 16059
rect 1066 14405 108874 14971
rect 1066 13317 108874 13883
rect 1066 12229 108874 12795
rect 1066 11141 108874 11707
rect 1066 10053 108874 10619
rect 1066 8965 108874 9531
rect 1066 7877 108874 8443
rect 1066 6789 108874 7355
rect 1066 5701 108874 6267
rect 1066 4613 108874 5179
rect 1066 3525 108874 4091
rect 1066 2437 108874 3003
<< obsli1 >>
rect 1104 2159 108836 107729
<< obsm1 >>
rect 1104 1844 109006 107760
<< obsm2 >>
rect 1584 1838 109000 107749
<< metal3 >>
rect 109200 106632 110000 106752
rect 109200 104048 110000 104168
rect 109200 101464 110000 101584
rect 109200 98880 110000 99000
rect 109200 96296 110000 96416
rect 109200 93712 110000 93832
rect 109200 91128 110000 91248
rect 109200 88544 110000 88664
rect 109200 85960 110000 86080
rect 109200 83376 110000 83496
rect 109200 80792 110000 80912
rect 109200 78208 110000 78328
rect 109200 75624 110000 75744
rect 109200 73040 110000 73160
rect 109200 70456 110000 70576
rect 109200 67872 110000 67992
rect 109200 65288 110000 65408
rect 109200 62704 110000 62824
rect 109200 60120 110000 60240
rect 109200 57536 110000 57656
rect 109200 54952 110000 55072
rect 109200 52368 110000 52488
rect 109200 49784 110000 49904
rect 109200 47200 110000 47320
rect 109200 44616 110000 44736
rect 109200 42032 110000 42152
rect 109200 39448 110000 39568
rect 109200 36864 110000 36984
rect 109200 34280 110000 34400
rect 109200 31696 110000 31816
rect 109200 29112 110000 29232
rect 109200 26528 110000 26648
rect 109200 23944 110000 24064
rect 109200 21360 110000 21480
rect 109200 18776 110000 18896
rect 109200 16192 110000 16312
rect 109200 13608 110000 13728
rect 109200 11024 110000 11144
rect 109200 8440 110000 8560
rect 109200 5856 110000 5976
rect 109200 3272 110000 3392
<< obsm3 >>
rect 2957 106832 109200 107745
rect 2957 106552 109120 106832
rect 2957 104248 109200 106552
rect 2957 103968 109120 104248
rect 2957 101664 109200 103968
rect 2957 101384 109120 101664
rect 2957 99080 109200 101384
rect 2957 98800 109120 99080
rect 2957 96496 109200 98800
rect 2957 96216 109120 96496
rect 2957 93912 109200 96216
rect 2957 93632 109120 93912
rect 2957 91328 109200 93632
rect 2957 91048 109120 91328
rect 2957 88744 109200 91048
rect 2957 88464 109120 88744
rect 2957 86160 109200 88464
rect 2957 85880 109120 86160
rect 2957 83576 109200 85880
rect 2957 83296 109120 83576
rect 2957 80992 109200 83296
rect 2957 80712 109120 80992
rect 2957 78408 109200 80712
rect 2957 78128 109120 78408
rect 2957 75824 109200 78128
rect 2957 75544 109120 75824
rect 2957 73240 109200 75544
rect 2957 72960 109120 73240
rect 2957 70656 109200 72960
rect 2957 70376 109120 70656
rect 2957 68072 109200 70376
rect 2957 67792 109120 68072
rect 2957 65488 109200 67792
rect 2957 65208 109120 65488
rect 2957 62904 109200 65208
rect 2957 62624 109120 62904
rect 2957 60320 109200 62624
rect 2957 60040 109120 60320
rect 2957 57736 109200 60040
rect 2957 57456 109120 57736
rect 2957 55152 109200 57456
rect 2957 54872 109120 55152
rect 2957 52568 109200 54872
rect 2957 52288 109120 52568
rect 2957 49984 109200 52288
rect 2957 49704 109120 49984
rect 2957 47400 109200 49704
rect 2957 47120 109120 47400
rect 2957 44816 109200 47120
rect 2957 44536 109120 44816
rect 2957 42232 109200 44536
rect 2957 41952 109120 42232
rect 2957 39648 109200 41952
rect 2957 39368 109120 39648
rect 2957 37064 109200 39368
rect 2957 36784 109120 37064
rect 2957 34480 109200 36784
rect 2957 34200 109120 34480
rect 2957 31896 109200 34200
rect 2957 31616 109120 31896
rect 2957 29312 109200 31616
rect 2957 29032 109120 29312
rect 2957 26728 109200 29032
rect 2957 26448 109120 26728
rect 2957 24144 109200 26448
rect 2957 23864 109120 24144
rect 2957 21560 109200 23864
rect 2957 21280 109120 21560
rect 2957 18976 109200 21280
rect 2957 18696 109120 18976
rect 2957 16392 109200 18696
rect 2957 16112 109120 16392
rect 2957 13808 109200 16112
rect 2957 13528 109120 13808
rect 2957 11224 109200 13528
rect 2957 10944 109120 11224
rect 2957 8640 109200 10944
rect 2957 8360 109120 8640
rect 2957 6056 109200 8360
rect 2957 5776 109120 6056
rect 2957 3472 109200 5776
rect 2957 3192 109120 3472
rect 2957 2143 109200 3192
<< metal4 >>
rect 4208 2128 4528 107760
rect 19568 2128 19888 107760
rect 34928 2128 35248 107760
rect 50288 2128 50608 107760
rect 65648 2128 65968 107760
rect 81008 2128 81328 107760
rect 96368 2128 96688 107760
<< obsm4 >>
rect 13491 2619 19488 106997
rect 19968 2619 34848 106997
rect 35328 2619 50208 106997
rect 50688 2619 65568 106997
rect 66048 2619 80928 106997
rect 81408 2619 96288 106997
rect 96768 2619 107581 106997
<< labels >>
rlabel metal3 s 109200 8440 110000 8560 6 i_addr[0]
port 1 nsew signal input
rlabel metal3 s 109200 16192 110000 16312 6 i_addr[1]
port 2 nsew signal input
rlabel metal3 s 109200 23944 110000 24064 6 i_addr[2]
port 3 nsew signal input
rlabel metal3 s 109200 31696 110000 31816 6 i_addr[3]
port 4 nsew signal input
rlabel metal3 s 109200 39448 110000 39568 6 i_addr[4]
port 5 nsew signal input
rlabel metal3 s 109200 47200 110000 47320 6 i_addr[5]
port 6 nsew signal input
rlabel metal3 s 109200 54952 110000 55072 6 i_addr[6]
port 7 nsew signal input
rlabel metal3 s 109200 3272 110000 3392 6 i_clk
port 8 nsew signal input
rlabel metal3 s 109200 11024 110000 11144 6 i_data[0]
port 9 nsew signal input
rlabel metal3 s 109200 78208 110000 78328 6 i_data[10]
port 10 nsew signal input
rlabel metal3 s 109200 83376 110000 83496 6 i_data[11]
port 11 nsew signal input
rlabel metal3 s 109200 88544 110000 88664 6 i_data[12]
port 12 nsew signal input
rlabel metal3 s 109200 93712 110000 93832 6 i_data[13]
port 13 nsew signal input
rlabel metal3 s 109200 98880 110000 99000 6 i_data[14]
port 14 nsew signal input
rlabel metal3 s 109200 104048 110000 104168 6 i_data[15]
port 15 nsew signal input
rlabel metal3 s 109200 18776 110000 18896 6 i_data[1]
port 16 nsew signal input
rlabel metal3 s 109200 26528 110000 26648 6 i_data[2]
port 17 nsew signal input
rlabel metal3 s 109200 34280 110000 34400 6 i_data[3]
port 18 nsew signal input
rlabel metal3 s 109200 42032 110000 42152 6 i_data[4]
port 19 nsew signal input
rlabel metal3 s 109200 49784 110000 49904 6 i_data[5]
port 20 nsew signal input
rlabel metal3 s 109200 57536 110000 57656 6 i_data[6]
port 21 nsew signal input
rlabel metal3 s 109200 62704 110000 62824 6 i_data[7]
port 22 nsew signal input
rlabel metal3 s 109200 67872 110000 67992 6 i_data[8]
port 23 nsew signal input
rlabel metal3 s 109200 73040 110000 73160 6 i_data[9]
port 24 nsew signal input
rlabel metal3 s 109200 5856 110000 5976 6 i_we
port 25 nsew signal input
rlabel metal3 s 109200 13608 110000 13728 6 o_data[0]
port 26 nsew signal output
rlabel metal3 s 109200 80792 110000 80912 6 o_data[10]
port 27 nsew signal output
rlabel metal3 s 109200 85960 110000 86080 6 o_data[11]
port 28 nsew signal output
rlabel metal3 s 109200 91128 110000 91248 6 o_data[12]
port 29 nsew signal output
rlabel metal3 s 109200 96296 110000 96416 6 o_data[13]
port 30 nsew signal output
rlabel metal3 s 109200 101464 110000 101584 6 o_data[14]
port 31 nsew signal output
rlabel metal3 s 109200 106632 110000 106752 6 o_data[15]
port 32 nsew signal output
rlabel metal3 s 109200 21360 110000 21480 6 o_data[1]
port 33 nsew signal output
rlabel metal3 s 109200 29112 110000 29232 6 o_data[2]
port 34 nsew signal output
rlabel metal3 s 109200 36864 110000 36984 6 o_data[3]
port 35 nsew signal output
rlabel metal3 s 109200 44616 110000 44736 6 o_data[4]
port 36 nsew signal output
rlabel metal3 s 109200 52368 110000 52488 6 o_data[5]
port 37 nsew signal output
rlabel metal3 s 109200 60120 110000 60240 6 o_data[6]
port 38 nsew signal output
rlabel metal3 s 109200 65288 110000 65408 6 o_data[7]
port 39 nsew signal output
rlabel metal3 s 109200 70456 110000 70576 6 o_data[8]
port 40 nsew signal output
rlabel metal3 s 109200 75624 110000 75744 6 o_data[9]
port 41 nsew signal output
rlabel metal4 s 4208 2128 4528 107760 6 vccd1
port 42 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 107760 6 vccd1
port 42 nsew power bidirectional
rlabel metal4 s 65648 2128 65968 107760 6 vccd1
port 42 nsew power bidirectional
rlabel metal4 s 96368 2128 96688 107760 6 vccd1
port 42 nsew power bidirectional
rlabel metal4 s 19568 2128 19888 107760 6 vssd1
port 43 nsew ground bidirectional
rlabel metal4 s 50288 2128 50608 107760 6 vssd1
port 43 nsew ground bidirectional
rlabel metal4 s 81008 2128 81328 107760 6 vssd1
port 43 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 110000 110000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 35221728
string GDS_FILE /home/piotro/caravel_user_project/openlane/int_ram/runs/22_12_31_01_20/results/signoff/int_ram.magic.gds
string GDS_START 493984
<< end >>

