VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO wb_cross_clk
  CLASS BLOCK ;
  FOREIGN wb_cross_clk ;
  ORIGIN 0.000 0.000 ;
  SIZE 200.000 BY 200.000 ;
  PIN clk_m
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 190.990 0.000 191.270 4.000 ;
    END
  END clk_m
  PIN clk_s
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 190.990 196.000 191.270 200.000 ;
    END
  END clk_s
  PIN m_rst
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 8.830 0.000 9.110 4.000 ;
    END
  END m_rst
  PIN m_wb_4_burst
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 11.590 0.000 11.870 4.000 ;
    END
  END m_wb_4_burst
  PIN m_wb_8_burst
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 14.350 0.000 14.630 4.000 ;
    END
  END m_wb_8_burst
  PIN m_wb_ack
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 17.110 0.000 17.390 4.000 ;
    END
  END m_wb_ack
  PIN m_wb_adr[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 19.870 0.000 20.150 4.000 ;
    END
  END m_wb_adr[0]
  PIN m_wb_adr[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 47.470 0.000 47.750 4.000 ;
    END
  END m_wb_adr[10]
  PIN m_wb_adr[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 50.230 0.000 50.510 4.000 ;
    END
  END m_wb_adr[11]
  PIN m_wb_adr[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 52.990 0.000 53.270 4.000 ;
    END
  END m_wb_adr[12]
  PIN m_wb_adr[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 55.750 0.000 56.030 4.000 ;
    END
  END m_wb_adr[13]
  PIN m_wb_adr[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 58.510 0.000 58.790 4.000 ;
    END
  END m_wb_adr[14]
  PIN m_wb_adr[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 61.270 0.000 61.550 4.000 ;
    END
  END m_wb_adr[15]
  PIN m_wb_adr[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 64.030 0.000 64.310 4.000 ;
    END
  END m_wb_adr[16]
  PIN m_wb_adr[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 66.790 0.000 67.070 4.000 ;
    END
  END m_wb_adr[17]
  PIN m_wb_adr[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 69.550 0.000 69.830 4.000 ;
    END
  END m_wb_adr[18]
  PIN m_wb_adr[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 72.310 0.000 72.590 4.000 ;
    END
  END m_wb_adr[19]
  PIN m_wb_adr[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 22.630 0.000 22.910 4.000 ;
    END
  END m_wb_adr[1]
  PIN m_wb_adr[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 75.070 0.000 75.350 4.000 ;
    END
  END m_wb_adr[20]
  PIN m_wb_adr[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 77.830 0.000 78.110 4.000 ;
    END
  END m_wb_adr[21]
  PIN m_wb_adr[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 80.590 0.000 80.870 4.000 ;
    END
  END m_wb_adr[22]
  PIN m_wb_adr[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 83.350 0.000 83.630 4.000 ;
    END
  END m_wb_adr[23]
  PIN m_wb_adr[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 25.390 0.000 25.670 4.000 ;
    END
  END m_wb_adr[2]
  PIN m_wb_adr[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 28.150 0.000 28.430 4.000 ;
    END
  END m_wb_adr[3]
  PIN m_wb_adr[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 30.910 0.000 31.190 4.000 ;
    END
  END m_wb_adr[4]
  PIN m_wb_adr[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 33.670 0.000 33.950 4.000 ;
    END
  END m_wb_adr[5]
  PIN m_wb_adr[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 36.430 0.000 36.710 4.000 ;
    END
  END m_wb_adr[6]
  PIN m_wb_adr[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 39.190 0.000 39.470 4.000 ;
    END
  END m_wb_adr[7]
  PIN m_wb_adr[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 41.950 0.000 42.230 4.000 ;
    END
  END m_wb_adr[8]
  PIN m_wb_adr[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 44.710 0.000 44.990 4.000 ;
    END
  END m_wb_adr[9]
  PIN m_wb_cyc
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 86.110 0.000 86.390 4.000 ;
    END
  END m_wb_cyc
  PIN m_wb_err
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 88.870 0.000 89.150 4.000 ;
    END
  END m_wb_err
  PIN m_wb_i_dat[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 91.630 0.000 91.910 4.000 ;
    END
  END m_wb_i_dat[0]
  PIN m_wb_i_dat[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 119.230 0.000 119.510 4.000 ;
    END
  END m_wb_i_dat[10]
  PIN m_wb_i_dat[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 121.990 0.000 122.270 4.000 ;
    END
  END m_wb_i_dat[11]
  PIN m_wb_i_dat[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 124.750 0.000 125.030 4.000 ;
    END
  END m_wb_i_dat[12]
  PIN m_wb_i_dat[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 127.510 0.000 127.790 4.000 ;
    END
  END m_wb_i_dat[13]
  PIN m_wb_i_dat[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 130.270 0.000 130.550 4.000 ;
    END
  END m_wb_i_dat[14]
  PIN m_wb_i_dat[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 133.030 0.000 133.310 4.000 ;
    END
  END m_wb_i_dat[15]
  PIN m_wb_i_dat[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 94.390 0.000 94.670 4.000 ;
    END
  END m_wb_i_dat[1]
  PIN m_wb_i_dat[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 97.150 0.000 97.430 4.000 ;
    END
  END m_wb_i_dat[2]
  PIN m_wb_i_dat[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 99.910 0.000 100.190 4.000 ;
    END
  END m_wb_i_dat[3]
  PIN m_wb_i_dat[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 102.670 0.000 102.950 4.000 ;
    END
  END m_wb_i_dat[4]
  PIN m_wb_i_dat[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 105.430 0.000 105.710 4.000 ;
    END
  END m_wb_i_dat[5]
  PIN m_wb_i_dat[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 108.190 0.000 108.470 4.000 ;
    END
  END m_wb_i_dat[6]
  PIN m_wb_i_dat[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 110.950 0.000 111.230 4.000 ;
    END
  END m_wb_i_dat[7]
  PIN m_wb_i_dat[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 113.710 0.000 113.990 4.000 ;
    END
  END m_wb_i_dat[8]
  PIN m_wb_i_dat[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 116.470 0.000 116.750 4.000 ;
    END
  END m_wb_i_dat[9]
  PIN m_wb_o_dat[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 135.790 0.000 136.070 4.000 ;
    END
  END m_wb_o_dat[0]
  PIN m_wb_o_dat[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 163.390 0.000 163.670 4.000 ;
    END
  END m_wb_o_dat[10]
  PIN m_wb_o_dat[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 166.150 0.000 166.430 4.000 ;
    END
  END m_wb_o_dat[11]
  PIN m_wb_o_dat[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 168.910 0.000 169.190 4.000 ;
    END
  END m_wb_o_dat[12]
  PIN m_wb_o_dat[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 171.670 0.000 171.950 4.000 ;
    END
  END m_wb_o_dat[13]
  PIN m_wb_o_dat[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 174.430 0.000 174.710 4.000 ;
    END
  END m_wb_o_dat[14]
  PIN m_wb_o_dat[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 177.190 0.000 177.470 4.000 ;
    END
  END m_wb_o_dat[15]
  PIN m_wb_o_dat[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 138.550 0.000 138.830 4.000 ;
    END
  END m_wb_o_dat[1]
  PIN m_wb_o_dat[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 141.310 0.000 141.590 4.000 ;
    END
  END m_wb_o_dat[2]
  PIN m_wb_o_dat[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 144.070 0.000 144.350 4.000 ;
    END
  END m_wb_o_dat[3]
  PIN m_wb_o_dat[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 146.830 0.000 147.110 4.000 ;
    END
  END m_wb_o_dat[4]
  PIN m_wb_o_dat[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 149.590 0.000 149.870 4.000 ;
    END
  END m_wb_o_dat[5]
  PIN m_wb_o_dat[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 152.350 0.000 152.630 4.000 ;
    END
  END m_wb_o_dat[6]
  PIN m_wb_o_dat[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 155.110 0.000 155.390 4.000 ;
    END
  END m_wb_o_dat[7]
  PIN m_wb_o_dat[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 157.870 0.000 158.150 4.000 ;
    END
  END m_wb_o_dat[8]
  PIN m_wb_o_dat[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 160.630 0.000 160.910 4.000 ;
    END
  END m_wb_o_dat[9]
  PIN m_wb_sel[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 179.950 0.000 180.230 4.000 ;
    END
  END m_wb_sel[0]
  PIN m_wb_sel[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 182.710 0.000 182.990 4.000 ;
    END
  END m_wb_sel[1]
  PIN m_wb_stb
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 185.470 0.000 185.750 4.000 ;
    END
  END m_wb_stb
  PIN m_wb_we
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 188.230 0.000 188.510 4.000 ;
    END
  END m_wb_we
  PIN s_rst
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 8.830 196.000 9.110 200.000 ;
    END
  END s_rst
  PIN s_wb_4_burst
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 11.590 196.000 11.870 200.000 ;
    END
  END s_wb_4_burst
  PIN s_wb_8_burst
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 14.350 196.000 14.630 200.000 ;
    END
  END s_wb_8_burst
  PIN s_wb_ack
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 17.110 196.000 17.390 200.000 ;
    END
  END s_wb_ack
  PIN s_wb_adr[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 19.870 196.000 20.150 200.000 ;
    END
  END s_wb_adr[0]
  PIN s_wb_adr[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 47.470 196.000 47.750 200.000 ;
    END
  END s_wb_adr[10]
  PIN s_wb_adr[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 50.230 196.000 50.510 200.000 ;
    END
  END s_wb_adr[11]
  PIN s_wb_adr[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 52.990 196.000 53.270 200.000 ;
    END
  END s_wb_adr[12]
  PIN s_wb_adr[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 55.750 196.000 56.030 200.000 ;
    END
  END s_wb_adr[13]
  PIN s_wb_adr[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 58.510 196.000 58.790 200.000 ;
    END
  END s_wb_adr[14]
  PIN s_wb_adr[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 61.270 196.000 61.550 200.000 ;
    END
  END s_wb_adr[15]
  PIN s_wb_adr[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 64.030 196.000 64.310 200.000 ;
    END
  END s_wb_adr[16]
  PIN s_wb_adr[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 66.790 196.000 67.070 200.000 ;
    END
  END s_wb_adr[17]
  PIN s_wb_adr[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 69.550 196.000 69.830 200.000 ;
    END
  END s_wb_adr[18]
  PIN s_wb_adr[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 72.310 196.000 72.590 200.000 ;
    END
  END s_wb_adr[19]
  PIN s_wb_adr[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 22.630 196.000 22.910 200.000 ;
    END
  END s_wb_adr[1]
  PIN s_wb_adr[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 75.070 196.000 75.350 200.000 ;
    END
  END s_wb_adr[20]
  PIN s_wb_adr[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 77.830 196.000 78.110 200.000 ;
    END
  END s_wb_adr[21]
  PIN s_wb_adr[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 80.590 196.000 80.870 200.000 ;
    END
  END s_wb_adr[22]
  PIN s_wb_adr[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 83.350 196.000 83.630 200.000 ;
    END
  END s_wb_adr[23]
  PIN s_wb_adr[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 25.390 196.000 25.670 200.000 ;
    END
  END s_wb_adr[2]
  PIN s_wb_adr[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 28.150 196.000 28.430 200.000 ;
    END
  END s_wb_adr[3]
  PIN s_wb_adr[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 30.910 196.000 31.190 200.000 ;
    END
  END s_wb_adr[4]
  PIN s_wb_adr[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 33.670 196.000 33.950 200.000 ;
    END
  END s_wb_adr[5]
  PIN s_wb_adr[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 36.430 196.000 36.710 200.000 ;
    END
  END s_wb_adr[6]
  PIN s_wb_adr[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 39.190 196.000 39.470 200.000 ;
    END
  END s_wb_adr[7]
  PIN s_wb_adr[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 41.950 196.000 42.230 200.000 ;
    END
  END s_wb_adr[8]
  PIN s_wb_adr[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 44.710 196.000 44.990 200.000 ;
    END
  END s_wb_adr[9]
  PIN s_wb_cyc
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 86.110 196.000 86.390 200.000 ;
    END
  END s_wb_cyc
  PIN s_wb_err
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 88.870 196.000 89.150 200.000 ;
    END
  END s_wb_err
  PIN s_wb_i_dat[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 91.630 196.000 91.910 200.000 ;
    END
  END s_wb_i_dat[0]
  PIN s_wb_i_dat[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 119.230 196.000 119.510 200.000 ;
    END
  END s_wb_i_dat[10]
  PIN s_wb_i_dat[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 121.990 196.000 122.270 200.000 ;
    END
  END s_wb_i_dat[11]
  PIN s_wb_i_dat[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 124.750 196.000 125.030 200.000 ;
    END
  END s_wb_i_dat[12]
  PIN s_wb_i_dat[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 127.510 196.000 127.790 200.000 ;
    END
  END s_wb_i_dat[13]
  PIN s_wb_i_dat[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 130.270 196.000 130.550 200.000 ;
    END
  END s_wb_i_dat[14]
  PIN s_wb_i_dat[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 133.030 196.000 133.310 200.000 ;
    END
  END s_wb_i_dat[15]
  PIN s_wb_i_dat[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 94.390 196.000 94.670 200.000 ;
    END
  END s_wb_i_dat[1]
  PIN s_wb_i_dat[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 97.150 196.000 97.430 200.000 ;
    END
  END s_wb_i_dat[2]
  PIN s_wb_i_dat[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 99.910 196.000 100.190 200.000 ;
    END
  END s_wb_i_dat[3]
  PIN s_wb_i_dat[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 102.670 196.000 102.950 200.000 ;
    END
  END s_wb_i_dat[4]
  PIN s_wb_i_dat[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 105.430 196.000 105.710 200.000 ;
    END
  END s_wb_i_dat[5]
  PIN s_wb_i_dat[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 108.190 196.000 108.470 200.000 ;
    END
  END s_wb_i_dat[6]
  PIN s_wb_i_dat[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 110.950 196.000 111.230 200.000 ;
    END
  END s_wb_i_dat[7]
  PIN s_wb_i_dat[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 113.710 196.000 113.990 200.000 ;
    END
  END s_wb_i_dat[8]
  PIN s_wb_i_dat[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 116.470 196.000 116.750 200.000 ;
    END
  END s_wb_i_dat[9]
  PIN s_wb_o_dat[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 135.790 196.000 136.070 200.000 ;
    END
  END s_wb_o_dat[0]
  PIN s_wb_o_dat[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 163.390 196.000 163.670 200.000 ;
    END
  END s_wb_o_dat[10]
  PIN s_wb_o_dat[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 166.150 196.000 166.430 200.000 ;
    END
  END s_wb_o_dat[11]
  PIN s_wb_o_dat[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 168.910 196.000 169.190 200.000 ;
    END
  END s_wb_o_dat[12]
  PIN s_wb_o_dat[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 171.670 196.000 171.950 200.000 ;
    END
  END s_wb_o_dat[13]
  PIN s_wb_o_dat[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 174.430 196.000 174.710 200.000 ;
    END
  END s_wb_o_dat[14]
  PIN s_wb_o_dat[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 177.190 196.000 177.470 200.000 ;
    END
  END s_wb_o_dat[15]
  PIN s_wb_o_dat[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 138.550 196.000 138.830 200.000 ;
    END
  END s_wb_o_dat[1]
  PIN s_wb_o_dat[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 141.310 196.000 141.590 200.000 ;
    END
  END s_wb_o_dat[2]
  PIN s_wb_o_dat[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 144.070 196.000 144.350 200.000 ;
    END
  END s_wb_o_dat[3]
  PIN s_wb_o_dat[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 146.830 196.000 147.110 200.000 ;
    END
  END s_wb_o_dat[4]
  PIN s_wb_o_dat[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 149.590 196.000 149.870 200.000 ;
    END
  END s_wb_o_dat[5]
  PIN s_wb_o_dat[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 152.350 196.000 152.630 200.000 ;
    END
  END s_wb_o_dat[6]
  PIN s_wb_o_dat[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 155.110 196.000 155.390 200.000 ;
    END
  END s_wb_o_dat[7]
  PIN s_wb_o_dat[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 157.870 196.000 158.150 200.000 ;
    END
  END s_wb_o_dat[8]
  PIN s_wb_o_dat[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 160.630 196.000 160.910 200.000 ;
    END
  END s_wb_o_dat[9]
  PIN s_wb_sel[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 179.950 196.000 180.230 200.000 ;
    END
  END s_wb_sel[0]
  PIN s_wb_sel[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 182.710 196.000 182.990 200.000 ;
    END
  END s_wb_sel[1]
  PIN s_wb_stb
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 185.470 196.000 185.750 200.000 ;
    END
  END s_wb_stb
  PIN s_wb_we
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 188.230 196.000 188.510 200.000 ;
    END
  END s_wb_we
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 187.920 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 187.920 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 187.920 ;
    END
  END vssd1
  OBS
      LAYER nwell ;
        RECT 5.330 186.265 194.310 187.870 ;
        RECT 5.330 180.825 194.310 183.655 ;
        RECT 5.330 175.385 194.310 178.215 ;
        RECT 5.330 169.945 194.310 172.775 ;
        RECT 5.330 164.505 194.310 167.335 ;
        RECT 5.330 159.065 194.310 161.895 ;
        RECT 5.330 153.625 194.310 156.455 ;
        RECT 5.330 148.185 194.310 151.015 ;
        RECT 5.330 142.745 194.310 145.575 ;
        RECT 5.330 137.305 194.310 140.135 ;
        RECT 5.330 131.865 194.310 134.695 ;
        RECT 5.330 126.425 194.310 129.255 ;
        RECT 5.330 120.985 194.310 123.815 ;
        RECT 5.330 115.545 194.310 118.375 ;
        RECT 5.330 110.105 194.310 112.935 ;
        RECT 5.330 104.665 194.310 107.495 ;
        RECT 5.330 99.225 194.310 102.055 ;
        RECT 5.330 93.785 194.310 96.615 ;
        RECT 5.330 88.345 194.310 91.175 ;
        RECT 5.330 82.905 194.310 85.735 ;
        RECT 5.330 77.465 194.310 80.295 ;
        RECT 5.330 72.025 194.310 74.855 ;
        RECT 5.330 66.585 194.310 69.415 ;
        RECT 5.330 61.145 194.310 63.975 ;
        RECT 5.330 55.705 194.310 58.535 ;
        RECT 5.330 50.265 194.310 53.095 ;
        RECT 5.330 44.825 194.310 47.655 ;
        RECT 5.330 39.385 194.310 42.215 ;
        RECT 5.330 33.945 194.310 36.775 ;
        RECT 5.330 28.505 194.310 31.335 ;
        RECT 5.330 23.065 194.310 25.895 ;
        RECT 5.330 17.625 194.310 20.455 ;
        RECT 5.330 12.185 194.310 15.015 ;
      LAYER li1 ;
        RECT 5.520 10.795 194.120 187.765 ;
      LAYER met1 ;
        RECT 5.520 6.840 194.120 188.660 ;
      LAYER met2 ;
        RECT 9.390 195.720 11.310 196.250 ;
        RECT 12.150 195.720 14.070 196.250 ;
        RECT 14.910 195.720 16.830 196.250 ;
        RECT 17.670 195.720 19.590 196.250 ;
        RECT 20.430 195.720 22.350 196.250 ;
        RECT 23.190 195.720 25.110 196.250 ;
        RECT 25.950 195.720 27.870 196.250 ;
        RECT 28.710 195.720 30.630 196.250 ;
        RECT 31.470 195.720 33.390 196.250 ;
        RECT 34.230 195.720 36.150 196.250 ;
        RECT 36.990 195.720 38.910 196.250 ;
        RECT 39.750 195.720 41.670 196.250 ;
        RECT 42.510 195.720 44.430 196.250 ;
        RECT 45.270 195.720 47.190 196.250 ;
        RECT 48.030 195.720 49.950 196.250 ;
        RECT 50.790 195.720 52.710 196.250 ;
        RECT 53.550 195.720 55.470 196.250 ;
        RECT 56.310 195.720 58.230 196.250 ;
        RECT 59.070 195.720 60.990 196.250 ;
        RECT 61.830 195.720 63.750 196.250 ;
        RECT 64.590 195.720 66.510 196.250 ;
        RECT 67.350 195.720 69.270 196.250 ;
        RECT 70.110 195.720 72.030 196.250 ;
        RECT 72.870 195.720 74.790 196.250 ;
        RECT 75.630 195.720 77.550 196.250 ;
        RECT 78.390 195.720 80.310 196.250 ;
        RECT 81.150 195.720 83.070 196.250 ;
        RECT 83.910 195.720 85.830 196.250 ;
        RECT 86.670 195.720 88.590 196.250 ;
        RECT 89.430 195.720 91.350 196.250 ;
        RECT 92.190 195.720 94.110 196.250 ;
        RECT 94.950 195.720 96.870 196.250 ;
        RECT 97.710 195.720 99.630 196.250 ;
        RECT 100.470 195.720 102.390 196.250 ;
        RECT 103.230 195.720 105.150 196.250 ;
        RECT 105.990 195.720 107.910 196.250 ;
        RECT 108.750 195.720 110.670 196.250 ;
        RECT 111.510 195.720 113.430 196.250 ;
        RECT 114.270 195.720 116.190 196.250 ;
        RECT 117.030 195.720 118.950 196.250 ;
        RECT 119.790 195.720 121.710 196.250 ;
        RECT 122.550 195.720 124.470 196.250 ;
        RECT 125.310 195.720 127.230 196.250 ;
        RECT 128.070 195.720 129.990 196.250 ;
        RECT 130.830 195.720 132.750 196.250 ;
        RECT 133.590 195.720 135.510 196.250 ;
        RECT 136.350 195.720 138.270 196.250 ;
        RECT 139.110 195.720 141.030 196.250 ;
        RECT 141.870 195.720 143.790 196.250 ;
        RECT 144.630 195.720 146.550 196.250 ;
        RECT 147.390 195.720 149.310 196.250 ;
        RECT 150.150 195.720 152.070 196.250 ;
        RECT 152.910 195.720 154.830 196.250 ;
        RECT 155.670 195.720 157.590 196.250 ;
        RECT 158.430 195.720 160.350 196.250 ;
        RECT 161.190 195.720 163.110 196.250 ;
        RECT 163.950 195.720 165.870 196.250 ;
        RECT 166.710 195.720 168.630 196.250 ;
        RECT 169.470 195.720 171.390 196.250 ;
        RECT 172.230 195.720 174.150 196.250 ;
        RECT 174.990 195.720 176.910 196.250 ;
        RECT 177.750 195.720 179.670 196.250 ;
        RECT 180.510 195.720 182.430 196.250 ;
        RECT 183.270 195.720 185.190 196.250 ;
        RECT 186.030 195.720 187.950 196.250 ;
        RECT 188.790 195.720 190.710 196.250 ;
        RECT 191.550 195.720 191.730 196.250 ;
        RECT 8.840 4.280 191.730 195.720 ;
        RECT 9.390 3.670 11.310 4.280 ;
        RECT 12.150 3.670 14.070 4.280 ;
        RECT 14.910 3.670 16.830 4.280 ;
        RECT 17.670 3.670 19.590 4.280 ;
        RECT 20.430 3.670 22.350 4.280 ;
        RECT 23.190 3.670 25.110 4.280 ;
        RECT 25.950 3.670 27.870 4.280 ;
        RECT 28.710 3.670 30.630 4.280 ;
        RECT 31.470 3.670 33.390 4.280 ;
        RECT 34.230 3.670 36.150 4.280 ;
        RECT 36.990 3.670 38.910 4.280 ;
        RECT 39.750 3.670 41.670 4.280 ;
        RECT 42.510 3.670 44.430 4.280 ;
        RECT 45.270 3.670 47.190 4.280 ;
        RECT 48.030 3.670 49.950 4.280 ;
        RECT 50.790 3.670 52.710 4.280 ;
        RECT 53.550 3.670 55.470 4.280 ;
        RECT 56.310 3.670 58.230 4.280 ;
        RECT 59.070 3.670 60.990 4.280 ;
        RECT 61.830 3.670 63.750 4.280 ;
        RECT 64.590 3.670 66.510 4.280 ;
        RECT 67.350 3.670 69.270 4.280 ;
        RECT 70.110 3.670 72.030 4.280 ;
        RECT 72.870 3.670 74.790 4.280 ;
        RECT 75.630 3.670 77.550 4.280 ;
        RECT 78.390 3.670 80.310 4.280 ;
        RECT 81.150 3.670 83.070 4.280 ;
        RECT 83.910 3.670 85.830 4.280 ;
        RECT 86.670 3.670 88.590 4.280 ;
        RECT 89.430 3.670 91.350 4.280 ;
        RECT 92.190 3.670 94.110 4.280 ;
        RECT 94.950 3.670 96.870 4.280 ;
        RECT 97.710 3.670 99.630 4.280 ;
        RECT 100.470 3.670 102.390 4.280 ;
        RECT 103.230 3.670 105.150 4.280 ;
        RECT 105.990 3.670 107.910 4.280 ;
        RECT 108.750 3.670 110.670 4.280 ;
        RECT 111.510 3.670 113.430 4.280 ;
        RECT 114.270 3.670 116.190 4.280 ;
        RECT 117.030 3.670 118.950 4.280 ;
        RECT 119.790 3.670 121.710 4.280 ;
        RECT 122.550 3.670 124.470 4.280 ;
        RECT 125.310 3.670 127.230 4.280 ;
        RECT 128.070 3.670 129.990 4.280 ;
        RECT 130.830 3.670 132.750 4.280 ;
        RECT 133.590 3.670 135.510 4.280 ;
        RECT 136.350 3.670 138.270 4.280 ;
        RECT 139.110 3.670 141.030 4.280 ;
        RECT 141.870 3.670 143.790 4.280 ;
        RECT 144.630 3.670 146.550 4.280 ;
        RECT 147.390 3.670 149.310 4.280 ;
        RECT 150.150 3.670 152.070 4.280 ;
        RECT 152.910 3.670 154.830 4.280 ;
        RECT 155.670 3.670 157.590 4.280 ;
        RECT 158.430 3.670 160.350 4.280 ;
        RECT 161.190 3.670 163.110 4.280 ;
        RECT 163.950 3.670 165.870 4.280 ;
        RECT 166.710 3.670 168.630 4.280 ;
        RECT 169.470 3.670 171.390 4.280 ;
        RECT 172.230 3.670 174.150 4.280 ;
        RECT 174.990 3.670 176.910 4.280 ;
        RECT 177.750 3.670 179.670 4.280 ;
        RECT 180.510 3.670 182.430 4.280 ;
        RECT 183.270 3.670 185.190 4.280 ;
        RECT 186.030 3.670 187.950 4.280 ;
        RECT 188.790 3.670 190.710 4.280 ;
        RECT 191.550 3.670 191.730 4.280 ;
      LAYER met3 ;
        RECT 21.050 8.335 191.755 187.845 ;
      LAYER met4 ;
        RECT 93.215 10.240 97.440 182.745 ;
        RECT 99.840 10.240 174.240 182.745 ;
        RECT 176.640 10.240 182.785 182.745 ;
        RECT 93.215 8.335 182.785 10.240 ;
  END
END wb_cross_clk
END LIBRARY

