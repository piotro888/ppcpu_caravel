magic
tech sky130B
magscale 1 2
timestamp 1663070636
<< obsli1 >>
rect 1104 2159 38824 37553
<< obsm1 >>
rect 14 2128 39362 37584
<< metal2 >>
rect 18 39200 74 40000
rect 662 39200 718 40000
rect 1950 39200 2006 40000
rect 2594 39200 2650 40000
rect 3238 39200 3294 40000
rect 4526 39200 4582 40000
rect 5170 39200 5226 40000
rect 5814 39200 5870 40000
rect 7102 39200 7158 40000
rect 7746 39200 7802 40000
rect 8390 39200 8446 40000
rect 9678 39200 9734 40000
rect 10322 39200 10378 40000
rect 10966 39200 11022 40000
rect 12254 39200 12310 40000
rect 12898 39200 12954 40000
rect 13542 39200 13598 40000
rect 14186 39200 14242 40000
rect 15474 39200 15530 40000
rect 16118 39200 16174 40000
rect 16762 39200 16818 40000
rect 18050 39200 18106 40000
rect 18694 39200 18750 40000
rect 19338 39200 19394 40000
rect 20626 39200 20682 40000
rect 21270 39200 21326 40000
rect 21914 39200 21970 40000
rect 23202 39200 23258 40000
rect 23846 39200 23902 40000
rect 24490 39200 24546 40000
rect 25778 39200 25834 40000
rect 26422 39200 26478 40000
rect 27066 39200 27122 40000
rect 28354 39200 28410 40000
rect 28998 39200 29054 40000
rect 29642 39200 29698 40000
rect 30930 39200 30986 40000
rect 31574 39200 31630 40000
rect 32218 39200 32274 40000
rect 33506 39200 33562 40000
rect 34150 39200 34206 40000
rect 34794 39200 34850 40000
rect 36082 39200 36138 40000
rect 36726 39200 36782 40000
rect 37370 39200 37426 40000
rect 38658 39200 38714 40000
rect 39302 39200 39358 40000
rect 18 0 74 800
rect 662 0 718 800
rect 1306 0 1362 800
rect 1950 0 2006 800
rect 3238 0 3294 800
rect 3882 0 3938 800
rect 4526 0 4582 800
rect 5814 0 5870 800
rect 6458 0 6514 800
rect 7102 0 7158 800
rect 8390 0 8446 800
rect 9034 0 9090 800
rect 9678 0 9734 800
rect 10966 0 11022 800
rect 11610 0 11666 800
rect 12254 0 12310 800
rect 13542 0 13598 800
rect 14186 0 14242 800
rect 14830 0 14886 800
rect 16118 0 16174 800
rect 16762 0 16818 800
rect 17406 0 17462 800
rect 18694 0 18750 800
rect 19338 0 19394 800
rect 19982 0 20038 800
rect 21270 0 21326 800
rect 21914 0 21970 800
rect 22558 0 22614 800
rect 23846 0 23902 800
rect 24490 0 24546 800
rect 25134 0 25190 800
rect 25778 0 25834 800
rect 27066 0 27122 800
rect 27710 0 27766 800
rect 28354 0 28410 800
rect 29642 0 29698 800
rect 30286 0 30342 800
rect 30930 0 30986 800
rect 32218 0 32274 800
rect 32862 0 32918 800
rect 33506 0 33562 800
rect 34794 0 34850 800
rect 35438 0 35494 800
rect 36082 0 36138 800
rect 37370 0 37426 800
rect 38014 0 38070 800
rect 38658 0 38714 800
<< obsm2 >>
rect 130 39144 606 39545
rect 774 39144 1894 39545
rect 2062 39144 2538 39545
rect 2706 39144 3182 39545
rect 3350 39144 4470 39545
rect 4638 39144 5114 39545
rect 5282 39144 5758 39545
rect 5926 39144 7046 39545
rect 7214 39144 7690 39545
rect 7858 39144 8334 39545
rect 8502 39144 9622 39545
rect 9790 39144 10266 39545
rect 10434 39144 10910 39545
rect 11078 39144 12198 39545
rect 12366 39144 12842 39545
rect 13010 39144 13486 39545
rect 13654 39144 14130 39545
rect 14298 39144 15418 39545
rect 15586 39144 16062 39545
rect 16230 39144 16706 39545
rect 16874 39144 17994 39545
rect 18162 39144 18638 39545
rect 18806 39144 19282 39545
rect 19450 39144 20570 39545
rect 20738 39144 21214 39545
rect 21382 39144 21858 39545
rect 22026 39144 23146 39545
rect 23314 39144 23790 39545
rect 23958 39144 24434 39545
rect 24602 39144 25722 39545
rect 25890 39144 26366 39545
rect 26534 39144 27010 39545
rect 27178 39144 28298 39545
rect 28466 39144 28942 39545
rect 29110 39144 29586 39545
rect 29754 39144 30874 39545
rect 31042 39144 31518 39545
rect 31686 39144 32162 39545
rect 32330 39144 33450 39545
rect 33618 39144 34094 39545
rect 34262 39144 34738 39545
rect 34906 39144 36026 39545
rect 36194 39144 36670 39545
rect 36838 39144 37314 39545
rect 37482 39144 38602 39545
rect 38770 39144 39246 39545
rect 20 856 39356 39144
rect 130 31 606 856
rect 774 31 1250 856
rect 1418 31 1894 856
rect 2062 31 3182 856
rect 3350 31 3826 856
rect 3994 31 4470 856
rect 4638 31 5758 856
rect 5926 31 6402 856
rect 6570 31 7046 856
rect 7214 31 8334 856
rect 8502 31 8978 856
rect 9146 31 9622 856
rect 9790 31 10910 856
rect 11078 31 11554 856
rect 11722 31 12198 856
rect 12366 31 13486 856
rect 13654 31 14130 856
rect 14298 31 14774 856
rect 14942 31 16062 856
rect 16230 31 16706 856
rect 16874 31 17350 856
rect 17518 31 18638 856
rect 18806 31 19282 856
rect 19450 31 19926 856
rect 20094 31 21214 856
rect 21382 31 21858 856
rect 22026 31 22502 856
rect 22670 31 23790 856
rect 23958 31 24434 856
rect 24602 31 25078 856
rect 25246 31 25722 856
rect 25890 31 27010 856
rect 27178 31 27654 856
rect 27822 31 28298 856
rect 28466 31 29586 856
rect 29754 31 30230 856
rect 30398 31 30874 856
rect 31042 31 32162 856
rect 32330 31 32806 856
rect 32974 31 33450 856
rect 33618 31 34738 856
rect 34906 31 35382 856
rect 35550 31 36026 856
rect 36194 31 37314 856
rect 37482 31 37958 856
rect 38126 31 38602 856
rect 38770 31 39356 856
<< metal3 >>
rect 0 39448 800 39568
rect 39200 39448 40000 39568
rect 39200 38768 40000 38888
rect 0 38088 800 38208
rect 0 37408 800 37528
rect 39200 37408 40000 37528
rect 0 36728 800 36848
rect 39200 36728 40000 36848
rect 39200 36048 40000 36168
rect 0 35368 800 35488
rect 0 34688 800 34808
rect 39200 34688 40000 34808
rect 0 34008 800 34128
rect 39200 34008 40000 34128
rect 39200 33328 40000 33448
rect 0 32648 800 32768
rect 0 31968 800 32088
rect 39200 31968 40000 32088
rect 0 31288 800 31408
rect 39200 31288 40000 31408
rect 39200 30608 40000 30728
rect 0 29928 800 30048
rect 0 29248 800 29368
rect 39200 29248 40000 29368
rect 0 28568 800 28688
rect 39200 28568 40000 28688
rect 39200 27888 40000 28008
rect 0 27208 800 27328
rect 0 26528 800 26648
rect 39200 26528 40000 26648
rect 0 25848 800 25968
rect 39200 25848 40000 25968
rect 0 25168 800 25288
rect 39200 25168 40000 25288
rect 0 23808 800 23928
rect 39200 23808 40000 23928
rect 0 23128 800 23248
rect 39200 23128 40000 23248
rect 0 22448 800 22568
rect 39200 22448 40000 22568
rect 0 21088 800 21208
rect 39200 21088 40000 21208
rect 0 20408 800 20528
rect 39200 20408 40000 20528
rect 0 19728 800 19848
rect 39200 19728 40000 19848
rect 0 18368 800 18488
rect 39200 18368 40000 18488
rect 0 17688 800 17808
rect 39200 17688 40000 17808
rect 0 17008 800 17128
rect 39200 17008 40000 17128
rect 0 15648 800 15768
rect 39200 15648 40000 15768
rect 0 14968 800 15088
rect 39200 14968 40000 15088
rect 0 14288 800 14408
rect 39200 14288 40000 14408
rect 0 12928 800 13048
rect 39200 12928 40000 13048
rect 0 12248 800 12368
rect 39200 12248 40000 12368
rect 0 11568 800 11688
rect 39200 11568 40000 11688
rect 39200 10888 40000 11008
rect 0 10208 800 10328
rect 0 9528 800 9648
rect 39200 9528 40000 9648
rect 0 8848 800 8968
rect 39200 8848 40000 8968
rect 39200 8168 40000 8288
rect 0 7488 800 7608
rect 0 6808 800 6928
rect 39200 6808 40000 6928
rect 0 6128 800 6248
rect 39200 6128 40000 6248
rect 39200 5448 40000 5568
rect 0 4768 800 4888
rect 0 4088 800 4208
rect 39200 4088 40000 4208
rect 0 3408 800 3528
rect 39200 3408 40000 3528
rect 39200 2728 40000 2848
rect 0 2048 800 2168
rect 0 1368 800 1488
rect 39200 1368 40000 1488
rect 0 688 800 808
rect 39200 688 40000 808
rect 39200 8 40000 128
<< obsm3 >>
rect 880 39368 39120 39541
rect 800 38968 39200 39368
rect 800 38688 39120 38968
rect 800 38288 39200 38688
rect 880 38008 39200 38288
rect 800 37608 39200 38008
rect 880 37328 39120 37608
rect 800 36928 39200 37328
rect 880 36648 39120 36928
rect 800 36248 39200 36648
rect 800 35968 39120 36248
rect 800 35568 39200 35968
rect 880 35288 39200 35568
rect 800 34888 39200 35288
rect 880 34608 39120 34888
rect 800 34208 39200 34608
rect 880 33928 39120 34208
rect 800 33528 39200 33928
rect 800 33248 39120 33528
rect 800 32848 39200 33248
rect 880 32568 39200 32848
rect 800 32168 39200 32568
rect 880 31888 39120 32168
rect 800 31488 39200 31888
rect 880 31208 39120 31488
rect 800 30808 39200 31208
rect 800 30528 39120 30808
rect 800 30128 39200 30528
rect 880 29848 39200 30128
rect 800 29448 39200 29848
rect 880 29168 39120 29448
rect 800 28768 39200 29168
rect 880 28488 39120 28768
rect 800 28088 39200 28488
rect 800 27808 39120 28088
rect 800 27408 39200 27808
rect 880 27128 39200 27408
rect 800 26728 39200 27128
rect 880 26448 39120 26728
rect 800 26048 39200 26448
rect 880 25768 39120 26048
rect 800 25368 39200 25768
rect 880 25088 39120 25368
rect 800 24008 39200 25088
rect 880 23728 39120 24008
rect 800 23328 39200 23728
rect 880 23048 39120 23328
rect 800 22648 39200 23048
rect 880 22368 39120 22648
rect 800 21288 39200 22368
rect 880 21008 39120 21288
rect 800 20608 39200 21008
rect 880 20328 39120 20608
rect 800 19928 39200 20328
rect 880 19648 39120 19928
rect 800 18568 39200 19648
rect 880 18288 39120 18568
rect 800 17888 39200 18288
rect 880 17608 39120 17888
rect 800 17208 39200 17608
rect 880 16928 39120 17208
rect 800 15848 39200 16928
rect 880 15568 39120 15848
rect 800 15168 39200 15568
rect 880 14888 39120 15168
rect 800 14488 39200 14888
rect 880 14208 39120 14488
rect 800 13128 39200 14208
rect 880 12848 39120 13128
rect 800 12448 39200 12848
rect 880 12168 39120 12448
rect 800 11768 39200 12168
rect 880 11488 39120 11768
rect 800 11088 39200 11488
rect 800 10808 39120 11088
rect 800 10408 39200 10808
rect 880 10128 39200 10408
rect 800 9728 39200 10128
rect 880 9448 39120 9728
rect 800 9048 39200 9448
rect 880 8768 39120 9048
rect 800 8368 39200 8768
rect 800 8088 39120 8368
rect 800 7688 39200 8088
rect 880 7408 39200 7688
rect 800 7008 39200 7408
rect 880 6728 39120 7008
rect 800 6328 39200 6728
rect 880 6048 39120 6328
rect 800 5648 39200 6048
rect 800 5368 39120 5648
rect 800 4968 39200 5368
rect 880 4688 39200 4968
rect 800 4288 39200 4688
rect 880 4008 39120 4288
rect 800 3608 39200 4008
rect 880 3328 39120 3608
rect 800 2928 39200 3328
rect 800 2648 39120 2928
rect 800 2248 39200 2648
rect 880 1968 39200 2248
rect 800 1568 39200 1968
rect 880 1288 39120 1568
rect 800 888 39200 1288
rect 880 608 39120 888
rect 800 208 39200 608
rect 800 35 39120 208
<< metal4 >>
rect 4208 2128 4528 37584
rect 19568 2128 19888 37584
rect 34928 2128 35248 37584
<< labels >>
rlabel metal2 s 30930 39200 30986 40000 6 b0_drv[0]
port 1 nsew signal output
rlabel metal2 s 25778 39200 25834 40000 6 b0_drv[10]
port 2 nsew signal output
rlabel metal2 s 36726 39200 36782 40000 6 b0_drv[11]
port 3 nsew signal output
rlabel metal3 s 0 7488 800 7608 6 b0_drv[12]
port 4 nsew signal output
rlabel metal2 s 9678 39200 9734 40000 6 b0_drv[13]
port 5 nsew signal output
rlabel metal2 s 39302 39200 39358 40000 6 b0_drv[14]
port 6 nsew signal output
rlabel metal2 s 30286 0 30342 800 6 b0_drv[15]
port 7 nsew signal output
rlabel metal2 s 12898 39200 12954 40000 6 b0_drv[16]
port 8 nsew signal output
rlabel metal3 s 0 37408 800 37528 6 b0_drv[17]
port 9 nsew signal output
rlabel metal3 s 39200 6808 40000 6928 6 b0_drv[18]
port 10 nsew signal output
rlabel metal2 s 18694 0 18750 800 6 b0_drv[19]
port 11 nsew signal output
rlabel metal3 s 39200 22448 40000 22568 6 b0_drv[1]
port 12 nsew signal output
rlabel metal2 s 7746 39200 7802 40000 6 b0_drv[20]
port 13 nsew signal output
rlabel metal2 s 7102 39200 7158 40000 6 b0_drv[21]
port 14 nsew signal output
rlabel metal2 s 3238 0 3294 800 6 b0_drv[22]
port 15 nsew signal output
rlabel metal2 s 12254 39200 12310 40000 6 b0_drv[23]
port 16 nsew signal output
rlabel metal3 s 0 28568 800 28688 6 b0_drv[24]
port 17 nsew signal output
rlabel metal3 s 0 21088 800 21208 6 b0_drv[25]
port 18 nsew signal output
rlabel metal2 s 10322 39200 10378 40000 6 b0_drv[26]
port 19 nsew signal output
rlabel metal3 s 0 4768 800 4888 6 b0_drv[27]
port 20 nsew signal output
rlabel metal3 s 39200 25848 40000 25968 6 b0_drv[28]
port 21 nsew signal output
rlabel metal2 s 24490 0 24546 800 6 b0_drv[29]
port 22 nsew signal output
rlabel metal3 s 0 38088 800 38208 6 b0_drv[2]
port 23 nsew signal output
rlabel metal2 s 21270 39200 21326 40000 6 b0_drv[30]
port 24 nsew signal output
rlabel metal3 s 39200 4088 40000 4208 6 b0_drv[31]
port 25 nsew signal output
rlabel metal2 s 34794 0 34850 800 6 b0_drv[32]
port 26 nsew signal output
rlabel metal3 s 0 19728 800 19848 6 b0_drv[33]
port 27 nsew signal output
rlabel metal2 s 2594 39200 2650 40000 6 b0_drv[34]
port 28 nsew signal output
rlabel metal2 s 33506 39200 33562 40000 6 b0_drv[35]
port 29 nsew signal output
rlabel metal2 s 20626 39200 20682 40000 6 b0_drv[36]
port 30 nsew signal output
rlabel metal2 s 29642 39200 29698 40000 6 b0_drv[37]
port 31 nsew signal output
rlabel metal3 s 0 6808 800 6928 6 b0_drv[38]
port 32 nsew signal output
rlabel metal3 s 0 1368 800 1488 6 b0_drv[39]
port 33 nsew signal output
rlabel metal3 s 39200 8848 40000 8968 6 b0_drv[3]
port 34 nsew signal output
rlabel metal2 s 14186 39200 14242 40000 6 b0_drv[40]
port 35 nsew signal output
rlabel metal3 s 39200 34688 40000 34808 6 b0_drv[41]
port 36 nsew signal output
rlabel metal3 s 0 8848 800 8968 6 b0_drv[42]
port 37 nsew signal output
rlabel metal3 s 39200 37408 40000 37528 6 b0_drv[43]
port 38 nsew signal output
rlabel metal3 s 0 29248 800 29368 6 b0_drv[44]
port 39 nsew signal output
rlabel metal2 s 9034 0 9090 800 6 b0_drv[45]
port 40 nsew signal output
rlabel metal2 s 6458 0 6514 800 6 b0_drv[46]
port 41 nsew signal output
rlabel metal3 s 39200 11568 40000 11688 6 b0_drv[47]
port 42 nsew signal output
rlabel metal2 s 23846 39200 23902 40000 6 b0_drv[48]
port 43 nsew signal output
rlabel metal3 s 0 36728 800 36848 6 b0_drv[49]
port 44 nsew signal output
rlabel metal3 s 0 23128 800 23248 6 b0_drv[4]
port 45 nsew signal output
rlabel metal3 s 0 25168 800 25288 6 b0_drv[50]
port 46 nsew signal output
rlabel metal2 s 8390 39200 8446 40000 6 b0_drv[51]
port 47 nsew signal output
rlabel metal3 s 0 14968 800 15088 6 b0_drv[52]
port 48 nsew signal output
rlabel metal3 s 0 4088 800 4208 6 b0_drv[53]
port 49 nsew signal output
rlabel metal3 s 39200 3408 40000 3528 6 b0_drv[54]
port 50 nsew signal output
rlabel metal2 s 16762 39200 16818 40000 6 b0_drv[55]
port 51 nsew signal output
rlabel metal2 s 11610 0 11666 800 6 b0_drv[56]
port 52 nsew signal output
rlabel metal3 s 39200 38768 40000 38888 6 b0_drv[57]
port 53 nsew signal output
rlabel metal3 s 39200 10888 40000 11008 6 b0_drv[58]
port 54 nsew signal output
rlabel metal3 s 39200 33328 40000 33448 6 b0_drv[59]
port 55 nsew signal output
rlabel metal3 s 39200 15648 40000 15768 6 b0_drv[5]
port 56 nsew signal output
rlabel metal2 s 15474 39200 15530 40000 6 b0_drv[60]
port 57 nsew signal output
rlabel metal2 s 28354 0 28410 800 6 b0_drv[61]
port 58 nsew signal output
rlabel metal3 s 39200 34008 40000 34128 6 b0_drv[62]
port 59 nsew signal output
rlabel metal2 s 27066 0 27122 800 6 b0_drv[63]
port 60 nsew signal output
rlabel metal2 s 34794 39200 34850 40000 6 b0_drv[64]
port 61 nsew signal output
rlabel metal2 s 36082 39200 36138 40000 6 b0_drv[65]
port 62 nsew signal output
rlabel metal2 s 37370 39200 37426 40000 6 b0_drv[66]
port 63 nsew signal output
rlabel metal2 s 16118 39200 16174 40000 6 b0_drv[67]
port 64 nsew signal output
rlabel metal2 s 17406 0 17462 800 6 b0_drv[68]
port 65 nsew signal output
rlabel metal3 s 0 12928 800 13048 6 b0_drv[69]
port 66 nsew signal output
rlabel metal2 s 34150 39200 34206 40000 6 b0_drv[6]
port 67 nsew signal output
rlabel metal3 s 39200 28568 40000 28688 6 b0_drv[70]
port 68 nsew signal output
rlabel metal2 s 10966 0 11022 800 6 b0_drv[71]
port 69 nsew signal output
rlabel metal2 s 32862 0 32918 800 6 b0_drv[72]
port 70 nsew signal output
rlabel metal3 s 0 39448 800 39568 6 b0_drv[73]
port 71 nsew signal output
rlabel metal3 s 0 15648 800 15768 6 b0_drv[74]
port 72 nsew signal output
rlabel metal3 s 39200 17688 40000 17808 6 b0_drv[75]
port 73 nsew signal output
rlabel metal3 s 39200 5448 40000 5568 6 b0_drv[76]
port 74 nsew signal output
rlabel metal2 s 37370 0 37426 800 6 b0_drv[77]
port 75 nsew signal output
rlabel metal3 s 39200 20408 40000 20528 6 b0_drv[78]
port 76 nsew signal output
rlabel metal3 s 0 688 800 808 6 b0_drv[79]
port 77 nsew signal output
rlabel metal2 s 25134 0 25190 800 6 b0_drv[7]
port 78 nsew signal output
rlabel metal2 s 13542 39200 13598 40000 6 b0_drv[80]
port 79 nsew signal output
rlabel metal2 s 29642 0 29698 800 6 b0_drv[81]
port 80 nsew signal output
rlabel metal2 s 31574 39200 31630 40000 6 b0_drv[82]
port 81 nsew signal output
rlabel metal2 s 21914 39200 21970 40000 6 b0_drv[8]
port 82 nsew signal output
rlabel metal3 s 39200 29248 40000 29368 6 b0_drv[9]
port 83 nsew signal output
rlabel metal2 s 1306 0 1362 800 6 cw_clk_i
port 84 nsew signal input
rlabel metal2 s 12254 0 12310 800 6 cw_clk_o
port 85 nsew signal output
rlabel metal3 s 39200 688 40000 808 6 cw_dir
port 86 nsew signal input
rlabel metal3 s 39200 8 40000 128 6 cw_dir_b_o
port 87 nsew signal input
rlabel metal2 s 14830 0 14886 800 6 cw_dir_b_oo
port 88 nsew signal output
rlabel metal3 s 0 22448 800 22568 6 cw_dir_o
port 89 nsew signal output
rlabel metal2 s 32218 0 32274 800 6 cw_req_i
port 90 nsew signal input
rlabel metal3 s 0 26528 800 26648 6 cw_req_o
port 91 nsew signal output
rlabel metal3 s 39200 19728 40000 19848 6 cw_rst_i
port 92 nsew signal input
rlabel metal2 s 662 39200 718 40000 6 cw_rst_o
port 93 nsew signal output
rlabel metal3 s 0 10208 800 10328 6 i_pin_rst
port 94 nsew signal input
rlabel metal2 s 26422 39200 26478 40000 6 i_wb_rst
port 95 nsew signal input
rlabel metal2 s 30930 0 30986 800 6 io_oeb_15_0[0]
port 96 nsew signal output
rlabel metal3 s 39200 36728 40000 36848 6 io_oeb_15_0[10]
port 97 nsew signal output
rlabel metal2 s 13542 0 13598 800 6 io_oeb_15_0[11]
port 98 nsew signal output
rlabel metal3 s 0 34008 800 34128 6 io_oeb_15_0[12]
port 99 nsew signal output
rlabel metal3 s 39200 31968 40000 32088 6 io_oeb_15_0[13]
port 100 nsew signal output
rlabel metal2 s 1950 39200 2006 40000 6 io_oeb_15_0[14]
port 101 nsew signal output
rlabel metal3 s 39200 12928 40000 13048 6 io_oeb_15_0[15]
port 102 nsew signal output
rlabel metal2 s 4526 39200 4582 40000 6 io_oeb_15_0[1]
port 103 nsew signal output
rlabel metal3 s 39200 21088 40000 21208 6 io_oeb_15_0[2]
port 104 nsew signal output
rlabel metal2 s 38658 0 38714 800 6 io_oeb_15_0[3]
port 105 nsew signal output
rlabel metal2 s 21270 0 21326 800 6 io_oeb_15_0[4]
port 106 nsew signal output
rlabel metal3 s 39200 23128 40000 23248 6 io_oeb_15_0[5]
port 107 nsew signal output
rlabel metal2 s 19982 0 20038 800 6 io_oeb_15_0[6]
port 108 nsew signal output
rlabel metal2 s 8390 0 8446 800 6 io_oeb_15_0[7]
port 109 nsew signal output
rlabel metal2 s 18050 39200 18106 40000 6 io_oeb_15_0[8]
port 110 nsew signal output
rlabel metal3 s 0 20408 800 20528 6 io_oeb_15_0[9]
port 111 nsew signal output
rlabel metal2 s 36082 0 36138 800 6 io_oeb_18_16[0]
port 112 nsew signal output
rlabel metal3 s 0 29928 800 30048 6 io_oeb_18_16[1]
port 113 nsew signal output
rlabel metal3 s 39200 14968 40000 15088 6 io_oeb_18_16[2]
port 114 nsew signal output
rlabel metal3 s 0 17008 800 17128 6 io_oeb_20_19[0]
port 115 nsew signal output
rlabel metal2 s 24490 39200 24546 40000 6 io_oeb_20_19[1]
port 116 nsew signal output
rlabel metal2 s 23202 39200 23258 40000 6 io_oeb_21
port 117 nsew signal output
rlabel metal3 s 0 31968 800 32088 6 io_oeb_22
port 118 nsew signal output
rlabel metal2 s 5814 0 5870 800 6 io_out[0]
port 119 nsew signal output
rlabel metal3 s 39200 6128 40000 6248 6 io_out[10]
port 120 nsew signal output
rlabel metal2 s 16762 0 16818 800 6 io_out[11]
port 121 nsew signal output
rlabel metal3 s 39200 31288 40000 31408 6 io_out[12]
port 122 nsew signal output
rlabel metal3 s 39200 23808 40000 23928 6 io_out[13]
port 123 nsew signal output
rlabel metal3 s 0 17688 800 17808 6 io_out[14]
port 124 nsew signal output
rlabel metal2 s 3882 0 3938 800 6 io_out[1]
port 125 nsew signal output
rlabel metal3 s 39200 9528 40000 9648 6 io_out[2]
port 126 nsew signal output
rlabel metal3 s 0 35368 800 35488 6 io_out[3]
port 127 nsew signal output
rlabel metal2 s 10966 39200 11022 40000 6 io_out[4]
port 128 nsew signal output
rlabel metal3 s 39200 17008 40000 17128 6 io_out[5]
port 129 nsew signal output
rlabel metal3 s 39200 1368 40000 1488 6 io_out[6]
port 130 nsew signal output
rlabel metal3 s 0 2048 800 2168 6 io_out[7]
port 131 nsew signal output
rlabel metal3 s 39200 30608 40000 30728 6 io_out[8]
port 132 nsew signal output
rlabel metal2 s 28998 39200 29054 40000 6 io_out[9]
port 133 nsew signal output
rlabel metal2 s 9678 0 9734 800 6 io_out_20_19[0]
port 134 nsew signal output
rlabel metal3 s 39200 12248 40000 12368 6 io_out_20_19[1]
port 135 nsew signal output
rlabel metal2 s 25778 0 25834 800 6 io_out_22
port 136 nsew signal output
rlabel metal3 s 39200 2728 40000 2848 6 la_data_out_16_17[0]
port 137 nsew signal output
rlabel metal2 s 3238 39200 3294 40000 6 la_data_out_16_17[1]
port 138 nsew signal output
rlabel metal2 s 33506 0 33562 800 6 la_data_out_21
port 139 nsew signal output
rlabel metal2 s 4526 0 4582 800 6 la_data_out_37_36[0]
port 140 nsew signal output
rlabel metal2 s 16118 0 16174 800 6 la_data_out_37_36[1]
port 141 nsew signal output
rlabel metal3 s 0 14288 800 14408 6 la_data_out_77_62[0]
port 142 nsew signal output
rlabel metal3 s 39200 36048 40000 36168 6 la_data_out_77_62[10]
port 143 nsew signal output
rlabel metal3 s 39200 25168 40000 25288 6 la_data_out_77_62[11]
port 144 nsew signal output
rlabel metal2 s 35438 0 35494 800 6 la_data_out_77_62[12]
port 145 nsew signal output
rlabel metal3 s 0 18368 800 18488 6 la_data_out_77_62[13]
port 146 nsew signal output
rlabel metal3 s 39200 14288 40000 14408 6 la_data_out_77_62[14]
port 147 nsew signal output
rlabel metal2 s 662 0 718 800 6 la_data_out_77_62[15]
port 148 nsew signal output
rlabel metal3 s 0 12248 800 12368 6 la_data_out_77_62[1]
port 149 nsew signal output
rlabel metal3 s 39200 39448 40000 39568 6 la_data_out_77_62[2]
port 150 nsew signal output
rlabel metal2 s 38014 0 38070 800 6 la_data_out_77_62[3]
port 151 nsew signal output
rlabel metal2 s 38658 39200 38714 40000 6 la_data_out_77_62[4]
port 152 nsew signal output
rlabel metal3 s 0 25848 800 25968 6 la_data_out_77_62[5]
port 153 nsew signal output
rlabel metal3 s 0 27208 800 27328 6 la_data_out_77_62[6]
port 154 nsew signal output
rlabel metal2 s 23846 0 23902 800 6 la_data_out_77_62[7]
port 155 nsew signal output
rlabel metal2 s 18 0 74 800 6 la_data_out_77_62[8]
port 156 nsew signal output
rlabel metal3 s 0 3408 800 3528 6 la_data_out_77_62[9]
port 157 nsew signal output
rlabel metal3 s 0 31288 800 31408 6 la_data_out_97_95[0]
port 158 nsew signal output
rlabel metal2 s 5170 39200 5226 40000 6 la_data_out_97_95[1]
port 159 nsew signal output
rlabel metal2 s 19338 39200 19394 40000 6 la_data_out_97_95[2]
port 160 nsew signal output
rlabel metal3 s 0 23808 800 23928 6 la_datb_i[0]
port 161 nsew signal input
rlabel metal3 s 0 11568 800 11688 6 la_datb_i[1]
port 162 nsew signal input
rlabel metal2 s 1950 0 2006 800 6 la_datb_i[2]
port 163 nsew signal input
rlabel metal2 s 27066 39200 27122 40000 6 la_datb_o[0]
port 164 nsew signal output
rlabel metal2 s 18694 39200 18750 40000 6 la_datb_o[1]
port 165 nsew signal output
rlabel metal2 s 19338 0 19394 800 6 la_datb_o[2]
port 166 nsew signal output
rlabel metal2 s 32218 39200 32274 40000 6 o_s_rst
port 167 nsew signal output
rlabel metal3 s 39200 8168 40000 8288 6 oeb_out[0]
port 168 nsew signal output
rlabel metal3 s 0 32648 800 32768 6 oeb_out[10]
port 169 nsew signal output
rlabel metal3 s 39200 27888 40000 28008 6 oeb_out[11]
port 170 nsew signal output
rlabel metal2 s 7102 0 7158 800 6 oeb_out[12]
port 171 nsew signal output
rlabel metal2 s 14186 0 14242 800 6 oeb_out[13]
port 172 nsew signal output
rlabel metal2 s 21914 0 21970 800 6 oeb_out[14]
port 173 nsew signal output
rlabel metal3 s 39200 26528 40000 26648 6 oeb_out[1]
port 174 nsew signal output
rlabel metal2 s 22558 0 22614 800 6 oeb_out[2]
port 175 nsew signal output
rlabel metal3 s 0 6128 800 6248 6 oeb_out[3]
port 176 nsew signal output
rlabel metal2 s 28354 39200 28410 40000 6 oeb_out[4]
port 177 nsew signal output
rlabel metal2 s 18 39200 74 40000 6 oeb_out[5]
port 178 nsew signal output
rlabel metal2 s 5814 39200 5870 40000 6 oeb_out[6]
port 179 nsew signal output
rlabel metal2 s 27710 0 27766 800 6 oeb_out[7]
port 180 nsew signal output
rlabel metal3 s 0 9528 800 9648 6 oeb_out[8]
port 181 nsew signal output
rlabel metal3 s 0 34688 800 34808 6 oeb_out[9]
port 182 nsew signal output
rlabel metal3 s 39200 18368 40000 18488 6 soft_rst
port 183 nsew signal input
rlabel metal4 s 4208 2128 4528 37584 6 vccd1
port 184 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 37584 6 vccd1
port 184 nsew power bidirectional
rlabel metal4 s 19568 2128 19888 37584 6 vssd1
port 185 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 40000 40000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 685570
string GDS_FILE /home/piotro/ppcpu_caravel/openlane/uprj_w_const/runs/22_09_13_14_02/results/signoff/uprj_w_const.magic.gds
string GDS_START 60140
<< end >>

