VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO core0
  CLASS BLOCK ;
  FOREIGN core0 ;
  ORIGIN 0.000 0.000 ;
  SIZE 400.000 BY 820.000 ;
  PIN dbg_pc[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 112.240 400.000 112.840 ;
    END
  END dbg_pc[0]
  PIN dbg_pc[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 513.440 400.000 514.040 ;
    END
  END dbg_pc[10]
  PIN dbg_pc[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 547.440 400.000 548.040 ;
    END
  END dbg_pc[11]
  PIN dbg_pc[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 581.440 400.000 582.040 ;
    END
  END dbg_pc[12]
  PIN dbg_pc[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 615.440 400.000 616.040 ;
    END
  END dbg_pc[13]
  PIN dbg_pc[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 649.440 400.000 650.040 ;
    END
  END dbg_pc[14]
  PIN dbg_pc[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 683.440 400.000 684.040 ;
    END
  END dbg_pc[15]
  PIN dbg_pc[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 156.440 400.000 157.040 ;
    END
  END dbg_pc[1]
  PIN dbg_pc[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 200.640 400.000 201.240 ;
    END
  END dbg_pc[2]
  PIN dbg_pc[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 241.440 400.000 242.040 ;
    END
  END dbg_pc[3]
  PIN dbg_pc[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 282.240 400.000 282.840 ;
    END
  END dbg_pc[4]
  PIN dbg_pc[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 323.040 400.000 323.640 ;
    END
  END dbg_pc[5]
  PIN dbg_pc[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 363.840 400.000 364.440 ;
    END
  END dbg_pc[6]
  PIN dbg_pc[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 404.640 400.000 405.240 ;
    END
  END dbg_pc[7]
  PIN dbg_pc[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 445.440 400.000 446.040 ;
    END
  END dbg_pc[8]
  PIN dbg_pc[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 479.440 400.000 480.040 ;
    END
  END dbg_pc[9]
  PIN dbg_r0[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 115.640 400.000 116.240 ;
    END
  END dbg_r0[0]
  PIN dbg_r0[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 516.840 400.000 517.440 ;
    END
  END dbg_r0[10]
  PIN dbg_r0[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 550.840 400.000 551.440 ;
    END
  END dbg_r0[11]
  PIN dbg_r0[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 584.840 400.000 585.440 ;
    END
  END dbg_r0[12]
  PIN dbg_r0[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 618.840 400.000 619.440 ;
    END
  END dbg_r0[13]
  PIN dbg_r0[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 652.840 400.000 653.440 ;
    END
  END dbg_r0[14]
  PIN dbg_r0[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 686.840 400.000 687.440 ;
    END
  END dbg_r0[15]
  PIN dbg_r0[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 159.840 400.000 160.440 ;
    END
  END dbg_r0[1]
  PIN dbg_r0[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 204.040 400.000 204.640 ;
    END
  END dbg_r0[2]
  PIN dbg_r0[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 244.840 400.000 245.440 ;
    END
  END dbg_r0[3]
  PIN dbg_r0[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 285.640 400.000 286.240 ;
    END
  END dbg_r0[4]
  PIN dbg_r0[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 326.440 400.000 327.040 ;
    END
  END dbg_r0[5]
  PIN dbg_r0[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 367.240 400.000 367.840 ;
    END
  END dbg_r0[6]
  PIN dbg_r0[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 408.040 400.000 408.640 ;
    END
  END dbg_r0[7]
  PIN dbg_r0[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 448.840 400.000 449.440 ;
    END
  END dbg_r0[8]
  PIN dbg_r0[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 482.840 400.000 483.440 ;
    END
  END dbg_r0[9]
  PIN i_clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 51.040 400.000 51.640 ;
    END
  END i_clk
  PIN i_core_int_sreg[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 119.040 400.000 119.640 ;
    END
  END i_core_int_sreg[0]
  PIN i_core_int_sreg[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 520.240 400.000 520.840 ;
    END
  END i_core_int_sreg[10]
  PIN i_core_int_sreg[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 554.240 400.000 554.840 ;
    END
  END i_core_int_sreg[11]
  PIN i_core_int_sreg[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 588.240 400.000 588.840 ;
    END
  END i_core_int_sreg[12]
  PIN i_core_int_sreg[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 622.240 400.000 622.840 ;
    END
  END i_core_int_sreg[13]
  PIN i_core_int_sreg[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 656.240 400.000 656.840 ;
    END
  END i_core_int_sreg[14]
  PIN i_core_int_sreg[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 690.240 400.000 690.840 ;
    END
  END i_core_int_sreg[15]
  PIN i_core_int_sreg[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 163.240 400.000 163.840 ;
    END
  END i_core_int_sreg[1]
  PIN i_core_int_sreg[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 207.440 400.000 208.040 ;
    END
  END i_core_int_sreg[2]
  PIN i_core_int_sreg[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 248.240 400.000 248.840 ;
    END
  END i_core_int_sreg[3]
  PIN i_core_int_sreg[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 289.040 400.000 289.640 ;
    END
  END i_core_int_sreg[4]
  PIN i_core_int_sreg[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 329.840 400.000 330.440 ;
    END
  END i_core_int_sreg[5]
  PIN i_core_int_sreg[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 370.640 400.000 371.240 ;
    END
  END i_core_int_sreg[6]
  PIN i_core_int_sreg[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 411.440 400.000 412.040 ;
    END
  END i_core_int_sreg[7]
  PIN i_core_int_sreg[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 452.240 400.000 452.840 ;
    END
  END i_core_int_sreg[8]
  PIN i_core_int_sreg[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 486.240 400.000 486.840 ;
    END
  END i_core_int_sreg[9]
  PIN i_disable
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 54.440 400.000 55.040 ;
    END
  END i_disable
  PIN i_irq
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 57.840 400.000 58.440 ;
    END
  END i_irq
  PIN i_mc_core_int
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 61.240 400.000 61.840 ;
    END
  END i_mc_core_int
  PIN i_mem_ack
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 64.640 400.000 65.240 ;
    END
  END i_mem_ack
  PIN i_mem_data[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 122.440 400.000 123.040 ;
    END
  END i_mem_data[0]
  PIN i_mem_data[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 523.640 400.000 524.240 ;
    END
  END i_mem_data[10]
  PIN i_mem_data[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 557.640 400.000 558.240 ;
    END
  END i_mem_data[11]
  PIN i_mem_data[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 591.640 400.000 592.240 ;
    END
  END i_mem_data[12]
  PIN i_mem_data[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 625.640 400.000 626.240 ;
    END
  END i_mem_data[13]
  PIN i_mem_data[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 659.640 400.000 660.240 ;
    END
  END i_mem_data[14]
  PIN i_mem_data[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 693.640 400.000 694.240 ;
    END
  END i_mem_data[15]
  PIN i_mem_data[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 166.640 400.000 167.240 ;
    END
  END i_mem_data[1]
  PIN i_mem_data[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 210.840 400.000 211.440 ;
    END
  END i_mem_data[2]
  PIN i_mem_data[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 251.640 400.000 252.240 ;
    END
  END i_mem_data[3]
  PIN i_mem_data[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 292.440 400.000 293.040 ;
    END
  END i_mem_data[4]
  PIN i_mem_data[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 333.240 400.000 333.840 ;
    END
  END i_mem_data[5]
  PIN i_mem_data[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 374.040 400.000 374.640 ;
    END
  END i_mem_data[6]
  PIN i_mem_data[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 414.840 400.000 415.440 ;
    END
  END i_mem_data[7]
  PIN i_mem_data[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 455.640 400.000 456.240 ;
    END
  END i_mem_data[8]
  PIN i_mem_data[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 489.640 400.000 490.240 ;
    END
  END i_mem_data[9]
  PIN i_mem_exception
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 68.040 400.000 68.640 ;
    END
  END i_mem_exception
  PIN i_req_data[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 125.840 400.000 126.440 ;
    END
  END i_req_data[0]
  PIN i_req_data[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 527.040 400.000 527.640 ;
    END
  END i_req_data[10]
  PIN i_req_data[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 561.040 400.000 561.640 ;
    END
  END i_req_data[11]
  PIN i_req_data[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 595.040 400.000 595.640 ;
    END
  END i_req_data[12]
  PIN i_req_data[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 629.040 400.000 629.640 ;
    END
  END i_req_data[13]
  PIN i_req_data[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 663.040 400.000 663.640 ;
    END
  END i_req_data[14]
  PIN i_req_data[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 697.040 400.000 697.640 ;
    END
  END i_req_data[15]
  PIN i_req_data[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 717.440 400.000 718.040 ;
    END
  END i_req_data[16]
  PIN i_req_data[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 720.840 400.000 721.440 ;
    END
  END i_req_data[17]
  PIN i_req_data[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 724.240 400.000 724.840 ;
    END
  END i_req_data[18]
  PIN i_req_data[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 727.640 400.000 728.240 ;
    END
  END i_req_data[19]
  PIN i_req_data[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 170.040 400.000 170.640 ;
    END
  END i_req_data[1]
  PIN i_req_data[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 731.040 400.000 731.640 ;
    END
  END i_req_data[20]
  PIN i_req_data[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 734.440 400.000 735.040 ;
    END
  END i_req_data[21]
  PIN i_req_data[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 737.840 400.000 738.440 ;
    END
  END i_req_data[22]
  PIN i_req_data[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 741.240 400.000 741.840 ;
    END
  END i_req_data[23]
  PIN i_req_data[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 744.640 400.000 745.240 ;
    END
  END i_req_data[24]
  PIN i_req_data[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 748.040 400.000 748.640 ;
    END
  END i_req_data[25]
  PIN i_req_data[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 751.440 400.000 752.040 ;
    END
  END i_req_data[26]
  PIN i_req_data[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 754.840 400.000 755.440 ;
    END
  END i_req_data[27]
  PIN i_req_data[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 758.240 400.000 758.840 ;
    END
  END i_req_data[28]
  PIN i_req_data[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 761.640 400.000 762.240 ;
    END
  END i_req_data[29]
  PIN i_req_data[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 214.240 400.000 214.840 ;
    END
  END i_req_data[2]
  PIN i_req_data[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 765.040 400.000 765.640 ;
    END
  END i_req_data[30]
  PIN i_req_data[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 768.440 400.000 769.040 ;
    END
  END i_req_data[31]
  PIN i_req_data[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 255.040 400.000 255.640 ;
    END
  END i_req_data[3]
  PIN i_req_data[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 295.840 400.000 296.440 ;
    END
  END i_req_data[4]
  PIN i_req_data[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 336.640 400.000 337.240 ;
    END
  END i_req_data[5]
  PIN i_req_data[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 377.440 400.000 378.040 ;
    END
  END i_req_data[6]
  PIN i_req_data[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 418.240 400.000 418.840 ;
    END
  END i_req_data[7]
  PIN i_req_data[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 459.040 400.000 459.640 ;
    END
  END i_req_data[8]
  PIN i_req_data[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 493.040 400.000 493.640 ;
    END
  END i_req_data[9]
  PIN i_req_data_valid
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 71.440 400.000 72.040 ;
    END
  END i_req_data_valid
  PIN i_rst
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 74.840 400.000 75.440 ;
    END
  END i_rst
  PIN o_c_data_page
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 78.240 400.000 78.840 ;
    END
  END o_c_data_page
  PIN o_c_instr_long
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 81.640 400.000 82.240 ;
    END
  END o_c_instr_long
  PIN o_c_instr_page
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 85.040 400.000 85.640 ;
    END
  END o_c_instr_page
  PIN o_icache_flush
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 88.440 400.000 89.040 ;
    END
  END o_icache_flush
  PIN o_instr_long_addr[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 129.240 400.000 129.840 ;
    END
  END o_instr_long_addr[0]
  PIN o_instr_long_addr[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 173.440 400.000 174.040 ;
    END
  END o_instr_long_addr[1]
  PIN o_instr_long_addr[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 217.640 400.000 218.240 ;
    END
  END o_instr_long_addr[2]
  PIN o_instr_long_addr[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 258.440 400.000 259.040 ;
    END
  END o_instr_long_addr[3]
  PIN o_instr_long_addr[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 299.240 400.000 299.840 ;
    END
  END o_instr_long_addr[4]
  PIN o_instr_long_addr[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 340.040 400.000 340.640 ;
    END
  END o_instr_long_addr[5]
  PIN o_instr_long_addr[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 380.840 400.000 381.440 ;
    END
  END o_instr_long_addr[6]
  PIN o_instr_long_addr[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 421.640 400.000 422.240 ;
    END
  END o_instr_long_addr[7]
  PIN o_mem_addr[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 132.640 400.000 133.240 ;
    END
  END o_mem_addr[0]
  PIN o_mem_addr[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 530.440 400.000 531.040 ;
    END
  END o_mem_addr[10]
  PIN o_mem_addr[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 564.440 400.000 565.040 ;
    END
  END o_mem_addr[11]
  PIN o_mem_addr[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 598.440 400.000 599.040 ;
    END
  END o_mem_addr[12]
  PIN o_mem_addr[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 632.440 400.000 633.040 ;
    END
  END o_mem_addr[13]
  PIN o_mem_addr[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 666.440 400.000 667.040 ;
    END
  END o_mem_addr[14]
  PIN o_mem_addr[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 700.440 400.000 701.040 ;
    END
  END o_mem_addr[15]
  PIN o_mem_addr[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 176.840 400.000 177.440 ;
    END
  END o_mem_addr[1]
  PIN o_mem_addr[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 221.040 400.000 221.640 ;
    END
  END o_mem_addr[2]
  PIN o_mem_addr[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 261.840 400.000 262.440 ;
    END
  END o_mem_addr[3]
  PIN o_mem_addr[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 302.640 400.000 303.240 ;
    END
  END o_mem_addr[4]
  PIN o_mem_addr[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 343.440 400.000 344.040 ;
    END
  END o_mem_addr[5]
  PIN o_mem_addr[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 384.240 400.000 384.840 ;
    END
  END o_mem_addr[6]
  PIN o_mem_addr[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 425.040 400.000 425.640 ;
    END
  END o_mem_addr[7]
  PIN o_mem_addr[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 462.440 400.000 463.040 ;
    END
  END o_mem_addr[8]
  PIN o_mem_addr[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 496.440 400.000 497.040 ;
    END
  END o_mem_addr[9]
  PIN o_mem_addr_high[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 136.040 400.000 136.640 ;
    END
  END o_mem_addr_high[0]
  PIN o_mem_addr_high[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 180.240 400.000 180.840 ;
    END
  END o_mem_addr_high[1]
  PIN o_mem_addr_high[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 224.440 400.000 225.040 ;
    END
  END o_mem_addr_high[2]
  PIN o_mem_addr_high[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 265.240 400.000 265.840 ;
    END
  END o_mem_addr_high[3]
  PIN o_mem_addr_high[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 306.040 400.000 306.640 ;
    END
  END o_mem_addr_high[4]
  PIN o_mem_addr_high[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 346.840 400.000 347.440 ;
    END
  END o_mem_addr_high[5]
  PIN o_mem_addr_high[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 387.640 400.000 388.240 ;
    END
  END o_mem_addr_high[6]
  PIN o_mem_addr_high[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 428.440 400.000 429.040 ;
    END
  END o_mem_addr_high[7]
  PIN o_mem_data[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 139.440 400.000 140.040 ;
    END
  END o_mem_data[0]
  PIN o_mem_data[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 533.840 400.000 534.440 ;
    END
  END o_mem_data[10]
  PIN o_mem_data[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 567.840 400.000 568.440 ;
    END
  END o_mem_data[11]
  PIN o_mem_data[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 601.840 400.000 602.440 ;
    END
  END o_mem_data[12]
  PIN o_mem_data[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 635.840 400.000 636.440 ;
    END
  END o_mem_data[13]
  PIN o_mem_data[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 669.840 400.000 670.440 ;
    END
  END o_mem_data[14]
  PIN o_mem_data[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 703.840 400.000 704.440 ;
    END
  END o_mem_data[15]
  PIN o_mem_data[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 183.640 400.000 184.240 ;
    END
  END o_mem_data[1]
  PIN o_mem_data[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 227.840 400.000 228.440 ;
    END
  END o_mem_data[2]
  PIN o_mem_data[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 268.640 400.000 269.240 ;
    END
  END o_mem_data[3]
  PIN o_mem_data[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 309.440 400.000 310.040 ;
    END
  END o_mem_data[4]
  PIN o_mem_data[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 350.240 400.000 350.840 ;
    END
  END o_mem_data[5]
  PIN o_mem_data[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 391.040 400.000 391.640 ;
    END
  END o_mem_data[6]
  PIN o_mem_data[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 431.840 400.000 432.440 ;
    END
  END o_mem_data[7]
  PIN o_mem_data[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 465.840 400.000 466.440 ;
    END
  END o_mem_data[8]
  PIN o_mem_data[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 499.840 400.000 500.440 ;
    END
  END o_mem_data[9]
  PIN o_mem_long
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 91.840 400.000 92.440 ;
    END
  END o_mem_long
  PIN o_mem_req
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 95.240 400.000 95.840 ;
    END
  END o_mem_req
  PIN o_mem_sel[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 142.840 400.000 143.440 ;
    END
  END o_mem_sel[0]
  PIN o_mem_sel[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 187.040 400.000 187.640 ;
    END
  END o_mem_sel[1]
  PIN o_mem_we
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 98.640 400.000 99.240 ;
    END
  END o_mem_we
  PIN o_req_active
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 102.040 400.000 102.640 ;
    END
  END o_req_active
  PIN o_req_addr[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 146.240 400.000 146.840 ;
    END
  END o_req_addr[0]
  PIN o_req_addr[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 537.240 400.000 537.840 ;
    END
  END o_req_addr[10]
  PIN o_req_addr[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 571.240 400.000 571.840 ;
    END
  END o_req_addr[11]
  PIN o_req_addr[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 605.240 400.000 605.840 ;
    END
  END o_req_addr[12]
  PIN o_req_addr[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 639.240 400.000 639.840 ;
    END
  END o_req_addr[13]
  PIN o_req_addr[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 673.240 400.000 673.840 ;
    END
  END o_req_addr[14]
  PIN o_req_addr[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 707.240 400.000 707.840 ;
    END
  END o_req_addr[15]
  PIN o_req_addr[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 190.440 400.000 191.040 ;
    END
  END o_req_addr[1]
  PIN o_req_addr[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 231.240 400.000 231.840 ;
    END
  END o_req_addr[2]
  PIN o_req_addr[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 272.040 400.000 272.640 ;
    END
  END o_req_addr[3]
  PIN o_req_addr[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 312.840 400.000 313.440 ;
    END
  END o_req_addr[4]
  PIN o_req_addr[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 353.640 400.000 354.240 ;
    END
  END o_req_addr[5]
  PIN o_req_addr[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 394.440 400.000 395.040 ;
    END
  END o_req_addr[6]
  PIN o_req_addr[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 435.240 400.000 435.840 ;
    END
  END o_req_addr[7]
  PIN o_req_addr[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 469.240 400.000 469.840 ;
    END
  END o_req_addr[8]
  PIN o_req_addr[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 503.240 400.000 503.840 ;
    END
  END o_req_addr[9]
  PIN o_req_ppl_submit
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 105.440 400.000 106.040 ;
    END
  END o_req_ppl_submit
  PIN sr_bus_addr[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 149.640 400.000 150.240 ;
    END
  END sr_bus_addr[0]
  PIN sr_bus_addr[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 540.640 400.000 541.240 ;
    END
  END sr_bus_addr[10]
  PIN sr_bus_addr[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 574.640 400.000 575.240 ;
    END
  END sr_bus_addr[11]
  PIN sr_bus_addr[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 608.640 400.000 609.240 ;
    END
  END sr_bus_addr[12]
  PIN sr_bus_addr[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 642.640 400.000 643.240 ;
    END
  END sr_bus_addr[13]
  PIN sr_bus_addr[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 676.640 400.000 677.240 ;
    END
  END sr_bus_addr[14]
  PIN sr_bus_addr[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 710.640 400.000 711.240 ;
    END
  END sr_bus_addr[15]
  PIN sr_bus_addr[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 193.840 400.000 194.440 ;
    END
  END sr_bus_addr[1]
  PIN sr_bus_addr[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 234.640 400.000 235.240 ;
    END
  END sr_bus_addr[2]
  PIN sr_bus_addr[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 275.440 400.000 276.040 ;
    END
  END sr_bus_addr[3]
  PIN sr_bus_addr[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 316.240 400.000 316.840 ;
    END
  END sr_bus_addr[4]
  PIN sr_bus_addr[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 357.040 400.000 357.640 ;
    END
  END sr_bus_addr[5]
  PIN sr_bus_addr[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 397.840 400.000 398.440 ;
    END
  END sr_bus_addr[6]
  PIN sr_bus_addr[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 438.640 400.000 439.240 ;
    END
  END sr_bus_addr[7]
  PIN sr_bus_addr[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 472.640 400.000 473.240 ;
    END
  END sr_bus_addr[8]
  PIN sr_bus_addr[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 506.640 400.000 507.240 ;
    END
  END sr_bus_addr[9]
  PIN sr_bus_data_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 153.040 400.000 153.640 ;
    END
  END sr_bus_data_o[0]
  PIN sr_bus_data_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 544.040 400.000 544.640 ;
    END
  END sr_bus_data_o[10]
  PIN sr_bus_data_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 578.040 400.000 578.640 ;
    END
  END sr_bus_data_o[11]
  PIN sr_bus_data_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 612.040 400.000 612.640 ;
    END
  END sr_bus_data_o[12]
  PIN sr_bus_data_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 646.040 400.000 646.640 ;
    END
  END sr_bus_data_o[13]
  PIN sr_bus_data_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 680.040 400.000 680.640 ;
    END
  END sr_bus_data_o[14]
  PIN sr_bus_data_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 714.040 400.000 714.640 ;
    END
  END sr_bus_data_o[15]
  PIN sr_bus_data_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 197.240 400.000 197.840 ;
    END
  END sr_bus_data_o[1]
  PIN sr_bus_data_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 238.040 400.000 238.640 ;
    END
  END sr_bus_data_o[2]
  PIN sr_bus_data_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 278.840 400.000 279.440 ;
    END
  END sr_bus_data_o[3]
  PIN sr_bus_data_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 319.640 400.000 320.240 ;
    END
  END sr_bus_data_o[4]
  PIN sr_bus_data_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 360.440 400.000 361.040 ;
    END
  END sr_bus_data_o[5]
  PIN sr_bus_data_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 401.240 400.000 401.840 ;
    END
  END sr_bus_data_o[6]
  PIN sr_bus_data_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 442.040 400.000 442.640 ;
    END
  END sr_bus_data_o[7]
  PIN sr_bus_data_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 476.040 400.000 476.640 ;
    END
  END sr_bus_data_o[8]
  PIN sr_bus_data_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 510.040 400.000 510.640 ;
    END
  END sr_bus_data_o[9]
  PIN sr_bus_we
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 108.840 400.000 109.440 ;
    END
  END sr_bus_we
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 808.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 808.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 328.240 10.640 329.840 808.080 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 808.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 251.440 10.640 253.040 808.080 ;
    END
  END vssd1
  OBS
      LAYER nwell ;
        RECT 5.330 806.425 394.410 808.030 ;
        RECT 5.330 800.985 394.410 803.815 ;
        RECT 5.330 795.545 394.410 798.375 ;
        RECT 5.330 790.105 394.410 792.935 ;
        RECT 5.330 784.665 394.410 787.495 ;
        RECT 5.330 779.225 394.410 782.055 ;
        RECT 5.330 773.785 394.410 776.615 ;
        RECT 5.330 768.345 394.410 771.175 ;
        RECT 5.330 762.905 394.410 765.735 ;
        RECT 5.330 757.465 394.410 760.295 ;
        RECT 5.330 752.025 394.410 754.855 ;
        RECT 5.330 746.585 394.410 749.415 ;
        RECT 5.330 741.145 394.410 743.975 ;
        RECT 5.330 735.705 394.410 738.535 ;
        RECT 5.330 730.265 394.410 733.095 ;
        RECT 5.330 724.825 394.410 727.655 ;
        RECT 5.330 719.385 394.410 722.215 ;
        RECT 5.330 713.945 394.410 716.775 ;
        RECT 5.330 708.505 394.410 711.335 ;
        RECT 5.330 703.065 394.410 705.895 ;
        RECT 5.330 697.625 394.410 700.455 ;
        RECT 5.330 692.185 394.410 695.015 ;
        RECT 5.330 686.745 394.410 689.575 ;
        RECT 5.330 681.305 394.410 684.135 ;
        RECT 5.330 675.865 394.410 678.695 ;
        RECT 5.330 670.425 394.410 673.255 ;
        RECT 5.330 664.985 394.410 667.815 ;
        RECT 5.330 659.545 394.410 662.375 ;
        RECT 5.330 654.105 394.410 656.935 ;
        RECT 5.330 648.665 394.410 651.495 ;
        RECT 5.330 643.225 394.410 646.055 ;
        RECT 5.330 637.785 394.410 640.615 ;
        RECT 5.330 632.345 394.410 635.175 ;
        RECT 5.330 626.905 394.410 629.735 ;
        RECT 5.330 621.465 394.410 624.295 ;
        RECT 5.330 616.025 394.410 618.855 ;
        RECT 5.330 610.585 394.410 613.415 ;
        RECT 5.330 605.145 394.410 607.975 ;
        RECT 5.330 599.705 394.410 602.535 ;
        RECT 5.330 594.265 394.410 597.095 ;
        RECT 5.330 588.825 394.410 591.655 ;
        RECT 5.330 583.385 394.410 586.215 ;
        RECT 5.330 577.945 394.410 580.775 ;
        RECT 5.330 572.505 394.410 575.335 ;
        RECT 5.330 567.065 394.410 569.895 ;
        RECT 5.330 561.625 394.410 564.455 ;
        RECT 5.330 556.185 394.410 559.015 ;
        RECT 5.330 550.745 394.410 553.575 ;
        RECT 5.330 545.305 394.410 548.135 ;
        RECT 5.330 539.865 394.410 542.695 ;
        RECT 5.330 534.425 394.410 537.255 ;
        RECT 5.330 528.985 394.410 531.815 ;
        RECT 5.330 523.545 394.410 526.375 ;
        RECT 5.330 518.105 394.410 520.935 ;
        RECT 5.330 512.665 394.410 515.495 ;
        RECT 5.330 507.225 394.410 510.055 ;
        RECT 5.330 501.785 394.410 504.615 ;
        RECT 5.330 496.345 394.410 499.175 ;
        RECT 5.330 490.905 394.410 493.735 ;
        RECT 5.330 485.465 394.410 488.295 ;
        RECT 5.330 480.025 394.410 482.855 ;
        RECT 5.330 474.585 394.410 477.415 ;
        RECT 5.330 469.145 394.410 471.975 ;
        RECT 5.330 463.705 394.410 466.535 ;
        RECT 5.330 458.265 394.410 461.095 ;
        RECT 5.330 452.825 394.410 455.655 ;
        RECT 5.330 447.385 394.410 450.215 ;
        RECT 5.330 441.945 394.410 444.775 ;
        RECT 5.330 436.505 394.410 439.335 ;
        RECT 5.330 431.065 394.410 433.895 ;
        RECT 5.330 425.625 394.410 428.455 ;
        RECT 5.330 420.185 394.410 423.015 ;
        RECT 5.330 414.745 394.410 417.575 ;
        RECT 5.330 409.305 394.410 412.135 ;
        RECT 5.330 403.865 394.410 406.695 ;
        RECT 5.330 398.425 394.410 401.255 ;
        RECT 5.330 392.985 394.410 395.815 ;
        RECT 5.330 387.545 394.410 390.375 ;
        RECT 5.330 382.105 394.410 384.935 ;
        RECT 5.330 376.665 394.410 379.495 ;
        RECT 5.330 371.225 394.410 374.055 ;
        RECT 5.330 365.785 394.410 368.615 ;
        RECT 5.330 360.345 394.410 363.175 ;
        RECT 5.330 354.905 394.410 357.735 ;
        RECT 5.330 349.465 394.410 352.295 ;
        RECT 5.330 344.025 394.410 346.855 ;
        RECT 5.330 338.585 394.410 341.415 ;
        RECT 5.330 333.145 394.410 335.975 ;
        RECT 5.330 327.705 394.410 330.535 ;
        RECT 5.330 322.265 394.410 325.095 ;
        RECT 5.330 316.825 394.410 319.655 ;
        RECT 5.330 311.385 394.410 314.215 ;
        RECT 5.330 305.945 394.410 308.775 ;
        RECT 5.330 300.505 394.410 303.335 ;
        RECT 5.330 295.065 394.410 297.895 ;
        RECT 5.330 289.625 394.410 292.455 ;
        RECT 5.330 284.185 394.410 287.015 ;
        RECT 5.330 278.745 394.410 281.575 ;
        RECT 5.330 273.305 394.410 276.135 ;
        RECT 5.330 267.865 394.410 270.695 ;
        RECT 5.330 262.425 394.410 265.255 ;
        RECT 5.330 256.985 394.410 259.815 ;
        RECT 5.330 251.545 394.410 254.375 ;
        RECT 5.330 246.105 394.410 248.935 ;
        RECT 5.330 240.665 394.410 243.495 ;
        RECT 5.330 235.225 394.410 238.055 ;
        RECT 5.330 229.785 394.410 232.615 ;
        RECT 5.330 224.345 394.410 227.175 ;
        RECT 5.330 218.905 394.410 221.735 ;
        RECT 5.330 213.465 394.410 216.295 ;
        RECT 5.330 208.025 394.410 210.855 ;
        RECT 5.330 202.585 394.410 205.415 ;
        RECT 5.330 197.145 394.410 199.975 ;
        RECT 5.330 191.705 394.410 194.535 ;
        RECT 5.330 186.265 394.410 189.095 ;
        RECT 5.330 180.825 394.410 183.655 ;
        RECT 5.330 175.385 394.410 178.215 ;
        RECT 5.330 169.945 394.410 172.775 ;
        RECT 5.330 164.505 394.410 167.335 ;
        RECT 5.330 159.065 394.410 161.895 ;
        RECT 5.330 153.625 394.410 156.455 ;
        RECT 5.330 148.185 394.410 151.015 ;
        RECT 5.330 142.745 394.410 145.575 ;
        RECT 5.330 137.305 394.410 140.135 ;
        RECT 5.330 131.865 394.410 134.695 ;
        RECT 5.330 126.425 394.410 129.255 ;
        RECT 5.330 120.985 394.410 123.815 ;
        RECT 5.330 115.545 394.410 118.375 ;
        RECT 5.330 110.105 394.410 112.935 ;
        RECT 5.330 104.665 394.410 107.495 ;
        RECT 5.330 99.225 394.410 102.055 ;
        RECT 5.330 93.785 394.410 96.615 ;
        RECT 5.330 88.345 394.410 91.175 ;
        RECT 5.330 82.905 394.410 85.735 ;
        RECT 5.330 77.465 394.410 80.295 ;
        RECT 5.330 72.025 394.410 74.855 ;
        RECT 5.330 66.585 394.410 69.415 ;
        RECT 5.330 61.145 394.410 63.975 ;
        RECT 5.330 55.705 394.410 58.535 ;
        RECT 5.330 50.265 394.410 53.095 ;
        RECT 5.330 44.825 394.410 47.655 ;
        RECT 5.330 39.385 394.410 42.215 ;
        RECT 5.330 33.945 394.410 36.775 ;
        RECT 5.330 28.505 394.410 31.335 ;
        RECT 5.330 23.065 394.410 25.895 ;
        RECT 5.330 17.625 394.410 20.455 ;
        RECT 5.330 12.185 394.410 15.015 ;
      LAYER li1 ;
        RECT 5.520 10.795 394.220 807.925 ;
      LAYER met1 ;
        RECT 5.520 10.640 399.670 808.080 ;
      LAYER met2 ;
        RECT 21.070 10.695 399.640 808.025 ;
      LAYER met3 ;
        RECT 21.050 769.440 397.835 808.005 ;
        RECT 21.050 768.040 395.600 769.440 ;
        RECT 21.050 766.040 397.835 768.040 ;
        RECT 21.050 764.640 395.600 766.040 ;
        RECT 21.050 762.640 397.835 764.640 ;
        RECT 21.050 761.240 395.600 762.640 ;
        RECT 21.050 759.240 397.835 761.240 ;
        RECT 21.050 757.840 395.600 759.240 ;
        RECT 21.050 755.840 397.835 757.840 ;
        RECT 21.050 754.440 395.600 755.840 ;
        RECT 21.050 752.440 397.835 754.440 ;
        RECT 21.050 751.040 395.600 752.440 ;
        RECT 21.050 749.040 397.835 751.040 ;
        RECT 21.050 747.640 395.600 749.040 ;
        RECT 21.050 745.640 397.835 747.640 ;
        RECT 21.050 744.240 395.600 745.640 ;
        RECT 21.050 742.240 397.835 744.240 ;
        RECT 21.050 740.840 395.600 742.240 ;
        RECT 21.050 738.840 397.835 740.840 ;
        RECT 21.050 737.440 395.600 738.840 ;
        RECT 21.050 735.440 397.835 737.440 ;
        RECT 21.050 734.040 395.600 735.440 ;
        RECT 21.050 732.040 397.835 734.040 ;
        RECT 21.050 730.640 395.600 732.040 ;
        RECT 21.050 728.640 397.835 730.640 ;
        RECT 21.050 727.240 395.600 728.640 ;
        RECT 21.050 725.240 397.835 727.240 ;
        RECT 21.050 723.840 395.600 725.240 ;
        RECT 21.050 721.840 397.835 723.840 ;
        RECT 21.050 720.440 395.600 721.840 ;
        RECT 21.050 718.440 397.835 720.440 ;
        RECT 21.050 717.040 395.600 718.440 ;
        RECT 21.050 715.040 397.835 717.040 ;
        RECT 21.050 713.640 395.600 715.040 ;
        RECT 21.050 711.640 397.835 713.640 ;
        RECT 21.050 710.240 395.600 711.640 ;
        RECT 21.050 708.240 397.835 710.240 ;
        RECT 21.050 706.840 395.600 708.240 ;
        RECT 21.050 704.840 397.835 706.840 ;
        RECT 21.050 703.440 395.600 704.840 ;
        RECT 21.050 701.440 397.835 703.440 ;
        RECT 21.050 700.040 395.600 701.440 ;
        RECT 21.050 698.040 397.835 700.040 ;
        RECT 21.050 696.640 395.600 698.040 ;
        RECT 21.050 694.640 397.835 696.640 ;
        RECT 21.050 693.240 395.600 694.640 ;
        RECT 21.050 691.240 397.835 693.240 ;
        RECT 21.050 689.840 395.600 691.240 ;
        RECT 21.050 687.840 397.835 689.840 ;
        RECT 21.050 686.440 395.600 687.840 ;
        RECT 21.050 684.440 397.835 686.440 ;
        RECT 21.050 683.040 395.600 684.440 ;
        RECT 21.050 681.040 397.835 683.040 ;
        RECT 21.050 679.640 395.600 681.040 ;
        RECT 21.050 677.640 397.835 679.640 ;
        RECT 21.050 676.240 395.600 677.640 ;
        RECT 21.050 674.240 397.835 676.240 ;
        RECT 21.050 672.840 395.600 674.240 ;
        RECT 21.050 670.840 397.835 672.840 ;
        RECT 21.050 669.440 395.600 670.840 ;
        RECT 21.050 667.440 397.835 669.440 ;
        RECT 21.050 666.040 395.600 667.440 ;
        RECT 21.050 664.040 397.835 666.040 ;
        RECT 21.050 662.640 395.600 664.040 ;
        RECT 21.050 660.640 397.835 662.640 ;
        RECT 21.050 659.240 395.600 660.640 ;
        RECT 21.050 657.240 397.835 659.240 ;
        RECT 21.050 655.840 395.600 657.240 ;
        RECT 21.050 653.840 397.835 655.840 ;
        RECT 21.050 652.440 395.600 653.840 ;
        RECT 21.050 650.440 397.835 652.440 ;
        RECT 21.050 649.040 395.600 650.440 ;
        RECT 21.050 647.040 397.835 649.040 ;
        RECT 21.050 645.640 395.600 647.040 ;
        RECT 21.050 643.640 397.835 645.640 ;
        RECT 21.050 642.240 395.600 643.640 ;
        RECT 21.050 640.240 397.835 642.240 ;
        RECT 21.050 638.840 395.600 640.240 ;
        RECT 21.050 636.840 397.835 638.840 ;
        RECT 21.050 635.440 395.600 636.840 ;
        RECT 21.050 633.440 397.835 635.440 ;
        RECT 21.050 632.040 395.600 633.440 ;
        RECT 21.050 630.040 397.835 632.040 ;
        RECT 21.050 628.640 395.600 630.040 ;
        RECT 21.050 626.640 397.835 628.640 ;
        RECT 21.050 625.240 395.600 626.640 ;
        RECT 21.050 623.240 397.835 625.240 ;
        RECT 21.050 621.840 395.600 623.240 ;
        RECT 21.050 619.840 397.835 621.840 ;
        RECT 21.050 618.440 395.600 619.840 ;
        RECT 21.050 616.440 397.835 618.440 ;
        RECT 21.050 615.040 395.600 616.440 ;
        RECT 21.050 613.040 397.835 615.040 ;
        RECT 21.050 611.640 395.600 613.040 ;
        RECT 21.050 609.640 397.835 611.640 ;
        RECT 21.050 608.240 395.600 609.640 ;
        RECT 21.050 606.240 397.835 608.240 ;
        RECT 21.050 604.840 395.600 606.240 ;
        RECT 21.050 602.840 397.835 604.840 ;
        RECT 21.050 601.440 395.600 602.840 ;
        RECT 21.050 599.440 397.835 601.440 ;
        RECT 21.050 598.040 395.600 599.440 ;
        RECT 21.050 596.040 397.835 598.040 ;
        RECT 21.050 594.640 395.600 596.040 ;
        RECT 21.050 592.640 397.835 594.640 ;
        RECT 21.050 591.240 395.600 592.640 ;
        RECT 21.050 589.240 397.835 591.240 ;
        RECT 21.050 587.840 395.600 589.240 ;
        RECT 21.050 585.840 397.835 587.840 ;
        RECT 21.050 584.440 395.600 585.840 ;
        RECT 21.050 582.440 397.835 584.440 ;
        RECT 21.050 581.040 395.600 582.440 ;
        RECT 21.050 579.040 397.835 581.040 ;
        RECT 21.050 577.640 395.600 579.040 ;
        RECT 21.050 575.640 397.835 577.640 ;
        RECT 21.050 574.240 395.600 575.640 ;
        RECT 21.050 572.240 397.835 574.240 ;
        RECT 21.050 570.840 395.600 572.240 ;
        RECT 21.050 568.840 397.835 570.840 ;
        RECT 21.050 567.440 395.600 568.840 ;
        RECT 21.050 565.440 397.835 567.440 ;
        RECT 21.050 564.040 395.600 565.440 ;
        RECT 21.050 562.040 397.835 564.040 ;
        RECT 21.050 560.640 395.600 562.040 ;
        RECT 21.050 558.640 397.835 560.640 ;
        RECT 21.050 557.240 395.600 558.640 ;
        RECT 21.050 555.240 397.835 557.240 ;
        RECT 21.050 553.840 395.600 555.240 ;
        RECT 21.050 551.840 397.835 553.840 ;
        RECT 21.050 550.440 395.600 551.840 ;
        RECT 21.050 548.440 397.835 550.440 ;
        RECT 21.050 547.040 395.600 548.440 ;
        RECT 21.050 545.040 397.835 547.040 ;
        RECT 21.050 543.640 395.600 545.040 ;
        RECT 21.050 541.640 397.835 543.640 ;
        RECT 21.050 540.240 395.600 541.640 ;
        RECT 21.050 538.240 397.835 540.240 ;
        RECT 21.050 536.840 395.600 538.240 ;
        RECT 21.050 534.840 397.835 536.840 ;
        RECT 21.050 533.440 395.600 534.840 ;
        RECT 21.050 531.440 397.835 533.440 ;
        RECT 21.050 530.040 395.600 531.440 ;
        RECT 21.050 528.040 397.835 530.040 ;
        RECT 21.050 526.640 395.600 528.040 ;
        RECT 21.050 524.640 397.835 526.640 ;
        RECT 21.050 523.240 395.600 524.640 ;
        RECT 21.050 521.240 397.835 523.240 ;
        RECT 21.050 519.840 395.600 521.240 ;
        RECT 21.050 517.840 397.835 519.840 ;
        RECT 21.050 516.440 395.600 517.840 ;
        RECT 21.050 514.440 397.835 516.440 ;
        RECT 21.050 513.040 395.600 514.440 ;
        RECT 21.050 511.040 397.835 513.040 ;
        RECT 21.050 509.640 395.600 511.040 ;
        RECT 21.050 507.640 397.835 509.640 ;
        RECT 21.050 506.240 395.600 507.640 ;
        RECT 21.050 504.240 397.835 506.240 ;
        RECT 21.050 502.840 395.600 504.240 ;
        RECT 21.050 500.840 397.835 502.840 ;
        RECT 21.050 499.440 395.600 500.840 ;
        RECT 21.050 497.440 397.835 499.440 ;
        RECT 21.050 496.040 395.600 497.440 ;
        RECT 21.050 494.040 397.835 496.040 ;
        RECT 21.050 492.640 395.600 494.040 ;
        RECT 21.050 490.640 397.835 492.640 ;
        RECT 21.050 489.240 395.600 490.640 ;
        RECT 21.050 487.240 397.835 489.240 ;
        RECT 21.050 485.840 395.600 487.240 ;
        RECT 21.050 483.840 397.835 485.840 ;
        RECT 21.050 482.440 395.600 483.840 ;
        RECT 21.050 480.440 397.835 482.440 ;
        RECT 21.050 479.040 395.600 480.440 ;
        RECT 21.050 477.040 397.835 479.040 ;
        RECT 21.050 475.640 395.600 477.040 ;
        RECT 21.050 473.640 397.835 475.640 ;
        RECT 21.050 472.240 395.600 473.640 ;
        RECT 21.050 470.240 397.835 472.240 ;
        RECT 21.050 468.840 395.600 470.240 ;
        RECT 21.050 466.840 397.835 468.840 ;
        RECT 21.050 465.440 395.600 466.840 ;
        RECT 21.050 463.440 397.835 465.440 ;
        RECT 21.050 462.040 395.600 463.440 ;
        RECT 21.050 460.040 397.835 462.040 ;
        RECT 21.050 458.640 395.600 460.040 ;
        RECT 21.050 456.640 397.835 458.640 ;
        RECT 21.050 455.240 395.600 456.640 ;
        RECT 21.050 453.240 397.835 455.240 ;
        RECT 21.050 451.840 395.600 453.240 ;
        RECT 21.050 449.840 397.835 451.840 ;
        RECT 21.050 448.440 395.600 449.840 ;
        RECT 21.050 446.440 397.835 448.440 ;
        RECT 21.050 445.040 395.600 446.440 ;
        RECT 21.050 443.040 397.835 445.040 ;
        RECT 21.050 441.640 395.600 443.040 ;
        RECT 21.050 439.640 397.835 441.640 ;
        RECT 21.050 438.240 395.600 439.640 ;
        RECT 21.050 436.240 397.835 438.240 ;
        RECT 21.050 434.840 395.600 436.240 ;
        RECT 21.050 432.840 397.835 434.840 ;
        RECT 21.050 431.440 395.600 432.840 ;
        RECT 21.050 429.440 397.835 431.440 ;
        RECT 21.050 428.040 395.600 429.440 ;
        RECT 21.050 426.040 397.835 428.040 ;
        RECT 21.050 424.640 395.600 426.040 ;
        RECT 21.050 422.640 397.835 424.640 ;
        RECT 21.050 421.240 395.600 422.640 ;
        RECT 21.050 419.240 397.835 421.240 ;
        RECT 21.050 417.840 395.600 419.240 ;
        RECT 21.050 415.840 397.835 417.840 ;
        RECT 21.050 414.440 395.600 415.840 ;
        RECT 21.050 412.440 397.835 414.440 ;
        RECT 21.050 411.040 395.600 412.440 ;
        RECT 21.050 409.040 397.835 411.040 ;
        RECT 21.050 407.640 395.600 409.040 ;
        RECT 21.050 405.640 397.835 407.640 ;
        RECT 21.050 404.240 395.600 405.640 ;
        RECT 21.050 402.240 397.835 404.240 ;
        RECT 21.050 400.840 395.600 402.240 ;
        RECT 21.050 398.840 397.835 400.840 ;
        RECT 21.050 397.440 395.600 398.840 ;
        RECT 21.050 395.440 397.835 397.440 ;
        RECT 21.050 394.040 395.600 395.440 ;
        RECT 21.050 392.040 397.835 394.040 ;
        RECT 21.050 390.640 395.600 392.040 ;
        RECT 21.050 388.640 397.835 390.640 ;
        RECT 21.050 387.240 395.600 388.640 ;
        RECT 21.050 385.240 397.835 387.240 ;
        RECT 21.050 383.840 395.600 385.240 ;
        RECT 21.050 381.840 397.835 383.840 ;
        RECT 21.050 380.440 395.600 381.840 ;
        RECT 21.050 378.440 397.835 380.440 ;
        RECT 21.050 377.040 395.600 378.440 ;
        RECT 21.050 375.040 397.835 377.040 ;
        RECT 21.050 373.640 395.600 375.040 ;
        RECT 21.050 371.640 397.835 373.640 ;
        RECT 21.050 370.240 395.600 371.640 ;
        RECT 21.050 368.240 397.835 370.240 ;
        RECT 21.050 366.840 395.600 368.240 ;
        RECT 21.050 364.840 397.835 366.840 ;
        RECT 21.050 363.440 395.600 364.840 ;
        RECT 21.050 361.440 397.835 363.440 ;
        RECT 21.050 360.040 395.600 361.440 ;
        RECT 21.050 358.040 397.835 360.040 ;
        RECT 21.050 356.640 395.600 358.040 ;
        RECT 21.050 354.640 397.835 356.640 ;
        RECT 21.050 353.240 395.600 354.640 ;
        RECT 21.050 351.240 397.835 353.240 ;
        RECT 21.050 349.840 395.600 351.240 ;
        RECT 21.050 347.840 397.835 349.840 ;
        RECT 21.050 346.440 395.600 347.840 ;
        RECT 21.050 344.440 397.835 346.440 ;
        RECT 21.050 343.040 395.600 344.440 ;
        RECT 21.050 341.040 397.835 343.040 ;
        RECT 21.050 339.640 395.600 341.040 ;
        RECT 21.050 337.640 397.835 339.640 ;
        RECT 21.050 336.240 395.600 337.640 ;
        RECT 21.050 334.240 397.835 336.240 ;
        RECT 21.050 332.840 395.600 334.240 ;
        RECT 21.050 330.840 397.835 332.840 ;
        RECT 21.050 329.440 395.600 330.840 ;
        RECT 21.050 327.440 397.835 329.440 ;
        RECT 21.050 326.040 395.600 327.440 ;
        RECT 21.050 324.040 397.835 326.040 ;
        RECT 21.050 322.640 395.600 324.040 ;
        RECT 21.050 320.640 397.835 322.640 ;
        RECT 21.050 319.240 395.600 320.640 ;
        RECT 21.050 317.240 397.835 319.240 ;
        RECT 21.050 315.840 395.600 317.240 ;
        RECT 21.050 313.840 397.835 315.840 ;
        RECT 21.050 312.440 395.600 313.840 ;
        RECT 21.050 310.440 397.835 312.440 ;
        RECT 21.050 309.040 395.600 310.440 ;
        RECT 21.050 307.040 397.835 309.040 ;
        RECT 21.050 305.640 395.600 307.040 ;
        RECT 21.050 303.640 397.835 305.640 ;
        RECT 21.050 302.240 395.600 303.640 ;
        RECT 21.050 300.240 397.835 302.240 ;
        RECT 21.050 298.840 395.600 300.240 ;
        RECT 21.050 296.840 397.835 298.840 ;
        RECT 21.050 295.440 395.600 296.840 ;
        RECT 21.050 293.440 397.835 295.440 ;
        RECT 21.050 292.040 395.600 293.440 ;
        RECT 21.050 290.040 397.835 292.040 ;
        RECT 21.050 288.640 395.600 290.040 ;
        RECT 21.050 286.640 397.835 288.640 ;
        RECT 21.050 285.240 395.600 286.640 ;
        RECT 21.050 283.240 397.835 285.240 ;
        RECT 21.050 281.840 395.600 283.240 ;
        RECT 21.050 279.840 397.835 281.840 ;
        RECT 21.050 278.440 395.600 279.840 ;
        RECT 21.050 276.440 397.835 278.440 ;
        RECT 21.050 275.040 395.600 276.440 ;
        RECT 21.050 273.040 397.835 275.040 ;
        RECT 21.050 271.640 395.600 273.040 ;
        RECT 21.050 269.640 397.835 271.640 ;
        RECT 21.050 268.240 395.600 269.640 ;
        RECT 21.050 266.240 397.835 268.240 ;
        RECT 21.050 264.840 395.600 266.240 ;
        RECT 21.050 262.840 397.835 264.840 ;
        RECT 21.050 261.440 395.600 262.840 ;
        RECT 21.050 259.440 397.835 261.440 ;
        RECT 21.050 258.040 395.600 259.440 ;
        RECT 21.050 256.040 397.835 258.040 ;
        RECT 21.050 254.640 395.600 256.040 ;
        RECT 21.050 252.640 397.835 254.640 ;
        RECT 21.050 251.240 395.600 252.640 ;
        RECT 21.050 249.240 397.835 251.240 ;
        RECT 21.050 247.840 395.600 249.240 ;
        RECT 21.050 245.840 397.835 247.840 ;
        RECT 21.050 244.440 395.600 245.840 ;
        RECT 21.050 242.440 397.835 244.440 ;
        RECT 21.050 241.040 395.600 242.440 ;
        RECT 21.050 239.040 397.835 241.040 ;
        RECT 21.050 237.640 395.600 239.040 ;
        RECT 21.050 235.640 397.835 237.640 ;
        RECT 21.050 234.240 395.600 235.640 ;
        RECT 21.050 232.240 397.835 234.240 ;
        RECT 21.050 230.840 395.600 232.240 ;
        RECT 21.050 228.840 397.835 230.840 ;
        RECT 21.050 227.440 395.600 228.840 ;
        RECT 21.050 225.440 397.835 227.440 ;
        RECT 21.050 224.040 395.600 225.440 ;
        RECT 21.050 222.040 397.835 224.040 ;
        RECT 21.050 220.640 395.600 222.040 ;
        RECT 21.050 218.640 397.835 220.640 ;
        RECT 21.050 217.240 395.600 218.640 ;
        RECT 21.050 215.240 397.835 217.240 ;
        RECT 21.050 213.840 395.600 215.240 ;
        RECT 21.050 211.840 397.835 213.840 ;
        RECT 21.050 210.440 395.600 211.840 ;
        RECT 21.050 208.440 397.835 210.440 ;
        RECT 21.050 207.040 395.600 208.440 ;
        RECT 21.050 205.040 397.835 207.040 ;
        RECT 21.050 203.640 395.600 205.040 ;
        RECT 21.050 201.640 397.835 203.640 ;
        RECT 21.050 200.240 395.600 201.640 ;
        RECT 21.050 198.240 397.835 200.240 ;
        RECT 21.050 196.840 395.600 198.240 ;
        RECT 21.050 194.840 397.835 196.840 ;
        RECT 21.050 193.440 395.600 194.840 ;
        RECT 21.050 191.440 397.835 193.440 ;
        RECT 21.050 190.040 395.600 191.440 ;
        RECT 21.050 188.040 397.835 190.040 ;
        RECT 21.050 186.640 395.600 188.040 ;
        RECT 21.050 184.640 397.835 186.640 ;
        RECT 21.050 183.240 395.600 184.640 ;
        RECT 21.050 181.240 397.835 183.240 ;
        RECT 21.050 179.840 395.600 181.240 ;
        RECT 21.050 177.840 397.835 179.840 ;
        RECT 21.050 176.440 395.600 177.840 ;
        RECT 21.050 174.440 397.835 176.440 ;
        RECT 21.050 173.040 395.600 174.440 ;
        RECT 21.050 171.040 397.835 173.040 ;
        RECT 21.050 169.640 395.600 171.040 ;
        RECT 21.050 167.640 397.835 169.640 ;
        RECT 21.050 166.240 395.600 167.640 ;
        RECT 21.050 164.240 397.835 166.240 ;
        RECT 21.050 162.840 395.600 164.240 ;
        RECT 21.050 160.840 397.835 162.840 ;
        RECT 21.050 159.440 395.600 160.840 ;
        RECT 21.050 157.440 397.835 159.440 ;
        RECT 21.050 156.040 395.600 157.440 ;
        RECT 21.050 154.040 397.835 156.040 ;
        RECT 21.050 152.640 395.600 154.040 ;
        RECT 21.050 150.640 397.835 152.640 ;
        RECT 21.050 149.240 395.600 150.640 ;
        RECT 21.050 147.240 397.835 149.240 ;
        RECT 21.050 145.840 395.600 147.240 ;
        RECT 21.050 143.840 397.835 145.840 ;
        RECT 21.050 142.440 395.600 143.840 ;
        RECT 21.050 140.440 397.835 142.440 ;
        RECT 21.050 139.040 395.600 140.440 ;
        RECT 21.050 137.040 397.835 139.040 ;
        RECT 21.050 135.640 395.600 137.040 ;
        RECT 21.050 133.640 397.835 135.640 ;
        RECT 21.050 132.240 395.600 133.640 ;
        RECT 21.050 130.240 397.835 132.240 ;
        RECT 21.050 128.840 395.600 130.240 ;
        RECT 21.050 126.840 397.835 128.840 ;
        RECT 21.050 125.440 395.600 126.840 ;
        RECT 21.050 123.440 397.835 125.440 ;
        RECT 21.050 122.040 395.600 123.440 ;
        RECT 21.050 120.040 397.835 122.040 ;
        RECT 21.050 118.640 395.600 120.040 ;
        RECT 21.050 116.640 397.835 118.640 ;
        RECT 21.050 115.240 395.600 116.640 ;
        RECT 21.050 113.240 397.835 115.240 ;
        RECT 21.050 111.840 395.600 113.240 ;
        RECT 21.050 109.840 397.835 111.840 ;
        RECT 21.050 108.440 395.600 109.840 ;
        RECT 21.050 106.440 397.835 108.440 ;
        RECT 21.050 105.040 395.600 106.440 ;
        RECT 21.050 103.040 397.835 105.040 ;
        RECT 21.050 101.640 395.600 103.040 ;
        RECT 21.050 99.640 397.835 101.640 ;
        RECT 21.050 98.240 395.600 99.640 ;
        RECT 21.050 96.240 397.835 98.240 ;
        RECT 21.050 94.840 395.600 96.240 ;
        RECT 21.050 92.840 397.835 94.840 ;
        RECT 21.050 91.440 395.600 92.840 ;
        RECT 21.050 89.440 397.835 91.440 ;
        RECT 21.050 88.040 395.600 89.440 ;
        RECT 21.050 86.040 397.835 88.040 ;
        RECT 21.050 84.640 395.600 86.040 ;
        RECT 21.050 82.640 397.835 84.640 ;
        RECT 21.050 81.240 395.600 82.640 ;
        RECT 21.050 79.240 397.835 81.240 ;
        RECT 21.050 77.840 395.600 79.240 ;
        RECT 21.050 75.840 397.835 77.840 ;
        RECT 21.050 74.440 395.600 75.840 ;
        RECT 21.050 72.440 397.835 74.440 ;
        RECT 21.050 71.040 395.600 72.440 ;
        RECT 21.050 69.040 397.835 71.040 ;
        RECT 21.050 67.640 395.600 69.040 ;
        RECT 21.050 65.640 397.835 67.640 ;
        RECT 21.050 64.240 395.600 65.640 ;
        RECT 21.050 62.240 397.835 64.240 ;
        RECT 21.050 60.840 395.600 62.240 ;
        RECT 21.050 58.840 397.835 60.840 ;
        RECT 21.050 57.440 395.600 58.840 ;
        RECT 21.050 55.440 397.835 57.440 ;
        RECT 21.050 54.040 395.600 55.440 ;
        RECT 21.050 52.040 397.835 54.040 ;
        RECT 21.050 50.640 395.600 52.040 ;
        RECT 21.050 10.715 397.835 50.640 ;
      LAYER met4 ;
        RECT 177.855 47.775 251.040 792.705 ;
        RECT 253.440 47.775 327.840 792.705 ;
        RECT 330.240 47.775 386.105 792.705 ;
  END
END core0
END LIBRARY

