magic
tech sky130A
magscale 1 2
timestamp 1672342418
<< obsli1 >>
rect 1104 2159 288880 277457
<< obsm1 >>
rect 290 2128 289970 277976
<< obsm2 >>
rect 296 2139 289966 278361
<< metal3 >>
rect 0 270512 800 270632
rect 0 268472 800 268592
rect 0 266432 800 266552
rect 0 264392 800 264512
rect 0 262352 800 262472
rect 0 260312 800 260432
rect 0 258272 800 258392
rect 0 256232 800 256352
rect 0 254192 800 254312
rect 0 252152 800 252272
rect 0 250112 800 250232
rect 0 248072 800 248192
rect 0 246032 800 246152
rect 0 243992 800 244112
rect 0 241952 800 242072
rect 0 239912 800 240032
rect 0 237872 800 237992
rect 0 235832 800 235952
rect 0 233792 800 233912
rect 0 231752 800 231872
rect 0 229712 800 229832
rect 0 227672 800 227792
rect 0 225632 800 225752
rect 0 223592 800 223712
rect 0 221552 800 221672
rect 0 219512 800 219632
rect 0 217472 800 217592
rect 0 215432 800 215552
rect 0 213392 800 213512
rect 0 211352 800 211472
rect 0 209312 800 209432
rect 0 207272 800 207392
rect 0 205232 800 205352
rect 0 203192 800 203312
rect 0 201152 800 201272
rect 0 199112 800 199232
rect 0 197072 800 197192
rect 0 195032 800 195152
rect 0 192992 800 193112
rect 0 190952 800 191072
rect 0 188912 800 189032
rect 0 186872 800 186992
rect 0 184832 800 184952
rect 0 182792 800 182912
rect 0 180752 800 180872
rect 0 178712 800 178832
rect 0 176672 800 176792
rect 0 174632 800 174752
rect 0 172592 800 172712
rect 0 170552 800 170672
rect 0 168512 800 168632
rect 0 166472 800 166592
rect 0 164432 800 164552
rect 0 162392 800 162512
rect 0 160352 800 160472
rect 0 158312 800 158432
rect 0 156272 800 156392
rect 0 154232 800 154352
rect 0 152192 800 152312
rect 0 150152 800 150272
rect 0 148112 800 148232
rect 0 146072 800 146192
rect 0 144032 800 144152
rect 0 141992 800 142112
rect 0 139952 800 140072
rect 0 137912 800 138032
rect 0 135872 800 135992
rect 0 133832 800 133952
rect 0 131792 800 131912
rect 0 129752 800 129872
rect 0 127712 800 127832
rect 0 125672 800 125792
rect 0 123632 800 123752
rect 0 121592 800 121712
rect 0 119552 800 119672
rect 0 117512 800 117632
rect 0 115472 800 115592
rect 0 113432 800 113552
rect 0 111392 800 111512
rect 0 109352 800 109472
rect 0 107312 800 107432
rect 0 105272 800 105392
rect 0 103232 800 103352
rect 0 101192 800 101312
rect 0 99152 800 99272
rect 0 97112 800 97232
rect 0 95072 800 95192
rect 0 93032 800 93152
rect 0 90992 800 91112
rect 0 88952 800 89072
rect 0 86912 800 87032
rect 0 84872 800 84992
rect 0 82832 800 82952
rect 0 80792 800 80912
rect 0 78752 800 78872
rect 0 76712 800 76832
rect 0 74672 800 74792
rect 0 72632 800 72752
rect 0 70592 800 70712
rect 0 68552 800 68672
rect 0 66512 800 66632
rect 0 64472 800 64592
rect 0 62432 800 62552
rect 0 60392 800 60512
rect 0 58352 800 58472
rect 0 56312 800 56432
rect 0 54272 800 54392
rect 0 52232 800 52352
rect 0 50192 800 50312
rect 0 48152 800 48272
rect 0 46112 800 46232
rect 0 44072 800 44192
rect 0 42032 800 42152
rect 0 39992 800 40112
rect 0 37952 800 38072
rect 0 35912 800 36032
rect 0 33872 800 33992
rect 0 31832 800 31952
rect 0 29792 800 29912
rect 0 27752 800 27872
rect 0 25712 800 25832
rect 0 23672 800 23792
rect 0 21632 800 21752
rect 0 19592 800 19712
rect 0 17552 800 17672
rect 0 15512 800 15632
rect 0 13472 800 13592
rect 0 11432 800 11552
rect 0 9392 800 9512
<< obsm3 >>
rect 422 270712 289971 278357
rect 880 270432 289971 270712
rect 422 268672 289971 270432
rect 880 268392 289971 268672
rect 422 266632 289971 268392
rect 880 266352 289971 266632
rect 422 264592 289971 266352
rect 880 264312 289971 264592
rect 422 262552 289971 264312
rect 880 262272 289971 262552
rect 422 260512 289971 262272
rect 880 260232 289971 260512
rect 422 258472 289971 260232
rect 880 258192 289971 258472
rect 422 256432 289971 258192
rect 880 256152 289971 256432
rect 422 254392 289971 256152
rect 880 254112 289971 254392
rect 422 252352 289971 254112
rect 880 252072 289971 252352
rect 422 250312 289971 252072
rect 880 250032 289971 250312
rect 422 248272 289971 250032
rect 880 247992 289971 248272
rect 422 246232 289971 247992
rect 880 245952 289971 246232
rect 422 244192 289971 245952
rect 880 243912 289971 244192
rect 422 242152 289971 243912
rect 880 241872 289971 242152
rect 422 240112 289971 241872
rect 880 239832 289971 240112
rect 422 238072 289971 239832
rect 880 237792 289971 238072
rect 422 236032 289971 237792
rect 880 235752 289971 236032
rect 422 233992 289971 235752
rect 880 233712 289971 233992
rect 422 231952 289971 233712
rect 880 231672 289971 231952
rect 422 229912 289971 231672
rect 880 229632 289971 229912
rect 422 227872 289971 229632
rect 880 227592 289971 227872
rect 422 225832 289971 227592
rect 880 225552 289971 225832
rect 422 223792 289971 225552
rect 880 223512 289971 223792
rect 422 221752 289971 223512
rect 880 221472 289971 221752
rect 422 219712 289971 221472
rect 880 219432 289971 219712
rect 422 217672 289971 219432
rect 880 217392 289971 217672
rect 422 215632 289971 217392
rect 880 215352 289971 215632
rect 422 213592 289971 215352
rect 880 213312 289971 213592
rect 422 211552 289971 213312
rect 880 211272 289971 211552
rect 422 209512 289971 211272
rect 880 209232 289971 209512
rect 422 207472 289971 209232
rect 880 207192 289971 207472
rect 422 205432 289971 207192
rect 880 205152 289971 205432
rect 422 203392 289971 205152
rect 880 203112 289971 203392
rect 422 201352 289971 203112
rect 880 201072 289971 201352
rect 422 199312 289971 201072
rect 880 199032 289971 199312
rect 422 197272 289971 199032
rect 880 196992 289971 197272
rect 422 195232 289971 196992
rect 880 194952 289971 195232
rect 422 193192 289971 194952
rect 880 192912 289971 193192
rect 422 191152 289971 192912
rect 880 190872 289971 191152
rect 422 189112 289971 190872
rect 880 188832 289971 189112
rect 422 187072 289971 188832
rect 880 186792 289971 187072
rect 422 185032 289971 186792
rect 880 184752 289971 185032
rect 422 182992 289971 184752
rect 880 182712 289971 182992
rect 422 180952 289971 182712
rect 880 180672 289971 180952
rect 422 178912 289971 180672
rect 880 178632 289971 178912
rect 422 176872 289971 178632
rect 880 176592 289971 176872
rect 422 174832 289971 176592
rect 880 174552 289971 174832
rect 422 172792 289971 174552
rect 880 172512 289971 172792
rect 422 170752 289971 172512
rect 880 170472 289971 170752
rect 422 168712 289971 170472
rect 880 168432 289971 168712
rect 422 166672 289971 168432
rect 880 166392 289971 166672
rect 422 164632 289971 166392
rect 880 164352 289971 164632
rect 422 162592 289971 164352
rect 880 162312 289971 162592
rect 422 160552 289971 162312
rect 880 160272 289971 160552
rect 422 158512 289971 160272
rect 880 158232 289971 158512
rect 422 156472 289971 158232
rect 880 156192 289971 156472
rect 422 154432 289971 156192
rect 880 154152 289971 154432
rect 422 152392 289971 154152
rect 880 152112 289971 152392
rect 422 150352 289971 152112
rect 880 150072 289971 150352
rect 422 148312 289971 150072
rect 880 148032 289971 148312
rect 422 146272 289971 148032
rect 880 145992 289971 146272
rect 422 144232 289971 145992
rect 880 143952 289971 144232
rect 422 142192 289971 143952
rect 880 141912 289971 142192
rect 422 140152 289971 141912
rect 880 139872 289971 140152
rect 422 138112 289971 139872
rect 880 137832 289971 138112
rect 422 136072 289971 137832
rect 880 135792 289971 136072
rect 422 134032 289971 135792
rect 880 133752 289971 134032
rect 422 131992 289971 133752
rect 880 131712 289971 131992
rect 422 129952 289971 131712
rect 880 129672 289971 129952
rect 422 127912 289971 129672
rect 880 127632 289971 127912
rect 422 125872 289971 127632
rect 880 125592 289971 125872
rect 422 123832 289971 125592
rect 880 123552 289971 123832
rect 422 121792 289971 123552
rect 880 121512 289971 121792
rect 422 119752 289971 121512
rect 880 119472 289971 119752
rect 422 117712 289971 119472
rect 880 117432 289971 117712
rect 422 115672 289971 117432
rect 880 115392 289971 115672
rect 422 113632 289971 115392
rect 880 113352 289971 113632
rect 422 111592 289971 113352
rect 880 111312 289971 111592
rect 422 109552 289971 111312
rect 880 109272 289971 109552
rect 422 107512 289971 109272
rect 880 107232 289971 107512
rect 422 105472 289971 107232
rect 880 105192 289971 105472
rect 422 103432 289971 105192
rect 880 103152 289971 103432
rect 422 101392 289971 103152
rect 880 101112 289971 101392
rect 422 99352 289971 101112
rect 880 99072 289971 99352
rect 422 97312 289971 99072
rect 880 97032 289971 97312
rect 422 95272 289971 97032
rect 880 94992 289971 95272
rect 422 93232 289971 94992
rect 880 92952 289971 93232
rect 422 91192 289971 92952
rect 880 90912 289971 91192
rect 422 89152 289971 90912
rect 880 88872 289971 89152
rect 422 87112 289971 88872
rect 880 86832 289971 87112
rect 422 85072 289971 86832
rect 880 84792 289971 85072
rect 422 83032 289971 84792
rect 880 82752 289971 83032
rect 422 80992 289971 82752
rect 880 80712 289971 80992
rect 422 78952 289971 80712
rect 880 78672 289971 78952
rect 422 76912 289971 78672
rect 880 76632 289971 76912
rect 422 74872 289971 76632
rect 880 74592 289971 74872
rect 422 72832 289971 74592
rect 880 72552 289971 72832
rect 422 70792 289971 72552
rect 880 70512 289971 70792
rect 422 68752 289971 70512
rect 880 68472 289971 68752
rect 422 66712 289971 68472
rect 880 66432 289971 66712
rect 422 64672 289971 66432
rect 880 64392 289971 64672
rect 422 62632 289971 64392
rect 880 62352 289971 62632
rect 422 60592 289971 62352
rect 880 60312 289971 60592
rect 422 58552 289971 60312
rect 880 58272 289971 58552
rect 422 56512 289971 58272
rect 880 56232 289971 56512
rect 422 54472 289971 56232
rect 880 54192 289971 54472
rect 422 52432 289971 54192
rect 880 52152 289971 52432
rect 422 50392 289971 52152
rect 880 50112 289971 50392
rect 422 48352 289971 50112
rect 880 48072 289971 48352
rect 422 46312 289971 48072
rect 880 46032 289971 46312
rect 422 44272 289971 46032
rect 880 43992 289971 44272
rect 422 42232 289971 43992
rect 880 41952 289971 42232
rect 422 40192 289971 41952
rect 880 39912 289971 40192
rect 422 38152 289971 39912
rect 880 37872 289971 38152
rect 422 36112 289971 37872
rect 880 35832 289971 36112
rect 422 34072 289971 35832
rect 880 33792 289971 34072
rect 422 32032 289971 33792
rect 880 31752 289971 32032
rect 422 29992 289971 31752
rect 880 29712 289971 29992
rect 422 27952 289971 29712
rect 880 27672 289971 27952
rect 422 25912 289971 27672
rect 880 25632 289971 25912
rect 422 23872 289971 25632
rect 880 23592 289971 23872
rect 422 21832 289971 23592
rect 880 21552 289971 21832
rect 422 19792 289971 21552
rect 880 19512 289971 19792
rect 422 17752 289971 19512
rect 880 17472 289971 17752
rect 422 15712 289971 17472
rect 880 15432 289971 15712
rect 422 13672 289971 15432
rect 880 13392 289971 13672
rect 422 11632 289971 13392
rect 880 11352 289971 11632
rect 422 9592 289971 11352
rect 880 9312 289971 9592
rect 422 2143 289971 9312
<< metal4 >>
rect 4208 2128 4528 277488
rect 19568 2128 19888 277488
rect 34928 2128 35248 277488
rect 50288 2128 50608 277488
rect 65648 2128 65968 277488
rect 81008 2128 81328 277488
rect 96368 2128 96688 277488
rect 111728 2128 112048 277488
rect 127088 2128 127408 277488
rect 142448 2128 142768 277488
rect 157808 2128 158128 277488
rect 173168 2128 173488 277488
rect 188528 2128 188848 277488
rect 203888 2128 204208 277488
rect 219248 2128 219568 277488
rect 234608 2128 234928 277488
rect 249968 2128 250288 277488
rect 265328 2128 265648 277488
rect 280688 2128 281008 277488
<< obsm4 >>
rect 427 277568 289189 278357
rect 427 5067 4128 277568
rect 4608 5067 19488 277568
rect 19968 5067 34848 277568
rect 35328 5067 50208 277568
rect 50688 5067 65568 277568
rect 66048 5067 80928 277568
rect 81408 5067 96288 277568
rect 96768 5067 111648 277568
rect 112128 5067 127008 277568
rect 127488 5067 142368 277568
rect 142848 5067 157728 277568
rect 158208 5067 173088 277568
rect 173568 5067 188448 277568
rect 188928 5067 203808 277568
rect 204288 5067 219168 277568
rect 219648 5067 234528 277568
rect 235008 5067 249888 277568
rect 250368 5067 265248 277568
rect 265728 5067 280608 277568
rect 281088 5067 289189 277568
<< labels >>
rlabel metal3 s 0 9392 800 9512 6 i_clk
port 1 nsew signal input
rlabel metal3 s 0 11432 800 11552 6 i_rst
port 2 nsew signal input
rlabel metal3 s 0 13472 800 13592 6 mem_ack
port 3 nsew signal output
rlabel metal3 s 0 35912 800 36032 6 mem_addr[0]
port 4 nsew signal input
rlabel metal3 s 0 166472 800 166592 6 mem_addr[10]
port 5 nsew signal input
rlabel metal3 s 0 178712 800 178832 6 mem_addr[11]
port 6 nsew signal input
rlabel metal3 s 0 190952 800 191072 6 mem_addr[12]
port 7 nsew signal input
rlabel metal3 s 0 203192 800 203312 6 mem_addr[13]
port 8 nsew signal input
rlabel metal3 s 0 215432 800 215552 6 mem_addr[14]
port 9 nsew signal input
rlabel metal3 s 0 227672 800 227792 6 mem_addr[15]
port 10 nsew signal input
rlabel metal3 s 0 239912 800 240032 6 mem_addr[16]
port 11 nsew signal input
rlabel metal3 s 0 243992 800 244112 6 mem_addr[17]
port 12 nsew signal input
rlabel metal3 s 0 248072 800 248192 6 mem_addr[18]
port 13 nsew signal input
rlabel metal3 s 0 252152 800 252272 6 mem_addr[19]
port 14 nsew signal input
rlabel metal3 s 0 52232 800 52352 6 mem_addr[1]
port 15 nsew signal input
rlabel metal3 s 0 256232 800 256352 6 mem_addr[20]
port 16 nsew signal input
rlabel metal3 s 0 260312 800 260432 6 mem_addr[21]
port 17 nsew signal input
rlabel metal3 s 0 264392 800 264512 6 mem_addr[22]
port 18 nsew signal input
rlabel metal3 s 0 268472 800 268592 6 mem_addr[23]
port 19 nsew signal input
rlabel metal3 s 0 68552 800 68672 6 mem_addr[2]
port 20 nsew signal input
rlabel metal3 s 0 80792 800 80912 6 mem_addr[3]
port 21 nsew signal input
rlabel metal3 s 0 93032 800 93152 6 mem_addr[4]
port 22 nsew signal input
rlabel metal3 s 0 105272 800 105392 6 mem_addr[5]
port 23 nsew signal input
rlabel metal3 s 0 117512 800 117632 6 mem_addr[6]
port 24 nsew signal input
rlabel metal3 s 0 129752 800 129872 6 mem_addr[7]
port 25 nsew signal input
rlabel metal3 s 0 141992 800 142112 6 mem_addr[8]
port 26 nsew signal input
rlabel metal3 s 0 154232 800 154352 6 mem_addr[9]
port 27 nsew signal input
rlabel metal3 s 0 15512 800 15632 6 mem_cache_enable
port 28 nsew signal input
rlabel metal3 s 0 17552 800 17672 6 mem_exception
port 29 nsew signal output
rlabel metal3 s 0 37952 800 38072 6 mem_i_data[0]
port 30 nsew signal input
rlabel metal3 s 0 168512 800 168632 6 mem_i_data[10]
port 31 nsew signal input
rlabel metal3 s 0 180752 800 180872 6 mem_i_data[11]
port 32 nsew signal input
rlabel metal3 s 0 192992 800 193112 6 mem_i_data[12]
port 33 nsew signal input
rlabel metal3 s 0 205232 800 205352 6 mem_i_data[13]
port 34 nsew signal input
rlabel metal3 s 0 217472 800 217592 6 mem_i_data[14]
port 35 nsew signal input
rlabel metal3 s 0 229712 800 229832 6 mem_i_data[15]
port 36 nsew signal input
rlabel metal3 s 0 54272 800 54392 6 mem_i_data[1]
port 37 nsew signal input
rlabel metal3 s 0 70592 800 70712 6 mem_i_data[2]
port 38 nsew signal input
rlabel metal3 s 0 82832 800 82952 6 mem_i_data[3]
port 39 nsew signal input
rlabel metal3 s 0 95072 800 95192 6 mem_i_data[4]
port 40 nsew signal input
rlabel metal3 s 0 107312 800 107432 6 mem_i_data[5]
port 41 nsew signal input
rlabel metal3 s 0 119552 800 119672 6 mem_i_data[6]
port 42 nsew signal input
rlabel metal3 s 0 131792 800 131912 6 mem_i_data[7]
port 43 nsew signal input
rlabel metal3 s 0 144032 800 144152 6 mem_i_data[8]
port 44 nsew signal input
rlabel metal3 s 0 156272 800 156392 6 mem_i_data[9]
port 45 nsew signal input
rlabel metal3 s 0 39992 800 40112 6 mem_o_data[0]
port 46 nsew signal output
rlabel metal3 s 0 170552 800 170672 6 mem_o_data[10]
port 47 nsew signal output
rlabel metal3 s 0 182792 800 182912 6 mem_o_data[11]
port 48 nsew signal output
rlabel metal3 s 0 195032 800 195152 6 mem_o_data[12]
port 49 nsew signal output
rlabel metal3 s 0 207272 800 207392 6 mem_o_data[13]
port 50 nsew signal output
rlabel metal3 s 0 219512 800 219632 6 mem_o_data[14]
port 51 nsew signal output
rlabel metal3 s 0 231752 800 231872 6 mem_o_data[15]
port 52 nsew signal output
rlabel metal3 s 0 56312 800 56432 6 mem_o_data[1]
port 53 nsew signal output
rlabel metal3 s 0 72632 800 72752 6 mem_o_data[2]
port 54 nsew signal output
rlabel metal3 s 0 84872 800 84992 6 mem_o_data[3]
port 55 nsew signal output
rlabel metal3 s 0 97112 800 97232 6 mem_o_data[4]
port 56 nsew signal output
rlabel metal3 s 0 109352 800 109472 6 mem_o_data[5]
port 57 nsew signal output
rlabel metal3 s 0 121592 800 121712 6 mem_o_data[6]
port 58 nsew signal output
rlabel metal3 s 0 133832 800 133952 6 mem_o_data[7]
port 59 nsew signal output
rlabel metal3 s 0 146072 800 146192 6 mem_o_data[8]
port 60 nsew signal output
rlabel metal3 s 0 158312 800 158432 6 mem_o_data[9]
port 61 nsew signal output
rlabel metal3 s 0 19592 800 19712 6 mem_req
port 62 nsew signal input
rlabel metal3 s 0 42032 800 42152 6 mem_sel[0]
port 63 nsew signal input
rlabel metal3 s 0 58352 800 58472 6 mem_sel[1]
port 64 nsew signal input
rlabel metal3 s 0 21632 800 21752 6 mem_we
port 65 nsew signal input
rlabel metal4 s 4208 2128 4528 277488 6 vccd1
port 66 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 277488 6 vccd1
port 66 nsew power bidirectional
rlabel metal4 s 65648 2128 65968 277488 6 vccd1
port 66 nsew power bidirectional
rlabel metal4 s 96368 2128 96688 277488 6 vccd1
port 66 nsew power bidirectional
rlabel metal4 s 127088 2128 127408 277488 6 vccd1
port 66 nsew power bidirectional
rlabel metal4 s 157808 2128 158128 277488 6 vccd1
port 66 nsew power bidirectional
rlabel metal4 s 188528 2128 188848 277488 6 vccd1
port 66 nsew power bidirectional
rlabel metal4 s 219248 2128 219568 277488 6 vccd1
port 66 nsew power bidirectional
rlabel metal4 s 249968 2128 250288 277488 6 vccd1
port 66 nsew power bidirectional
rlabel metal4 s 280688 2128 281008 277488 6 vccd1
port 66 nsew power bidirectional
rlabel metal4 s 19568 2128 19888 277488 6 vssd1
port 67 nsew ground bidirectional
rlabel metal4 s 50288 2128 50608 277488 6 vssd1
port 67 nsew ground bidirectional
rlabel metal4 s 81008 2128 81328 277488 6 vssd1
port 67 nsew ground bidirectional
rlabel metal4 s 111728 2128 112048 277488 6 vssd1
port 67 nsew ground bidirectional
rlabel metal4 s 142448 2128 142768 277488 6 vssd1
port 67 nsew ground bidirectional
rlabel metal4 s 173168 2128 173488 277488 6 vssd1
port 67 nsew ground bidirectional
rlabel metal4 s 203888 2128 204208 277488 6 vssd1
port 67 nsew ground bidirectional
rlabel metal4 s 234608 2128 234928 277488 6 vssd1
port 67 nsew ground bidirectional
rlabel metal4 s 265328 2128 265648 277488 6 vssd1
port 67 nsew ground bidirectional
rlabel metal3 s 0 23672 800 23792 6 wb_4_burst
port 68 nsew signal output
rlabel metal3 s 0 25712 800 25832 6 wb_ack
port 69 nsew signal input
rlabel metal3 s 0 44072 800 44192 6 wb_adr[0]
port 70 nsew signal output
rlabel metal3 s 0 172592 800 172712 6 wb_adr[10]
port 71 nsew signal output
rlabel metal3 s 0 184832 800 184952 6 wb_adr[11]
port 72 nsew signal output
rlabel metal3 s 0 197072 800 197192 6 wb_adr[12]
port 73 nsew signal output
rlabel metal3 s 0 209312 800 209432 6 wb_adr[13]
port 74 nsew signal output
rlabel metal3 s 0 221552 800 221672 6 wb_adr[14]
port 75 nsew signal output
rlabel metal3 s 0 233792 800 233912 6 wb_adr[15]
port 76 nsew signal output
rlabel metal3 s 0 241952 800 242072 6 wb_adr[16]
port 77 nsew signal output
rlabel metal3 s 0 246032 800 246152 6 wb_adr[17]
port 78 nsew signal output
rlabel metal3 s 0 250112 800 250232 6 wb_adr[18]
port 79 nsew signal output
rlabel metal3 s 0 254192 800 254312 6 wb_adr[19]
port 80 nsew signal output
rlabel metal3 s 0 60392 800 60512 6 wb_adr[1]
port 81 nsew signal output
rlabel metal3 s 0 258272 800 258392 6 wb_adr[20]
port 82 nsew signal output
rlabel metal3 s 0 262352 800 262472 6 wb_adr[21]
port 83 nsew signal output
rlabel metal3 s 0 266432 800 266552 6 wb_adr[22]
port 84 nsew signal output
rlabel metal3 s 0 270512 800 270632 6 wb_adr[23]
port 85 nsew signal output
rlabel metal3 s 0 74672 800 74792 6 wb_adr[2]
port 86 nsew signal output
rlabel metal3 s 0 86912 800 87032 6 wb_adr[3]
port 87 nsew signal output
rlabel metal3 s 0 99152 800 99272 6 wb_adr[4]
port 88 nsew signal output
rlabel metal3 s 0 111392 800 111512 6 wb_adr[5]
port 89 nsew signal output
rlabel metal3 s 0 123632 800 123752 6 wb_adr[6]
port 90 nsew signal output
rlabel metal3 s 0 135872 800 135992 6 wb_adr[7]
port 91 nsew signal output
rlabel metal3 s 0 148112 800 148232 6 wb_adr[8]
port 92 nsew signal output
rlabel metal3 s 0 160352 800 160472 6 wb_adr[9]
port 93 nsew signal output
rlabel metal3 s 0 27752 800 27872 6 wb_cyc
port 94 nsew signal output
rlabel metal3 s 0 29792 800 29912 6 wb_err
port 95 nsew signal input
rlabel metal3 s 0 46112 800 46232 6 wb_i_dat[0]
port 96 nsew signal input
rlabel metal3 s 0 174632 800 174752 6 wb_i_dat[10]
port 97 nsew signal input
rlabel metal3 s 0 186872 800 186992 6 wb_i_dat[11]
port 98 nsew signal input
rlabel metal3 s 0 199112 800 199232 6 wb_i_dat[12]
port 99 nsew signal input
rlabel metal3 s 0 211352 800 211472 6 wb_i_dat[13]
port 100 nsew signal input
rlabel metal3 s 0 223592 800 223712 6 wb_i_dat[14]
port 101 nsew signal input
rlabel metal3 s 0 235832 800 235952 6 wb_i_dat[15]
port 102 nsew signal input
rlabel metal3 s 0 62432 800 62552 6 wb_i_dat[1]
port 103 nsew signal input
rlabel metal3 s 0 76712 800 76832 6 wb_i_dat[2]
port 104 nsew signal input
rlabel metal3 s 0 88952 800 89072 6 wb_i_dat[3]
port 105 nsew signal input
rlabel metal3 s 0 101192 800 101312 6 wb_i_dat[4]
port 106 nsew signal input
rlabel metal3 s 0 113432 800 113552 6 wb_i_dat[5]
port 107 nsew signal input
rlabel metal3 s 0 125672 800 125792 6 wb_i_dat[6]
port 108 nsew signal input
rlabel metal3 s 0 137912 800 138032 6 wb_i_dat[7]
port 109 nsew signal input
rlabel metal3 s 0 150152 800 150272 6 wb_i_dat[8]
port 110 nsew signal input
rlabel metal3 s 0 162392 800 162512 6 wb_i_dat[9]
port 111 nsew signal input
rlabel metal3 s 0 48152 800 48272 6 wb_o_dat[0]
port 112 nsew signal output
rlabel metal3 s 0 176672 800 176792 6 wb_o_dat[10]
port 113 nsew signal output
rlabel metal3 s 0 188912 800 189032 6 wb_o_dat[11]
port 114 nsew signal output
rlabel metal3 s 0 201152 800 201272 6 wb_o_dat[12]
port 115 nsew signal output
rlabel metal3 s 0 213392 800 213512 6 wb_o_dat[13]
port 116 nsew signal output
rlabel metal3 s 0 225632 800 225752 6 wb_o_dat[14]
port 117 nsew signal output
rlabel metal3 s 0 237872 800 237992 6 wb_o_dat[15]
port 118 nsew signal output
rlabel metal3 s 0 64472 800 64592 6 wb_o_dat[1]
port 119 nsew signal output
rlabel metal3 s 0 78752 800 78872 6 wb_o_dat[2]
port 120 nsew signal output
rlabel metal3 s 0 90992 800 91112 6 wb_o_dat[3]
port 121 nsew signal output
rlabel metal3 s 0 103232 800 103352 6 wb_o_dat[4]
port 122 nsew signal output
rlabel metal3 s 0 115472 800 115592 6 wb_o_dat[5]
port 123 nsew signal output
rlabel metal3 s 0 127712 800 127832 6 wb_o_dat[6]
port 124 nsew signal output
rlabel metal3 s 0 139952 800 140072 6 wb_o_dat[7]
port 125 nsew signal output
rlabel metal3 s 0 152192 800 152312 6 wb_o_dat[8]
port 126 nsew signal output
rlabel metal3 s 0 164432 800 164552 6 wb_o_dat[9]
port 127 nsew signal output
rlabel metal3 s 0 50192 800 50312 6 wb_sel[0]
port 128 nsew signal output
rlabel metal3 s 0 66512 800 66632 6 wb_sel[1]
port 129 nsew signal output
rlabel metal3 s 0 31832 800 31952 6 wb_stb
port 130 nsew signal output
rlabel metal3 s 0 33872 800 33992 6 wb_we
port 131 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 290000 280000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 225307784
string GDS_FILE /home/piotro/caravel_user_project/openlane/dcache/runs/22_12_29_19_29/results/signoff/dcache.magic.gds
string GDS_START 836450
<< end >>

