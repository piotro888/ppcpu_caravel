magic
tech sky130B
magscale 1 2
timestamp 1663071165
<< obsli1 >>
rect 1104 2159 158884 157777
<< obsm1 >>
rect 1104 2048 159054 157808
<< obsm2 >>
rect 1320 2042 159050 157797
<< metal3 >>
rect 0 157360 800 157480
rect 159200 155592 160000 155712
rect 0 153280 800 153400
rect 159200 152736 160000 152856
rect 159200 149880 160000 150000
rect 0 149200 800 149320
rect 159200 147024 160000 147144
rect 0 145120 800 145240
rect 159200 144168 160000 144288
rect 159200 141312 160000 141432
rect 0 141040 800 141160
rect 159200 138456 160000 138576
rect 0 136960 800 137080
rect 159200 135600 160000 135720
rect 0 132880 800 133000
rect 159200 132744 160000 132864
rect 159200 129888 160000 130008
rect 0 128800 800 128920
rect 159200 127032 160000 127152
rect 0 124720 800 124840
rect 159200 124176 160000 124296
rect 159200 121320 160000 121440
rect 0 120640 800 120760
rect 159200 118464 160000 118584
rect 0 116560 800 116680
rect 159200 115608 160000 115728
rect 159200 112752 160000 112872
rect 0 112480 800 112600
rect 159200 109896 160000 110016
rect 0 108400 800 108520
rect 159200 107040 160000 107160
rect 0 104320 800 104440
rect 159200 104184 160000 104304
rect 159200 101328 160000 101448
rect 0 100240 800 100360
rect 159200 98472 160000 98592
rect 0 96160 800 96280
rect 159200 95616 160000 95736
rect 159200 92760 160000 92880
rect 0 92080 800 92200
rect 159200 89904 160000 90024
rect 0 88000 800 88120
rect 159200 87048 160000 87168
rect 159200 84192 160000 84312
rect 0 83920 800 84040
rect 159200 81336 160000 81456
rect 0 79840 800 79960
rect 159200 78480 160000 78600
rect 0 75760 800 75880
rect 159200 75624 160000 75744
rect 159200 72768 160000 72888
rect 0 71680 800 71800
rect 159200 69912 160000 70032
rect 0 67600 800 67720
rect 159200 67056 160000 67176
rect 159200 64200 160000 64320
rect 0 63520 800 63640
rect 159200 61344 160000 61464
rect 0 59440 800 59560
rect 159200 58488 160000 58608
rect 159200 55632 160000 55752
rect 0 55360 800 55480
rect 159200 52776 160000 52896
rect 0 51280 800 51400
rect 159200 49920 160000 50040
rect 0 47200 800 47320
rect 159200 47064 160000 47184
rect 159200 44208 160000 44328
rect 0 43120 800 43240
rect 159200 41352 160000 41472
rect 0 39040 800 39160
rect 159200 38496 160000 38616
rect 159200 35640 160000 35760
rect 0 34960 800 35080
rect 159200 32784 160000 32904
rect 0 30880 800 31000
rect 159200 29928 160000 30048
rect 159200 27072 160000 27192
rect 0 26800 800 26920
rect 159200 24216 160000 24336
rect 0 22720 800 22840
rect 159200 21360 160000 21480
rect 0 18640 800 18760
rect 159200 18504 160000 18624
rect 159200 15648 160000 15768
rect 0 14560 800 14680
rect 159200 12792 160000 12912
rect 0 10480 800 10600
rect 159200 9936 160000 10056
rect 159200 7080 160000 7200
rect 0 6400 800 6520
rect 159200 4224 160000 4344
rect 0 2320 800 2440
<< obsm3 >>
rect 800 157560 159282 157793
rect 880 157280 159282 157560
rect 800 155792 159282 157280
rect 800 155512 159120 155792
rect 800 153480 159282 155512
rect 880 153200 159282 153480
rect 800 152936 159282 153200
rect 800 152656 159120 152936
rect 800 150080 159282 152656
rect 800 149800 159120 150080
rect 800 149400 159282 149800
rect 880 149120 159282 149400
rect 800 147224 159282 149120
rect 800 146944 159120 147224
rect 800 145320 159282 146944
rect 880 145040 159282 145320
rect 800 144368 159282 145040
rect 800 144088 159120 144368
rect 800 141512 159282 144088
rect 800 141240 159120 141512
rect 880 141232 159120 141240
rect 880 140960 159282 141232
rect 800 138656 159282 140960
rect 800 138376 159120 138656
rect 800 137160 159282 138376
rect 880 136880 159282 137160
rect 800 135800 159282 136880
rect 800 135520 159120 135800
rect 800 133080 159282 135520
rect 880 132944 159282 133080
rect 880 132800 159120 132944
rect 800 132664 159120 132800
rect 800 130088 159282 132664
rect 800 129808 159120 130088
rect 800 129000 159282 129808
rect 880 128720 159282 129000
rect 800 127232 159282 128720
rect 800 126952 159120 127232
rect 800 124920 159282 126952
rect 880 124640 159282 124920
rect 800 124376 159282 124640
rect 800 124096 159120 124376
rect 800 121520 159282 124096
rect 800 121240 159120 121520
rect 800 120840 159282 121240
rect 880 120560 159282 120840
rect 800 118664 159282 120560
rect 800 118384 159120 118664
rect 800 116760 159282 118384
rect 880 116480 159282 116760
rect 800 115808 159282 116480
rect 800 115528 159120 115808
rect 800 112952 159282 115528
rect 800 112680 159120 112952
rect 880 112672 159120 112680
rect 880 112400 159282 112672
rect 800 110096 159282 112400
rect 800 109816 159120 110096
rect 800 108600 159282 109816
rect 880 108320 159282 108600
rect 800 107240 159282 108320
rect 800 106960 159120 107240
rect 800 104520 159282 106960
rect 880 104384 159282 104520
rect 880 104240 159120 104384
rect 800 104104 159120 104240
rect 800 101528 159282 104104
rect 800 101248 159120 101528
rect 800 100440 159282 101248
rect 880 100160 159282 100440
rect 800 98672 159282 100160
rect 800 98392 159120 98672
rect 800 96360 159282 98392
rect 880 96080 159282 96360
rect 800 95816 159282 96080
rect 800 95536 159120 95816
rect 800 92960 159282 95536
rect 800 92680 159120 92960
rect 800 92280 159282 92680
rect 880 92000 159282 92280
rect 800 90104 159282 92000
rect 800 89824 159120 90104
rect 800 88200 159282 89824
rect 880 87920 159282 88200
rect 800 87248 159282 87920
rect 800 86968 159120 87248
rect 800 84392 159282 86968
rect 800 84120 159120 84392
rect 880 84112 159120 84120
rect 880 83840 159282 84112
rect 800 81536 159282 83840
rect 800 81256 159120 81536
rect 800 80040 159282 81256
rect 880 79760 159282 80040
rect 800 78680 159282 79760
rect 800 78400 159120 78680
rect 800 75960 159282 78400
rect 880 75824 159282 75960
rect 880 75680 159120 75824
rect 800 75544 159120 75680
rect 800 72968 159282 75544
rect 800 72688 159120 72968
rect 800 71880 159282 72688
rect 880 71600 159282 71880
rect 800 70112 159282 71600
rect 800 69832 159120 70112
rect 800 67800 159282 69832
rect 880 67520 159282 67800
rect 800 67256 159282 67520
rect 800 66976 159120 67256
rect 800 64400 159282 66976
rect 800 64120 159120 64400
rect 800 63720 159282 64120
rect 880 63440 159282 63720
rect 800 61544 159282 63440
rect 800 61264 159120 61544
rect 800 59640 159282 61264
rect 880 59360 159282 59640
rect 800 58688 159282 59360
rect 800 58408 159120 58688
rect 800 55832 159282 58408
rect 800 55560 159120 55832
rect 880 55552 159120 55560
rect 880 55280 159282 55552
rect 800 52976 159282 55280
rect 800 52696 159120 52976
rect 800 51480 159282 52696
rect 880 51200 159282 51480
rect 800 50120 159282 51200
rect 800 49840 159120 50120
rect 800 47400 159282 49840
rect 880 47264 159282 47400
rect 880 47120 159120 47264
rect 800 46984 159120 47120
rect 800 44408 159282 46984
rect 800 44128 159120 44408
rect 800 43320 159282 44128
rect 880 43040 159282 43320
rect 800 41552 159282 43040
rect 800 41272 159120 41552
rect 800 39240 159282 41272
rect 880 38960 159282 39240
rect 800 38696 159282 38960
rect 800 38416 159120 38696
rect 800 35840 159282 38416
rect 800 35560 159120 35840
rect 800 35160 159282 35560
rect 880 34880 159282 35160
rect 800 32984 159282 34880
rect 800 32704 159120 32984
rect 800 31080 159282 32704
rect 880 30800 159282 31080
rect 800 30128 159282 30800
rect 800 29848 159120 30128
rect 800 27272 159282 29848
rect 800 27000 159120 27272
rect 880 26992 159120 27000
rect 880 26720 159282 26992
rect 800 24416 159282 26720
rect 800 24136 159120 24416
rect 800 22920 159282 24136
rect 880 22640 159282 22920
rect 800 21560 159282 22640
rect 800 21280 159120 21560
rect 800 18840 159282 21280
rect 880 18704 159282 18840
rect 880 18560 159120 18704
rect 800 18424 159120 18560
rect 800 15848 159282 18424
rect 800 15568 159120 15848
rect 800 14760 159282 15568
rect 880 14480 159282 14760
rect 800 12992 159282 14480
rect 800 12712 159120 12992
rect 800 10680 159282 12712
rect 880 10400 159282 10680
rect 800 10136 159282 10400
rect 800 9856 159120 10136
rect 800 7280 159282 9856
rect 800 7000 159120 7280
rect 800 6600 159282 7000
rect 880 6320 159282 6600
rect 800 4424 159282 6320
rect 800 4144 159120 4424
rect 800 2520 159282 4144
rect 880 2240 159282 2520
rect 800 2143 159282 2240
<< metal4 >>
rect 4208 2128 4528 157808
rect 19568 2128 19888 157808
rect 34928 2128 35248 157808
rect 50288 2128 50608 157808
rect 65648 2128 65968 157808
rect 81008 2128 81328 157808
rect 96368 2128 96688 157808
rect 111728 2128 112048 157808
rect 127088 2128 127408 157808
rect 142448 2128 142768 157808
rect 157808 2128 158128 157808
<< obsm4 >>
rect 1899 2347 4128 154597
rect 4608 2347 19488 154597
rect 19968 2347 34848 154597
rect 35328 2347 50208 154597
rect 50688 2347 65568 154597
rect 66048 2347 80928 154597
rect 81408 2347 96288 154597
rect 96768 2347 111648 154597
rect 112128 2347 127008 154597
rect 127488 2347 142368 154597
rect 142848 2347 157261 154597
<< labels >>
rlabel metal3 s 159200 152736 160000 152856 6 i_clk
port 1 nsew signal input
rlabel metal3 s 159200 155592 160000 155712 6 i_rst
port 2 nsew signal input
rlabel metal3 s 159200 4224 160000 4344 6 mem_ack
port 3 nsew signal output
rlabel metal3 s 159200 7080 160000 7200 6 mem_addr[0]
port 4 nsew signal input
rlabel metal3 s 159200 35640 160000 35760 6 mem_addr[10]
port 5 nsew signal input
rlabel metal3 s 159200 38496 160000 38616 6 mem_addr[11]
port 6 nsew signal input
rlabel metal3 s 159200 41352 160000 41472 6 mem_addr[12]
port 7 nsew signal input
rlabel metal3 s 159200 44208 160000 44328 6 mem_addr[13]
port 8 nsew signal input
rlabel metal3 s 159200 47064 160000 47184 6 mem_addr[14]
port 9 nsew signal input
rlabel metal3 s 159200 49920 160000 50040 6 mem_addr[15]
port 10 nsew signal input
rlabel metal3 s 159200 9936 160000 10056 6 mem_addr[1]
port 11 nsew signal input
rlabel metal3 s 159200 12792 160000 12912 6 mem_addr[2]
port 12 nsew signal input
rlabel metal3 s 159200 15648 160000 15768 6 mem_addr[3]
port 13 nsew signal input
rlabel metal3 s 159200 18504 160000 18624 6 mem_addr[4]
port 14 nsew signal input
rlabel metal3 s 159200 21360 160000 21480 6 mem_addr[5]
port 15 nsew signal input
rlabel metal3 s 159200 24216 160000 24336 6 mem_addr[6]
port 16 nsew signal input
rlabel metal3 s 159200 27072 160000 27192 6 mem_addr[7]
port 17 nsew signal input
rlabel metal3 s 159200 29928 160000 30048 6 mem_addr[8]
port 18 nsew signal input
rlabel metal3 s 159200 32784 160000 32904 6 mem_addr[9]
port 19 nsew signal input
rlabel metal3 s 159200 52776 160000 52896 6 mem_cache_flush
port 20 nsew signal input
rlabel metal3 s 159200 55632 160000 55752 6 mem_data[0]
port 21 nsew signal output
rlabel metal3 s 159200 84192 160000 84312 6 mem_data[10]
port 22 nsew signal output
rlabel metal3 s 159200 87048 160000 87168 6 mem_data[11]
port 23 nsew signal output
rlabel metal3 s 159200 89904 160000 90024 6 mem_data[12]
port 24 nsew signal output
rlabel metal3 s 159200 92760 160000 92880 6 mem_data[13]
port 25 nsew signal output
rlabel metal3 s 159200 95616 160000 95736 6 mem_data[14]
port 26 nsew signal output
rlabel metal3 s 159200 98472 160000 98592 6 mem_data[15]
port 27 nsew signal output
rlabel metal3 s 159200 101328 160000 101448 6 mem_data[16]
port 28 nsew signal output
rlabel metal3 s 159200 104184 160000 104304 6 mem_data[17]
port 29 nsew signal output
rlabel metal3 s 159200 107040 160000 107160 6 mem_data[18]
port 30 nsew signal output
rlabel metal3 s 159200 109896 160000 110016 6 mem_data[19]
port 31 nsew signal output
rlabel metal3 s 159200 58488 160000 58608 6 mem_data[1]
port 32 nsew signal output
rlabel metal3 s 159200 112752 160000 112872 6 mem_data[20]
port 33 nsew signal output
rlabel metal3 s 159200 115608 160000 115728 6 mem_data[21]
port 34 nsew signal output
rlabel metal3 s 159200 118464 160000 118584 6 mem_data[22]
port 35 nsew signal output
rlabel metal3 s 159200 121320 160000 121440 6 mem_data[23]
port 36 nsew signal output
rlabel metal3 s 159200 124176 160000 124296 6 mem_data[24]
port 37 nsew signal output
rlabel metal3 s 159200 127032 160000 127152 6 mem_data[25]
port 38 nsew signal output
rlabel metal3 s 159200 129888 160000 130008 6 mem_data[26]
port 39 nsew signal output
rlabel metal3 s 159200 132744 160000 132864 6 mem_data[27]
port 40 nsew signal output
rlabel metal3 s 159200 135600 160000 135720 6 mem_data[28]
port 41 nsew signal output
rlabel metal3 s 159200 138456 160000 138576 6 mem_data[29]
port 42 nsew signal output
rlabel metal3 s 159200 61344 160000 61464 6 mem_data[2]
port 43 nsew signal output
rlabel metal3 s 159200 141312 160000 141432 6 mem_data[30]
port 44 nsew signal output
rlabel metal3 s 159200 144168 160000 144288 6 mem_data[31]
port 45 nsew signal output
rlabel metal3 s 159200 64200 160000 64320 6 mem_data[3]
port 46 nsew signal output
rlabel metal3 s 159200 67056 160000 67176 6 mem_data[4]
port 47 nsew signal output
rlabel metal3 s 159200 69912 160000 70032 6 mem_data[5]
port 48 nsew signal output
rlabel metal3 s 159200 72768 160000 72888 6 mem_data[6]
port 49 nsew signal output
rlabel metal3 s 159200 75624 160000 75744 6 mem_data[7]
port 50 nsew signal output
rlabel metal3 s 159200 78480 160000 78600 6 mem_data[8]
port 51 nsew signal output
rlabel metal3 s 159200 81336 160000 81456 6 mem_data[9]
port 52 nsew signal output
rlabel metal3 s 159200 147024 160000 147144 6 mem_ppl_submit
port 53 nsew signal input
rlabel metal3 s 159200 149880 160000 150000 6 mem_req
port 54 nsew signal input
rlabel metal4 s 4208 2128 4528 157808 6 vccd1
port 55 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 157808 6 vccd1
port 55 nsew power bidirectional
rlabel metal4 s 65648 2128 65968 157808 6 vccd1
port 55 nsew power bidirectional
rlabel metal4 s 96368 2128 96688 157808 6 vccd1
port 55 nsew power bidirectional
rlabel metal4 s 127088 2128 127408 157808 6 vccd1
port 55 nsew power bidirectional
rlabel metal4 s 157808 2128 158128 157808 6 vccd1
port 55 nsew power bidirectional
rlabel metal4 s 19568 2128 19888 157808 6 vssd1
port 56 nsew ground bidirectional
rlabel metal4 s 50288 2128 50608 157808 6 vssd1
port 56 nsew ground bidirectional
rlabel metal4 s 81008 2128 81328 157808 6 vssd1
port 56 nsew ground bidirectional
rlabel metal4 s 111728 2128 112048 157808 6 vssd1
port 56 nsew ground bidirectional
rlabel metal4 s 142448 2128 142768 157808 6 vssd1
port 56 nsew ground bidirectional
rlabel metal3 s 0 2320 800 2440 6 wb_ack
port 57 nsew signal input
rlabel metal3 s 0 6400 800 6520 6 wb_adr[0]
port 58 nsew signal output
rlabel metal3 s 0 47200 800 47320 6 wb_adr[10]
port 59 nsew signal output
rlabel metal3 s 0 51280 800 51400 6 wb_adr[11]
port 60 nsew signal output
rlabel metal3 s 0 55360 800 55480 6 wb_adr[12]
port 61 nsew signal output
rlabel metal3 s 0 59440 800 59560 6 wb_adr[13]
port 62 nsew signal output
rlabel metal3 s 0 63520 800 63640 6 wb_adr[14]
port 63 nsew signal output
rlabel metal3 s 0 67600 800 67720 6 wb_adr[15]
port 64 nsew signal output
rlabel metal3 s 0 10480 800 10600 6 wb_adr[1]
port 65 nsew signal output
rlabel metal3 s 0 14560 800 14680 6 wb_adr[2]
port 66 nsew signal output
rlabel metal3 s 0 18640 800 18760 6 wb_adr[3]
port 67 nsew signal output
rlabel metal3 s 0 22720 800 22840 6 wb_adr[4]
port 68 nsew signal output
rlabel metal3 s 0 26800 800 26920 6 wb_adr[5]
port 69 nsew signal output
rlabel metal3 s 0 30880 800 31000 6 wb_adr[6]
port 70 nsew signal output
rlabel metal3 s 0 34960 800 35080 6 wb_adr[7]
port 71 nsew signal output
rlabel metal3 s 0 39040 800 39160 6 wb_adr[8]
port 72 nsew signal output
rlabel metal3 s 0 43120 800 43240 6 wb_adr[9]
port 73 nsew signal output
rlabel metal3 s 0 71680 800 71800 6 wb_cyc
port 74 nsew signal output
rlabel metal3 s 0 75760 800 75880 6 wb_err
port 75 nsew signal input
rlabel metal3 s 0 79840 800 79960 6 wb_i_dat[0]
port 76 nsew signal input
rlabel metal3 s 0 120640 800 120760 6 wb_i_dat[10]
port 77 nsew signal input
rlabel metal3 s 0 124720 800 124840 6 wb_i_dat[11]
port 78 nsew signal input
rlabel metal3 s 0 128800 800 128920 6 wb_i_dat[12]
port 79 nsew signal input
rlabel metal3 s 0 132880 800 133000 6 wb_i_dat[13]
port 80 nsew signal input
rlabel metal3 s 0 136960 800 137080 6 wb_i_dat[14]
port 81 nsew signal input
rlabel metal3 s 0 141040 800 141160 6 wb_i_dat[15]
port 82 nsew signal input
rlabel metal3 s 0 83920 800 84040 6 wb_i_dat[1]
port 83 nsew signal input
rlabel metal3 s 0 88000 800 88120 6 wb_i_dat[2]
port 84 nsew signal input
rlabel metal3 s 0 92080 800 92200 6 wb_i_dat[3]
port 85 nsew signal input
rlabel metal3 s 0 96160 800 96280 6 wb_i_dat[4]
port 86 nsew signal input
rlabel metal3 s 0 100240 800 100360 6 wb_i_dat[5]
port 87 nsew signal input
rlabel metal3 s 0 104320 800 104440 6 wb_i_dat[6]
port 88 nsew signal input
rlabel metal3 s 0 108400 800 108520 6 wb_i_dat[7]
port 89 nsew signal input
rlabel metal3 s 0 112480 800 112600 6 wb_i_dat[8]
port 90 nsew signal input
rlabel metal3 s 0 116560 800 116680 6 wb_i_dat[9]
port 91 nsew signal input
rlabel metal3 s 0 145120 800 145240 6 wb_sel[0]
port 92 nsew signal output
rlabel metal3 s 0 149200 800 149320 6 wb_sel[1]
port 93 nsew signal output
rlabel metal3 s 0 153280 800 153400 6 wb_stb
port 94 nsew signal output
rlabel metal3 s 0 157360 800 157480 6 wb_we
port 95 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 160000 160000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 76045352
string GDS_FILE /home/piotro/ppcpu_caravel/openlane/icache/runs/22_09_13_13_55/results/signoff/icache.magic.gds
string GDS_START 604212
<< end >>

