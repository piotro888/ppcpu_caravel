* NGSPICE file created from core0.ext - technology: gf180mcuD

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__antenna abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__antenna I VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__filltie abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__filltie VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fill_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fill_2 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fill_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fill_1 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dffq_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dffq_1 D CLK Q VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi21_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi21_1 A1 A2 B ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_8 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_8 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_16 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_16 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_4 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand3_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand3_2 A1 A2 A3 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai21_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai21_1 A1 A2 B ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor2_1 A1 A2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_64 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_64 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__inv_3 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__inv_3 I ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_32 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_32 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand2_2 A1 A2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand2_1 A1 A2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_1 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi22_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi22_1 A1 A2 B1 B2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and2_1 A1 A2 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dffq_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dffq_4 D CLK Q VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dffq_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dffq_2 D CLK Q VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_2 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai211_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai211_2 A1 A2 B C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__endcap abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__endcap VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand3_1 A1 A2 A3 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor3_1 A1 A2 A3 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__mux2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__mux2_2 I0 I1 S Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor2_2 A1 A2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai211_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai211_4 A1 A2 B C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkinv_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkinv_1 I ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand4_1 A1 A2 A3 A4 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_4 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai21_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai21_2 A1 A2 B ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai221_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai221_4 A1 A2 B1 B2 C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi21_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi21_2 A1 A2 B ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor2_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor2_4 A1 A2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi211_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi211_1 A1 A2 B C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi221_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi221_4 A1 A2 B1 B2 C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai211_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai211_1 A1 A2 B C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor4_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor4_4 A1 A2 A3 A4 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xor2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xor2_1 A1 A2 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi21_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi21_4 A1 A2 B ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi211_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi211_4 A1 A2 B C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_3 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_3 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and3_1 A1 A2 A3 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand2_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand2_4 A1 A2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or2_1 A1 A2 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dlya_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dlya_2 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor3_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor3_4 A1 A2 A3 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand4_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand4_2 A1 A2 A3 A4 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__inv_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__inv_1 I ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai21_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai21_4 A1 A2 B ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand4_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand4_4 A1 A2 A3 A4 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai22_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai22_1 A1 A2 B1 B2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or4_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or4_2 A1 A2 A3 A4 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai32_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai32_2 A1 A2 A3 B1 B2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai31_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai31_4 A1 A2 A3 B ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor3_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor3_2 A1 A2 A3 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xnor2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xnor2_1 A1 A2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi22_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi22_2 A1 A2 B1 B2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xor2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xor2_2 A1 A2 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and2_2 A1 A2 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or3_1 A1 A2 A3 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai222_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai222_1 A1 A2 B1 B2 C1 C2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi221_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi221_2 A1 A2 B1 B2 C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi222_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi222_4 A1 A2 B1 B2 C1 C2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkinv_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkinv_2 I ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xor3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xor3_1 A1 A2 A3 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or3_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or3_2 A1 A2 A3 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and3_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and3_2 A1 A2 A3 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi222_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi222_1 A1 A2 B1 B2 C1 C2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi211_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi211_2 A1 A2 B C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or4_1 A1 A2 A3 A4 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi221_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi221_1 A1 A2 B1 B2 C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand3_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand3_4 A1 A2 A3 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_8 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_8 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or2_2 A1 A2 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai31_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai31_2 A1 A2 A3 B ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai221_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai221_1 A1 A2 B1 B2 C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__mux2_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__mux2_4 I0 I1 S Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi22_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi22_4 A1 A2 B1 B2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai22_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai22_4 A1 A2 B1 B2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai32_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai32_1 A1 A2 A3 B1 B2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkinv_3 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkinv_3 I ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkinv_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkinv_4 I ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__inv_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__inv_4 I ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__inv_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__inv_2 I ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi222_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi222_2 A1 A2 B1 B2 C1 C2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and4_1 A1 A2 A3 A4 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and4_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and4_2 A1 A2 A3 A4 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__mux4_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__mux4_4 I0 I1 I2 I3 S0 S1 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or2_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or2_4 A1 A2 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai221_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai221_2 A1 A2 B1 B2 C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and2_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and2_4 A1 A2 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xor3_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xor3_2 A1 A2 A3 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or4_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or4_4 A1 A2 A3 A4 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor4_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor4_2 A1 A2 A3 A4 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai22_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai22_2 A1 A2 B1 B2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__tiel abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__tiel ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai31_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai31_1 A1 A2 A3 B ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__mux4_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__mux4_2 I0 I1 I2 I3 S0 S1 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and3_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and3_4 A1 A2 A3 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xor2_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xor2_4 A1 A2 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__mux4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__mux4_1 I0 I1 I2 I3 S0 S1 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dlyc_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dlyc_4 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai222_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai222_4 A1 A2 B1 B2 C1 C2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or3_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or3_4 A1 A2 A3 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai32_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai32_4 A1 A2 A3 B1 B2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkinv_8 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkinv_8 I ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xnor3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xnor3_1 A1 A2 A3 ZN VDD VNW VPW VSS
.ends

.subckt core0 dbg_pc[0] dbg_pc[10] dbg_pc[11] dbg_pc[12] dbg_pc[13] dbg_pc[14] dbg_pc[15]
+ dbg_pc[1] dbg_pc[2] dbg_pc[3] dbg_pc[4] dbg_pc[5] dbg_pc[6] dbg_pc[7] dbg_pc[8]
+ dbg_pc[9] dbg_r0[0] dbg_r0[10] dbg_r0[11] dbg_r0[12] dbg_r0[13] dbg_r0[14] dbg_r0[15]
+ dbg_r0[1] dbg_r0[2] dbg_r0[3] dbg_r0[4] dbg_r0[5] dbg_r0[6] dbg_r0[7] dbg_r0[8]
+ dbg_r0[9] i_clk i_core_int_sreg[0] i_core_int_sreg[10] i_core_int_sreg[11] i_core_int_sreg[12]
+ i_core_int_sreg[13] i_core_int_sreg[14] i_core_int_sreg[15] i_core_int_sreg[1] i_core_int_sreg[2]
+ i_core_int_sreg[3] i_core_int_sreg[4] i_core_int_sreg[5] i_core_int_sreg[6] i_core_int_sreg[7]
+ i_core_int_sreg[8] i_core_int_sreg[9] i_disable i_irq i_mc_core_int i_mem_ack i_mem_data[0]
+ i_mem_data[10] i_mem_data[11] i_mem_data[12] i_mem_data[13] i_mem_data[14] i_mem_data[15]
+ i_mem_data[1] i_mem_data[2] i_mem_data[3] i_mem_data[4] i_mem_data[5] i_mem_data[6]
+ i_mem_data[7] i_mem_data[8] i_mem_data[9] i_mem_exception i_req_data[0] i_req_data[10]
+ i_req_data[11] i_req_data[12] i_req_data[13] i_req_data[14] i_req_data[15] i_req_data[16]
+ i_req_data[17] i_req_data[18] i_req_data[19] i_req_data[1] i_req_data[20] i_req_data[21]
+ i_req_data[22] i_req_data[23] i_req_data[24] i_req_data[25] i_req_data[26] i_req_data[27]
+ i_req_data[28] i_req_data[29] i_req_data[2] i_req_data[30] i_req_data[31] i_req_data[3]
+ i_req_data[4] i_req_data[5] i_req_data[6] i_req_data[7] i_req_data[8] i_req_data[9]
+ i_req_data_valid i_rst o_c_data_page o_c_instr_long o_c_instr_page o_icache_flush
+ o_instr_long_addr[0] o_instr_long_addr[1] o_instr_long_addr[2] o_instr_long_addr[3]
+ o_instr_long_addr[4] o_instr_long_addr[5] o_instr_long_addr[6] o_instr_long_addr[7]
+ o_mem_addr[0] o_mem_addr[10] o_mem_addr[11] o_mem_addr[12] o_mem_addr[13] o_mem_addr[14]
+ o_mem_addr[15] o_mem_addr[1] o_mem_addr[2] o_mem_addr[3] o_mem_addr[4] o_mem_addr[5]
+ o_mem_addr[6] o_mem_addr[7] o_mem_addr[8] o_mem_addr[9] o_mem_addr_high[0] o_mem_addr_high[1]
+ o_mem_addr_high[2] o_mem_addr_high[3] o_mem_addr_high[4] o_mem_addr_high[5] o_mem_addr_high[6]
+ o_mem_data[0] o_mem_data[10] o_mem_data[11] o_mem_data[12] o_mem_data[13] o_mem_data[14]
+ o_mem_data[15] o_mem_data[1] o_mem_data[2] o_mem_data[3] o_mem_data[4] o_mem_data[5]
+ o_mem_data[6] o_mem_data[7] o_mem_data[8] o_mem_data[9] o_mem_long o_mem_req o_mem_sel[0]
+ o_mem_sel[1] o_mem_we o_req_active o_req_addr[0] o_req_addr[10] o_req_addr[11] o_req_addr[12]
+ o_req_addr[13] o_req_addr[14] o_req_addr[15] o_req_addr[1] o_req_addr[2] o_req_addr[3]
+ o_req_addr[4] o_req_addr[5] o_req_addr[6] o_req_addr[7] o_req_addr[8] o_req_addr[9]
+ o_req_ppl_submit sr_bus_addr[0] sr_bus_addr[10] sr_bus_addr[11] sr_bus_addr[12]
+ sr_bus_addr[13] sr_bus_addr[14] sr_bus_addr[15] sr_bus_addr[1] sr_bus_addr[2] sr_bus_addr[3]
+ sr_bus_addr[4] sr_bus_addr[5] sr_bus_addr[6] sr_bus_addr[7] sr_bus_addr[8] sr_bus_addr[9]
+ sr_bus_data_o[0] sr_bus_data_o[10] sr_bus_data_o[11] sr_bus_data_o[12] sr_bus_data_o[13]
+ sr_bus_data_o[14] sr_bus_data_o[15] sr_bus_data_o[1] sr_bus_data_o[2] sr_bus_data_o[3]
+ sr_bus_data_o[4] sr_bus_data_o[5] sr_bus_data_o[6] sr_bus_data_o[7] sr_bus_data_o[8]
+ sr_bus_data_o[9] sr_bus_we vccd1 vssd1 o_mem_addr_high[7]
XANTENNA__6209__A2 _2409_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7406__A1 _1357_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_2_538 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_222_732 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_118_95 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7963_ _0141_ clknet_leaf_22_i_clk net104 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_38_968 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6914_ _2983_ _3129_ _3142_ _0342_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_7894_ _0085_ clknet_leaf_71_i_clk core_0.decode.i_imm_pass\[3\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_221_286 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4373__C _0963_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4640__A1 net181 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7709__A2 _1098_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_347 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_159_2418 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_76_144 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6845_ _2990_ _3087_ _3102_ _0313_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_147_522 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_175_831 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_175_842 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_64_317 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_147_555 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_734 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5196__A2 _1435_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_91_125 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6776_ _2996_ _3043_ _3062_ _0284_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_3988_ _0533_ core_0.execute.rf.reg_outputs\[4\]\[9\] net230 _0618_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_0_9_477 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_91_136 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_419 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_147_588 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5485__B _1367_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_91_158 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5727_ _2126_ _2127_ _1689_ _2128_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_73_862 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_134_227 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_17_255 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_115_430 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6145__A1 core_0.execute.pc_high_out\[6\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_5_650 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_60_523 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5658_ _1754_ _1585_ _2059_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_143_772 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_32_247 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_130_400 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_211_3040 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_102_102 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_103_625 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_32_258 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_5_694 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6696__A2 _3006_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4609_ _1169_ _1170_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__inv_3
XFILLER_0_20_409 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_170_591 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5589_ _1988_ _1989_ _1990_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__5705__S _1819_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7328_ _2384_ _2434_ _3501_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_102_157 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_130_477 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7645__A1 _3732_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6448__A2 _1386_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7259_ net85 _3426_ net86 _3440_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_183_2703 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_244_301 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4459__A1 core_0.decode.oc_alu_mode\[1\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_183_2714 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_110_190 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_217_559 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5120__A2 _1486_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6536__S _2906_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5671__A3 _1994_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_225_570 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5959__A1 core_0.execute.sreg_scratch.o_d\[2\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_222_3180 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_68_601 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5959__B2 net9 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_212_242 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_169_135 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_169_146 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_240_573 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_197_466 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_169_157 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_197_488 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_185_628 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_807 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_68_667 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_509 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_155 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_678 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_103_1749 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_140_2190 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_184_138 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_166_853 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_194_2843 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_82_103 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7594__C _3672_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6384__A1 _1501_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_83_648 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_193_683 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_391 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_125_205 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_126_728 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_82_147 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5395__B _1817_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_192_171 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_82_158 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4934__A2 _1394_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_715 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_24_737 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xrebuffer7 net228 net229 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_106_452 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_134_761 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_180_366 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_236 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_58_1206 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6687__A2 _3006_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_121_422 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_133_282 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6938__C _1225_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_236_802 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_37 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_114_1878 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7636__A1 core_0.execute.pc_high_buff_out\[4\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_225_3209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_120_i_clk clknet_4_3__leaf_i_clk clknet_leaf_120_i_clk vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_235_378 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_69_1335 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_188_422 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_69_1346 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_207_2997 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6998__I0 _2001_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_231_562 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_58_100 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6611__A2 _2956_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4960_ core_0.execute.sreg_priv_control.o_d\[9\] _1394_ _1415_ _1391_ _1416_ vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_TAPCELL_ROW_35_927 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_82_1502 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_35_938 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_3911_ core_0.dec_r_reg_sel\[1\] _0518_ _0547_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_58_155 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3976__A3 _0520_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_157_842 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4891_ _0726_ _1146_ _1359_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_58_166 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_317 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_104_31 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_236_3349 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6630_ _2936_ _2972_ _2973_ _0227_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__6375__A1 net74 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5178__A2 _1615_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_129_566 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_156_352 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_659 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6375__B2 _2537_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_542 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_171_300 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_15_695 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_73_158 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6561_ _2921_ _0210_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_144_547 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_27_586 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_54_372 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8300_ _0476_ clknet_leaf_16_i_clk net185 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_4
X_5512_ _1841_ _1719_ _1944_ _0138_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_154_2359 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6492_ core_0.ew_data\[14\] _2486_ _2871_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_120_30 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_125_772 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_131_208 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_247 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_70_865 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8231_ _0407_ clknet_leaf_13_i_clk core_0.execute.sreg_irq_pc.o_d\[3\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_30_718 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6678__A2 _2999_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5443_ _1374_ _1880_ _1881_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_140_731 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_152_591 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_93_1631 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_8162_ _0338_ clknet_leaf_89_i_clk net99 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_4
XFILLER_0_196_34 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_10_420 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_100_617 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5374_ _1809_ _1822_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_140_797 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7627__A1 net221 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7113_ _1226_ _1491_ _3321_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4325_ _0725_ _0817_ _0943_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_8093_ _0269_ clknet_leaf_92_i_clk core_0.execute.rf.reg_outputs\[4\]\[0\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_226_312 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7044_ _1592_ _3209_ _3257_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_129_72 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4256_ _0726_ _0727_ _0813_ _0874_ _0875_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai211_2
XANTENNA__5102__A2 net178 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4187_ core_0.ew_mem_access core_0.ew_submit _0806_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_165_2488 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_241_337 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_167_606 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_179_466 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7946_ _0124_ clknet_leaf_5_i_clk core_0.execute.alu_mul_div.div_cur\[2\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_49_122 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_49_133 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_194_425 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_38_807 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__3967__A3 net231 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7877_ _0068_ clknet_leaf_47_i_clk core_0.decode.i_instr_l\[2\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_4
XFILLER_0_65_615 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_92_401 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_148_864 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_147_352 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_42_1018 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6828_ _2961_ _3086_ _3093_ _0305_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_92_434 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_9_274 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_107_216 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6759_ _2977_ _3042_ _3053_ _0276_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_80_629 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_174_193 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_60_331 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_122_219 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6669__A2 _3000_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_103_422 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_115_282 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_131_753 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7330__A3 _3502_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5341__A2 _1509_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_103_477 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7618__A1 _0739_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_53_1147 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_217_356 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_129_2063 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6841__A2 _3087_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7589__C _1950_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_189_208 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5170__S _1446_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4852__A1 core_0.decode.i_imm_pass\[2\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_52_i_clk clknet_4_14__leaf_i_clk clknet_leaf_52_i_clk vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_197_230 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_197_263 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_158_639 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_197_296 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_67_i_clk clknet_4_15__leaf_i_clk clknet_leaf_67_i_clk vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_28_306 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_139_842 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_EDGE_ROW_1_Left_248 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_173_609 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_64_1276 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6357__A1 _1137_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_138_352 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_55_136 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_166_672 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_147 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_138_374 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_607 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_49 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_153_322 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_629 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_83_489 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_12_654 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_70_117 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6109__A1 _2244_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_40_996 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_3_417 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_63_180 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5580__A2 _0177_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_116_1907 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_181_697 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_865 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_153_399 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_231_3279 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_24_578 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_134_591 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_293 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_386 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5868__B1 _2260_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_58 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_121_274 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_208_301 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_clkbuf_leaf_74_i_clk_I clknet_4_13__leaf_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4110_ _0728_ _0729_ _0730_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__7085__A2 _1568_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_166_37 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5090_ _1536_ _1537_ _1538_ _1539_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__5096__A1 _0789_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_235_142 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_235_153 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_223_304 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4041_ _0516_ core_0.execute.rf.reg_outputs\[3\]\[5\] _0548_ _0667_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__6832__A2 _3086_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_75_68 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_246_70 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_188_241 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_78_228 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7800_ _1039_ _1048_ _1069_ _3864_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_0_182_47 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6596__A1 _2929_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5992_ _1676_ _1456_ _2295_ _2382_ _2383_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__5399__A2 _1811_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_188_274 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7793__B1 _3802_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_149_639 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7731_ net179 core_0.decode.i_imm_pass\[10\] _1946_ _3817_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4943_ _1400_ _1403_ _1404_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__3949__A3 _0544_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4071__A2 _0523_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_47_626 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6703__I _3020_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_115_96 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_191_406 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_129_352 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7662_ _1132_ _1048_ _3767_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_4874_ core_0.decode.i_imm_pass\[12\] _1341_ _1351_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_144_300 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6613_ net31 _1149_ _2959_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6899__A2 _3130_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7593_ net205 _3674_ _3712_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__7735__S _1946_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6544_ net129 _2652_ _2906_ _2913_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_132_517 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5571__A2 _0733_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_70_640 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6859__B _3098_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_172_697 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_15_556 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_70_651 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_132_539 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_93 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_113_720 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_171_196 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6475_ _2839_ _2840_ _2851_ _2853_ _2854_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai211_4
X_8214_ _0390_ clknet_leaf_35_i_clk net86 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_2
X_5426_ core_0.execute.alu_mul_div.div_cur\[9\] _1811_ _1866_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__6520__A1 _1380_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_2_461 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_559 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_64_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_112_285 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8145_ _0321_ clknet_leaf_114_i_clk core_0.execute.rf.reg_outputs\[1\]\[4\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_2
XTAP_TAPCELL_ROW_167_2517 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_5357_ _1796_ _1802_ _1804_ _1797_ _1805_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai211_2
XPHY_EDGE_ROW_206_Left_453 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__3885__A2 _0520_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_239_492 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_227_632 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4308_ _0889_ _0843_ _0884_ _0926_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_10_294 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_8076_ _0252_ clknet_leaf_77_i_clk core_0.execute.rf.reg_outputs\[6\]\[15\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_2
X_5288_ _1414_ _1732_ _1736_ _1737_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA_input36_I i_mem_data[9] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7027_ _1371_ _1939_ core_0.execute.alu_mul_div.mul_res\[6\] _3241_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_227_698 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4239_ core_0.fetch.out_buffer_data_instr\[18\] _0858_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__6823__A2 _3086_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_214_326 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4834__A1 _1280_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_241_123 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_199_539 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_241_134 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_97_504 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_69_206 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6036__B1 _2146_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_241_178 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_228 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_179_241 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6587__A1 net35 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8225__CLK clknet_leaf_12_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_210_521 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_210_543 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_84_209 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_167_436 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7929_ _0107_ clknet_leaf_24_i_clk core_0.execute.sreg_priv_control.o_d\[0\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_139_138 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4842__B _1170_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_195_767 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_178_2646 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_215_Left_462 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_37_103 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_78_795 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_194_266 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_100_1708 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_136_801 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6339__A1 _1379_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_191_2802 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_65_489 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_137_Right_137 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_151_815 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5562__A2 _1957_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_61_640 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_865 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6769__B _3057_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_150_314 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_162_174 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_116_580 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4770__B1 _0881_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_104_753 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_60_172 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_131_550 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5314__A2 _1761_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6511__A1 core_0.execute.alu_mul_div.i_mul vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_224_Left_471 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_189_2775 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_189_2786 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_111_1848 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_245_451 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_217_142 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_205_304 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6814__A2 _3065_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_205_337 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_221_808 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_220_307 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_88_537 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_204_2956 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_66_1305 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6578__A1 _2930_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_17_713 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_233_Left_480 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_216_84 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_198_583 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_198_594 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_56_401 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_784 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4053__A2 _0578_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5250__A1 _1693_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_122_1977 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_233_3308 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_185_288 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_232_61 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_126_311 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_71_426 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_37_681 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_142_804 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_154_664 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_4_704 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_104_Right_104 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
X_4590_ core_0.ew_data\[1\] core_0.ew_data\[9\] _1150_ _1160_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__5553__A2 _1955_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6750__A1 _2956_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6679__B _3004_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4600__I1 core_0.ew_data\[14\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_3_214 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_4_737 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_126_399 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_151_2329 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_3_225 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_662 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_673 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_51_150 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_77_1434 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_51_172 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_12_537 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6260_ _2629_ _2631_ _2636_ _2644_ _2645_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai211_2
XANTENNA__6502__A1 _1689_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5211_ _0782_ _0768_ _0776_ core_0.execute.rf.reg_outputs\[2\]\[3\] _1660_ vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_0_86_34 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_110_745 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_177_47 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_209_610 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6191_ _2264_ _2577_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_209_632 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_20_592 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_244_3437 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_5142_ net102 _1492_ _1590_ _1591_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_236_440 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5069__A1 _1466_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_72 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6805__A2 _3065_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5073_ net94 _0521_ _0538_ _0552_ _1461_ _1522_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai221_4
XFILLER_0_208_197 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4024_ _0532_ core_0.execute.rf.reg_outputs\[4\]\[6\] _0519_ _0651_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_2
XTAP_TAPCELL_ROW_162_2458 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_79_526 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4292__A2 _0857_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_88_1563 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_239_Right_239 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_79_548 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_88_1574 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_79_559 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_204_381 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_149_414 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_177_734 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5975_ _2004_ _2284_ _2365_ _2366_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XANTENNA__4044__A2 _0578_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_261 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_710 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_192_704 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7714_ _2251_ _0514_ _3808_ _0476_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4926_ _1381_ _1389_ _1390_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_0_191_203 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_19_136 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_176_277 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_192_737 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5792__A2 _1604_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_47_456 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_75_776 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_47_478 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_75_787 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7645_ _3732_ _3753_ _3754_ _0461_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_4857_ core_0.decode.i_imm_pass\[4\] _1341_ _1342_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_34_139 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7576_ _3682_ _3695_ _3696_ _3697_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_0_117_377 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_133_826 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4788_ _1290_ _1298_ _0060_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__5544__A2 _1957_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_43_640 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_388 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_865 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_173_2587 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_132_325 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_144_185 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6527_ core_0.ew_addr\[0\] _2190_ _2904_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__4888__I net37 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_70_470 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_160_667 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_132_369 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7297__A2 _3391_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_70_492 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6458_ core_0.ew_data\[13\] _2486_ _2838_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_101_734 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_219_418 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5409_ _1233_ _1845_ _1851_ _1822_ _1852_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_6389_ _1061_ _1701_ _2068_ _1109_ _2741_ _2770_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_0_100_233 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5713__S _2113_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_208_3012 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_8128_ _0304_ clknet_leaf_94_i_clk core_0.execute.rf.reg_outputs\[2\]\[3\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_50_1117 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_8059_ _0235_ clknet_leaf_99_i_clk core_0.execute.rf.reg_outputs\[7\]\[14\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__4807__A1 _0869_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_214_123 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_126_2022 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_242_443 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_98_802 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_215_668 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_199_347 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_82_Left_329 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_242_465 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_199_358 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5480__A1 _1909_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6544__S _2906_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_206_Right_206 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_97_367 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_85_518 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7221__A2 core_0.execute.sreg_irq_pc.o_d\[3\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_195_553 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_22_i_clk_I clknet_4_8__leaf_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_168_789 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_219_3141 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_195_586 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_155_417 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_445 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5783__A2 _2183_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_183_748 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_108_311 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_93_562 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_61_1246 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_182_247 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_489 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_19_670 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_108_333 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_53_426 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_136_653 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_124_804 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_182_269 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_25_139 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_19_692 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_137_2151 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_22_771 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_22_782 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6732__A1 _2990_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_91_Left_338 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_137_2162 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_151_623 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4594__I0 core_0.ew_data\[3\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_662 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_150 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4889__A4 core_0.ew_submit vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_312 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_150_155 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_61_492 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_21_334 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_0_206 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_150_177 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_367 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_246_760 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_56_37 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_72_1375 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6799__A1 _2981_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_148_2291 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7460__A2 _3546_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_88_301 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5471__A1 _1375_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_186_520 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_88_367 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7212__A2 _1739_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_202_863 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4026__A2 _0523_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5223__A1 _0771_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_159_767 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_159_778 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_174_715 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5760_ _2148_ _2150_ _2160_ _2161_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_29_434 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_317 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_186_597 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_174_737 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_242 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_158_299 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_173_225 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_139_480 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4711_ _1252_ _1237_ _1254_ _0027_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_173_236 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_573 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5691_ _1720_ _2092_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_17_629 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_122_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_7430_ _0637_ _3544_ _3545_ _3588_ _3589_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_154_450 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4702__S _1246_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_16_139 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_72_757 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4642_ net187 net192 _1199_ _1200_ _1201_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_0_154_461 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_44_459 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_126_163 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_4_512 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6574__I1 core_0.ew_reg_ie\[7\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_112_75 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_112_86 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7361_ _2565_ _2606_ _3530_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_4573_ _1151_ net139 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_130_807 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_142_667 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6312_ _2633_ _2694_ _2166_ _2695_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_0_97_33 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7279__A2 _3393_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_12_334 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7292_ net75 _3398_ _3399_ _3468_ _3469_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_188_68 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_141_188 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_122_380 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_12_378 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6243_ _2026_ _2034_ _2628_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_122_391 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_0_784 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6174_ _1600_ _2374_ _2560_ _1479_ _2561_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XPHY_EDGE_ROW_139_Left_386 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_110_597 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5125_ core_0.execute.rf.reg_outputs\[7\]\[10\] net232 _1443_ core_0.execute.rf.reg_outputs\[3\]\[10\]
+ _1574_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_224_454 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5056_ _1466_ net193 _1505_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_137_72 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_212_605 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_27_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4007_ net102 _0578_ _0636_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_79_323 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_211_115 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_196_317 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_95_816 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7203__A2 _1381_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4017__A2 _0523_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1_72 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_220_671 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_0_499 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_148_Left_395 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_109_108 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_137_417 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_149_288 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_164_214 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_175_2616 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_5958_ core_0.execute.irq_en _1385_ _2249_ core_0.execute.pc_high_buff_out\[2\] _2349_
+ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_47_242 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_776 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_702 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4909_ _1373_ _1374_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_164_247 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_275 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_201 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5889_ _2280_ _2281_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_118_653 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_426 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5708__S _1819_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_106_804 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_145_450 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7628_ core_0.execute.pc_high_buff_out\[2\] _3731_ _1216_ _3742_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__6714__A1 core_0.execute.rf.reg_outputs\[5\]\[4\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_90_554 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_133_623 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_90_565 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_145_483 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_106_859 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_132_111 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_172_291 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_150 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_214_3082 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_7559_ _3681_ _3682_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_43_481 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_31_632 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_132_177 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_31_676 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_31_698 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_132_2092 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_30_186 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_186_2745 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7690__A2 _1092_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_234_229 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7442__A2 _3546_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_188_807 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6782__B _3057_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4256__A2 _0727_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5453__A1 core_0.execute.alu_mul_div.div_cur\[12\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_97_142 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_230_457 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_230_468 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_201_2926 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_27_841 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4008__A2 _0635_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_210_170 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_197_2874 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_128_417 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5756__A2 _2019_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6953__A1 core_0.execute.alu_mul_div.mul_res\[0\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_156_737 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_168_597 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_66_551 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_264 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_404 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_26_415 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_212 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_297 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5618__S _1492_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_26_437 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_183_578 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_53_223 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_124_601 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_163 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6556__I1 _2859_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_53_267 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_170_239 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_109 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_124_645 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_610 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_112_807 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_34_470 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6181__A2 _2567_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_124_667 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_492 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_74_1404 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_123_188 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_142 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_153 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_104_380 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7130__A1 _2855_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_67_69 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7681__A2 _1056_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5692__A1 _1714_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_241_3407 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_246_590 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5152__I _1600_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_174_37 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_233_240 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_206_465 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5444__A1 _1233_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_83_57 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_233_273 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_206_498 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6930_ _1221_ _3150_ _3151_ _0349_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_88_120 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_178_317 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_107_53 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_85_1533 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6861_ _0722_ _3112_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_159_542 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_186_350 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5812_ _2202_ _2208_ _2210_ _0171_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_119_417 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6792_ core_0.execute.rf.reg_outputs\[3\]\[5\] _3070_ _3072_ _3073_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_146_203 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5747__A2 _2146_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6944__A1 _1915_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_174_523 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_648 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_702 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_125 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_57_562 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5743_ _1653_ _2142_ _2143_ _2144_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_146_247 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_32_61 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_426 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_174_589 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5674_ _1701_ _1501_ _2075_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_161_228 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_127_494 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7413_ core_0.execute.sreg_irq_pc.o_d\[5\] _3542_ _3516_ _3575_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4625_ core_0.dec_jump_cond_code\[2\] _1182_ _1183_ _1184_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_0_142_442 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_199_78 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6172__A2 net223 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_170_2557 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_25_492 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_13_632 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_4_364 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4183__A1 core_0.decode.o_submit vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7344_ _3514_ _2888_ _3502_ _3515_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_96_1662 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_102_317 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4556_ _1078_ _1092_ _1138_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_114_177 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6867__B _3112_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7275_ net73 net87 _3439_ _3454_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and3_1
XANTENNA__7121__A1 _2797_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4487_ _1056_ _1073_ _1080_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_6226_ _2586_ _2611_ _2356_ _2612_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__5490__C _1226_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_229_568 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__7672__A2 _1053_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_244_527 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4486__A2 _1072_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6157_ _2244_ _2542_ _2543_ _2544_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_99_407 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_5_569 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_5108_ net95 _0521_ _0703_ _0708_ _1460_ _1557_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai221_4
XANTENNA__7424__A2 _3544_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6088_ _2295_ _2459_ _2476_ _2477_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XANTENNA__4238__A2 net48 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5435__A1 _1233_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_240_733 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_212_424 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5039_ _0789_ core_0.execute.rf.reg_outputs\[4\]\[13\] _0779_ _1488_ vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_79_120 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_181_2686 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_196_103 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_164_70 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_212_457 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_67_304 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_79_164 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_156_Left_403 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_164_92 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_94_101 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_24_800 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output105_I net105 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4406__I net82 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_67_348 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6935__A1 _1915_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_138_737 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_45_1049 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_216_3100 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_82_329 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_165_556 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4410__A2 _0966_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_153_718 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_192_364 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6538__I1 _2526_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7735__I0 net181 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_152_228 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_105_100 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_35_267 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_134_2121 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_50_215 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7360__A1 _2477_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_106_667 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_44_790 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_133_464 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_166 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_165_Left_412 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_105_177 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_120_103 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5910__A2 _1491_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_105_199 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_462 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_208_708 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7953__CLK clknet_leaf_4_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_56_1189 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7663__A2 _3766_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput75 net75 dbg_pc[12] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XTAP_TAPCELL_ROW_227_3240 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
Xoutput86 net86 dbg_pc[8] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA__5674__A1 _1701_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4477__A2 _1068_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput97 net97 dbg_r0[3] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_207_218 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_108_1809 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_145_2250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4229__A2 _0843_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5426__A1 core_0.execute.alu_mul_div.div_cur\[9\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_199_2903 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7401__B _3553_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_174_Left_421 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_231_733 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_231_744 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_16 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_98_451 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_59_816 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3988__A1 _0533_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_187_158 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7179__A1 _1748_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6926__A1 _2996_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_551 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_86_679 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_168_383 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_562 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_702 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_184_843 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_195_191 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_184_865 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6531__I _2189_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_80_1474 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_143_206 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_156_589 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_543 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_863 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_171_537 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_26_267 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_119_1938 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_30_869 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_156_2390 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_183_Left_430 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__7351__A1 net213 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4410_ _1013_ _0966_ _1015_ _1016_ _0877_ net171 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XANTENNA__7790__C _1950_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_151_261 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5390_ _1747_ _1830_ _1835_ _0125_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_1
XANTENNA__6687__B _3004_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_78_57 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_4341_ _0946_ _0959_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA__4986__I _1434_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7060_ _2648_ _3181_ _3272_ _0358_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4272_ core_0.fetch.prev_request_pc\[9\] _0890_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_238_387 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_226_527 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6011_ core_0.dec_sreg_irt _2400_ _2401_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_94_34 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_241_508 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7406__A2 _1013_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_241_519 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_118_74 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_27_72 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_2_539 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_7962_ _0140_ clknet_leaf_77_i_clk core_0.de_jmp_pred vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_221_232 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_38_969 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3979__A1 _0568_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6913_ net103 _3135_ _3139_ _3142_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_7893_ _0084_ clknet_leaf_71_i_clk core_0.decode.i_imm_pass\[2\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_2
XANTENNA__4640__A2 net184 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_194_629 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_159_2419 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_221_298 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6844_ core_0.execute.rf.reg_outputs\[2\]\[12\] _3092_ _3098_ _3102_ vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__6917__A1 net90 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_147_534 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_119_236 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_69_i_clk_I clknet_4_15__leaf_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_18_724 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_92_638 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7590__A1 core_0.execute.pc_high_out\[5\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_190_802 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3987_ core_0.execute.rf.reg_outputs\[7\]\[9\] _0530_ _0617_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6775_ core_0.execute.rf.reg_outputs\[4\]\[15\] _3041_ _3057_ _3062_ vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_119_269 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_17_223 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_489 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5726_ _1124_ _1541_ _2127_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_17_245 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_94_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_17_267 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_162_559 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_72_373 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6145__A2 _2257_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5657_ _2056_ _2057_ _2058_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_4
XANTENNA__7342__A1 _3510_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_211_3041 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_115_475 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_130_412 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4608_ _0726_ _0727_ _0813_ _1168_ _1169_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai211_4
XFILLER_0_4_172 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5588_ _1711_ _1719_ _1989_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_103_648 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_input66_I i_req_data[6] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4539_ _1123_ _1124_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
X_7327_ _2477_ _2521_ _3500_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_229_343 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7258_ net86 net85 _3426_ _3439_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and3_1
XTAP_TAPCELL_ROW_183_2704 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_245_836 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5656__A1 _1789_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4459__A2 _1053_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_244_324 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6209_ _1600_ _2409_ _2595_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or2_1
X_7189_ _1748_ _3379_ _0380_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__5721__S _2102_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_245_28 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5408__A1 _1232_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6616__I _2935_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5520__I _1051_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5959__A2 _2254_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_222_3181 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_197_434 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_213_766 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_240_563 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_68_646 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_140_2191 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_138_545 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_165_331 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_194_2844 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_165_342 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_166_865 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_36_521 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6384__A2 _1455_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_153_504 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7581__A1 _3673_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_181_813 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_193_695 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_64_863 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_565 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_51_502 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_727 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_513 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6136__A2 _2332_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7333__A1 _2777_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_90_170 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xrebuffer8 net228 net230 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlya_2
XFILLER_0_140_209 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_58_1207 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_161_570 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_51_579 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3924__B _0520_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_210_97 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7097__B1 _3300_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_121_489 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_114_1879 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7636__A2 _3731_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_208_527 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_219_84 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_64_37 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4870__A2 _1341_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4247__S _0725_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_69_1336 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_235_50 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8281__CLK clknet_leaf_29_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_207_2998 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_235_61 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6072__A1 _2013_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_235_72 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_203_276 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_148_309 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_35_928 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4046__I _0671_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_98_292 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_668 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3910_ _0539_ core_0.execute.rf.reg_outputs\[4\]\[15\] _0520_ _0546_ vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_4890_ _0806_ _1358_ _1284_ _0102_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_86_476 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_70_i_clk_I clknet_4_15__leaf_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_74_627 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_156_331 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_236_3339 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6375__A2 _2531_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_172_802 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7572__A1 core_0.execute.pc_high_out\[2\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_392 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_15_696 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7999__CLK clknet_leaf_119_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6560_ core_0.dec_rf_ie\[0\] core_0.ew_reg_ie\[0\] _1985_ _2921_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_183_183 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5511_ core_0.execute.alu_mul_div.div_cur\[0\] _1812_ _1943_ _1841_ _1944_ vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_171_356 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_42_524 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_54_384 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_125_751 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6491_ _0563_ _2869_ _2241_ _2870_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_202_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_70_855 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_89_67 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5442_ _1879_ _1791_ _1880_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_8230_ _0406_ clknet_leaf_13_i_clk core_0.execute.sreg_irq_pc.o_d\[2\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5886__A1 core_0.ew_data\[1\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_93_1632 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_5373_ _1374_ _1820_ _1821_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_8161_ _0337_ clknet_leaf_88_i_clk net98 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_4
XFILLER_0_1_142 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_1_164 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4324_ _0872_ _0939_ _0941_ _0942_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_4
X_7112_ _3319_ _3320_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_8092_ _0268_ clknet_leaf_77_i_clk core_0.execute.rf.reg_outputs\[5\]\[15\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_239_696 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7043_ _2587_ _3181_ _3256_ _0357_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_227_858 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4255_ _0864_ _0867_ _0868_ _0873_ _0874_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_0_38_71 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_129_84 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4186_ net156 _0805_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__inv_1
XTAP_TAPCELL_ROW_165_2489 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4861__A2 _1341_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_241_349 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4384__C _0877_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6063__A1 net82 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_179_434 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6063__B2 _2245_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7945_ _0123_ clknet_leaf_7_i_clk core_0.execute.alu_mul_div.div_cur\[1\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_49_112 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_145_94 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_118_Right_118 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
X_7876_ _0067_ clknet_leaf_83_i_clk core_0.decode.i_instr_l\[1\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_64_104 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_65_627 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_77_487 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_92_413 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6827_ core_0.execute.rf.reg_outputs\[2\]\[4\] _3092_ _3083_ _3093_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__7563__A1 net201 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6366__A2 core_0.execute.alu_mul_div.mul_res\[11\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_42_1019 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_18_521 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_137 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_206 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_108_729 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4377__A1 _0837_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_92_457 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__8004__CLK clknet_leaf_48_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_46_863 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_190_632 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6758_ core_0.execute.rf.reg_outputs\[4\]\[7\] _3049_ _3045_ _3053_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_135_537 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_373 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5709_ _2106_ _2109_ _2102_ _2110_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__7315__A1 _2893_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6689_ core_0.execute.rf.reg_outputs\[6\]\[10\] _3006_ _3004_ _3013_ vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__4129__A1 core_0.execute.pc_high_out\[5\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_5_492 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5877__A1 core_0.dec_sreg_irt vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output172_I net172 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_60_387 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_130_242 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_131_765 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6120__B _2013_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_590 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5515__I _1063_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_103_489 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_245_600 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5629__A1 _1761_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_53_1148 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_129_2064 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_233_839 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4852__A2 _1307_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_225_390 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_198_732 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_142_2220 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_87_229 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_198_776 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4065__B1 _0521_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_158_607 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_68_454 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_96_763 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_465 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_200_257 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_154_802 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7554__A1 core_0.execute.pc_high_out\[0\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_64_1277 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6357__A2 _1568_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_181_632 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_193_492 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_36_351 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_165_183 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_12_655 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_153_345 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_384 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_524 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_63_170 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_113_209 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_40_997 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_52_855 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_116_1908 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_122_710 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_229 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5868__B2 net1 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4540__A1 _1066_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_17_i_clk_I clknet_4_8__leaf_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_208_313 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_209_847 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_102_Left_349 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__6457__S _2242_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_235_132 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4040_ _0515_ _0523_ _0525_ core_0.execute.rf.reg_outputs\[2\]\[5\] _0666_ vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_0_208_379 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_236_699 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_235_187 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4843__A2 _1333_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_189_743 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6045__A1 _2281_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_410 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5991_ _2294_ _2381_ _2382_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__7793__A1 core_0.decode.i_instr_l\[15\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_152_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_182_59 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_59_432 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_149_629 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_231_382 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7793__B2 core_0.decode.i_instr_l\[12\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8027__CLK clknet_leaf_53_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7730_ _3816_ _0484_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4942_ net204 _1403_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_86_251 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_87_774 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_148_139 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4932__C _1395_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_307 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4071__A3 _0526_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_487 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_86_262 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_111_Left_358 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_157_640 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_46_104 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_74_413 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_46_115 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_74_424 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7661_ _1132_ _3766_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
X_4873_ _0854_ _1321_ _1350_ _0093_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__7545__A1 net77 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_7_702 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_117_504 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_74_457 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6612_ net24 _1148_ _2958_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_144_312 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_863 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_537 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_156_172 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7592_ core_0.execute.pc_high_buff_out\[5\] _3682_ _3710_ _3711_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_184_492 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_171_120 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8177__CLK clknet_leaf_129_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6543_ _2912_ _0201_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_171_142 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_54_181 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_70_663 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_505 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6474_ _1993_ _2178_ _2852_ _2853_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_8213_ _0389_ clknet_leaf_33_i_clk net85 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_4
XFILLER_0_42_387 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_527 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_140_540 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput210 net210 sr_bus_we vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XPHY_EDGE_ROW_12_Right_12 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
X_5425_ _1812_ _1864_ _1865_ _0130_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_113_776 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_140_584 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4531__A1 _1117_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_120_Left_367 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_11_763 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8144_ _0320_ clknet_leaf_118_i_clk core_0.execute.rf.reg_outputs\[1\]\[3\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5356_ core_0.execute.alu_mul_div.div_cur\[12\] _1803_ _1799_ _1804_ vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
XTAP_TAPCELL_ROW_167_2518 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6875__B _3112_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5874__A4 _2266_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_10_273 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4307_ core_0.fetch.prev_request_pc\[15\] _0827_ _0886_ core_0.fetch.prev_request_pc\[14\]
+ _0925_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_8075_ _0251_ clknet_leaf_77_i_clk core_0.execute.rf.reg_outputs\[6\]\[14\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5287_ _1735_ _1736_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XANTENNA__5087__A2 _1484_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4238_ _0824_ net48 _0856_ _0857_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_4
X_7026_ _1620_ _3178_ _3240_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA_input29_I i_mem_data[2] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4834__A2 net41 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4169_ core_0.ew_reg_ie\[5\] _0779_ _0788_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6036__A1 _1121_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6036__B2 _1107_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_21_Right_21 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_195_702 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4047__B1 _0662_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_195_713 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7784__A1 _1136_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_179_264 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_195_724 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_179_286 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7928_ _0106_ clknet_leaf_129_i_clk core_0.execute.alu_mul_div.cbit\[3\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_77_240 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_78_763 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_210_555 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_38_605 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_195_757 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_194_234 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_178_2647 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_38_638 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7859_ _0051_ clknet_leaf_61_i_clk core_0.fetch.prev_request_pc\[2\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_2
XANTENNA__6115__B _2010_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_100_1709 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_37_137 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_191_2803 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_148_684 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_182_429 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_65_457 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_92_243 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_163_610 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_619 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_135_334 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_310 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_190_473 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_395 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_150_304 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_855 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_163_698 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4770__A1 core_0.fetch.prev_request_pc\[3\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_104_721 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4770__B2 net170 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_30_Right_30 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA_output97_I net97 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_376 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_60_162 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_398 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_765 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6511__A2 core_0.execute.alu_mul_div.mul_res\[15\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_131_573 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_29_18 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_189_2776 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_111_1849 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6275__A1 _2447_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_245_463 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_233_625 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_206_839 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_205_349 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6027__A1 _1601_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_66_1306 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_213_360 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_204_2957 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4038__B1 _0662_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6578__A2 _1985_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7775__A1 core_0.decode.i_instr_l\[7\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_17_714 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_185_212 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_68_251 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_711 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_627 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_104 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_139_640 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_115 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_126 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_435 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_122_1978 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_233_3309 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_194_790 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_56_479 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_37_693 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_24_310 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_24_321 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_126_378 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6750__A2 _3042_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_153_164 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_151_2319 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_12_516 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_77_1435 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_24_387 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_12_527 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_101_66 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5210_ _0771_ _0768_ _0776_ core_0.execute.rf.reg_outputs\[6\]\[3\] _1659_ vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_0_177_26 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4513__A1 core_0.decode.i_instr_l\[3\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_228_419 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6190_ _2201_ _2576_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_86_57 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5141_ _1586_ _1587_ _1588_ _1589_ _1590_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_0_110_779 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_244_3438 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_208_121 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5069__A2 net189 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6266__A1 core_0.execute.alu_mul_div.div_cur\[8\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
X_5072_ _1467_ net184 _1521_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_4023_ core_0.execute.rf.reg_outputs\[7\]\[6\] _0529_ _0650_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_162_2459 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_126_41 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_88_1564 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_189_562 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_177_702 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_126_74 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_220_831 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_72 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_126_85 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_149_426 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_94_519 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_177_746 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5974_ _1596_ _2005_ _2365_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_59_273 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7713_ core_0.decode.i_imm_pass\[1\] _1064_ _3808_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4925_ _0810_ _1388_ _1389_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__7518__A1 _0637_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_74_221 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_75_766 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_243 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7644_ core_0.execute.pc_high_buff_out\[6\] _3731_ _1216_ _3754_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_191_237 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_159 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_28_660 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_117_323 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_145_632 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_157_492 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4856_ _1305_ _1341_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_34_107 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_191_259 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7575_ core_0.execute.pc_high_out\[3\] _3688_ _3696_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_4787_ core_0.fetch.prev_request_pc\[11\] net225 _0880_ net163 _1298_ vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_0_16_855 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_133_838 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_160_635 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_173_2588 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4752__A1 net61 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6526_ _2576_ _2902_ _2903_ _0193_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xclkbuf_leaf_51_i_clk clknet_4_12__leaf_i_clk clknet_leaf_51_i_clk vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_42_162 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_31_836 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_30_302 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_42_173 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_313 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6457_ _0580_ _2836_ _2242_ _2837_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_31_858 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_101_702 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_113_562 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_113_573 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4504__A1 _1046_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_30_368 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5408_ _1232_ _1850_ _1851_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_140_381 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_30_379 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6388_ _2080_ _2175_ _2769_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_208_3013 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_66_i_clk clknet_4_15__leaf_i_clk clknet_leaf_66_i_clk vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_8127_ _0303_ clknet_leaf_110_i_clk core_0.execute.rf.reg_outputs\[2\]\[2\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5339_ core_0.execute.alu_mul_div.div_cur\[9\] _1754_ _1787_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_50_1107 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6257__A1 _2412_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_50_1118 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_8058_ _0234_ clknet_leaf_99_i_clk core_0.execute.rf.reg_outputs\[7\]\[13\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_214_102 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_215_636 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4807__A2 core_0.fetch.submitable vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_126_2023 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output135_I net135 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_199_326 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7009_ _3183_ _3184_ _1229_ _3225_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_215_658 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_170_Right_170 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__5480__A2 _1576_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_97_324 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_168_702 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_183_80 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_195_510 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_168_724 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_211_842 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_167_212 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_222_190 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_195_543 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4035__A3 _0518_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_219_3142 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7509__A1 net227 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_65_221 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_457 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6560__S _1985_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_66_777 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_176_790 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_53_405 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_61_1247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_93_574 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_202_43 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_135_142 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_137_2152 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_151_602 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_34_630 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_22_772 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6732__A2 _3022_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_19_i_clk clknet_4_8__leaf_i_clk clknet_leaf_19_i_clk vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__4594__I1 core_0.ew_data\[11\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_123_348 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_346 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7693__B1 _1092_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_72_1376 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_56_49 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_246_794 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_206_636 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6799__A2 _3064_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_233_422 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_206_647 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_148_2292 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_205_135 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_205_146 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_88_313 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_89_836 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_89_858 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_72_37 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_198_381 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_159_735 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7212__A3 _1734_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_186_543 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_201_352 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4026__A3 _0526_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_186_554 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5223__A2 _0768_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6420__A1 _1803_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_56_210 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_766 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_17_608 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_72_703 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4710_ net40 _1253_ _1254_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__7793__C _1133_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_139_492 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5690_ net211 _2091_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_16_107 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4989__I _1437_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_56_298 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4641_ net193 net180 net179 net182 _1200_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or4_2
XFILLER_0_142_613 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6723__A2 _3027_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_25_641 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_115_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_4_524 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_71_257 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4572_ core_0.ew_data\[0\] net157 _1151_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
X_7360_ _2477_ _2521_ _3529_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_142_646 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_112_98 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_12_302 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_13_836 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6311_ _2036_ _2040_ _2694_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
X_7291_ _3466_ _3467_ _3468_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_13_858 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_97_56 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8215__CLK clknet_leaf_36_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6242_ _1831_ _1700_ _1721_ _2133_ _2114_ _2627_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai32_2
X_6173_ _1600_ _2370_ _2560_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_110_587 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_237_772 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5124_ _0782_ core_0.execute.rf.reg_outputs\[4\]\[10\] _0778_ _1573_ vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_236_271 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_209_485 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5055_ _0630_ _0635_ _0636_ _1460_ _1504_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai31_4
XFILLER_0_137_84 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4006_ _0631_ _0632_ _0633_ _0634_ _0635_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_4
XANTENNA__5462__A2 _1817_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_211_105 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_79_335 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_79_368 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_149_223 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_177_543 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6411__A1 _1380_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4017__A3 _0526_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_153_72 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_733 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_94_349 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_149_278 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5957_ core_0.execute.sreg_irq_flags.o_d\[2\] _2250_ _2257_ core_0.execute.pc_high_out\[2\]
+ _2348_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_TAPCELL_ROW_175_2617 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_192_524 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_192_535 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_47_1080 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_118_621 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4908_ _1372_ _1367_ _1227_ _1230_ _1373_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor4_4
XANTENNA__4973__B2 _1390_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5888_ core_0.execute.alu_mul_div.i_mul _2280_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_8_863 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_522 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7627_ net221 _3733_ _3740_ _3741_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_117_142 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4839_ _1328_ _1330_ _0079_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6714__A2 _3027_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_62_257 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7558_ _3637_ _1953_ _1205_ _3681_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_2
XTAP_TAPCELL_ROW_214_3083 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_133_679 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6509_ _1719_ _1455_ _2887_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_7489_ core_0.execute.sreg_jtr_buff.o_d\[1\] _1398_ _1206_ _3636_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__6478__A1 _1088_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_113_381 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_101_543 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_132_2093 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_219_227 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7224__B _3409_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_186_2746 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5150__A1 _1467_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_243_720 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_227_271 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_215_411 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_227_282 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_215_422 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_230_403 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_188_819 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5453__A2 _1812_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_187_307 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_97_121 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_202_149 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_201_2927 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_27_831 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_27_842 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_58_519 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_86_839 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6402__A1 core_0.execute.alu_mul_div.div_cur\[12\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_211_683 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_733 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_349 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_197_2875 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_195_395 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4964__A1 _1301_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_183_557 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_449 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_109_676 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6705__A2 _3022_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_136_473 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_191_590 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4716__A1 net42 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_163_292 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_62_780 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_599 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_151_454 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_123_156 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_74_1405 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6469__A1 _1137_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6469__B2 _1109_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5516__I0 core_0.de_jmp_pred vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_10_839 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7130__A2 _1941_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4758__B _1280_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_120_863 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_219_772 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5692__A2 _1592_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_241_3408 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6641__A1 _2936_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_83_69 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3888__I _0523_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_89_655 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_85_1534 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_221_469 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_74 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6860_ _2951_ _3107_ _3111_ _0319_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_190_37 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5811_ net133 _2209_ _2210_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_9_616 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_232_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_57_530 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6791_ _1963_ _3072_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_8_104 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6944__A2 _1803_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4955__A1 _1400_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5742_ _1558_ _1652_ _2143_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_57_574 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_360 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_213 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_162_719 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5673_ _2072_ _2073_ _2074_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_45_769 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_127_484 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7412_ net227 _3544_ _3573_ _3574_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XPHY_EDGE_ROW_6_Right_6 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
X_4624_ core_0.dec_jump_cond_code\[1\] core_0.dec_jump_cond_code\[0\] core_0.execute.alu_flag_reg.o_d\[0\]
+ _1183_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
XTAP_TAPCELL_ROW_170_2547 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6172__A3 _1555_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_142_454 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_170_2558 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4183__A2 _0801_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5380__A1 _1232_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7343_ net202 _3514_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_12_121 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4555_ core_0.decode.oc_alu_mode\[2\] _1137_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XTAP_TAPCELL_ROW_96_1663 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_4_387 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7274_ net87 _3439_ net73 _3453_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__7121__A2 _3328_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4486_ _1078_ _1072_ _1079_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5132__A1 _0789_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6225_ _2608_ _2609_ _2610_ _2611_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_4
XANTENNA_clkbuf_leaf_65_i_clk_I clknet_4_15__leaf_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_110_373 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6880__A1 _2988_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6156_ _2455_ _2495_ _2541_ _2543_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_225_720 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_209_282 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_225_742 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_209_293 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5107_ _1466_ net185 _1556_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_99_419 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_224_241 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6087_ _2464_ _2475_ _2476_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_224_252 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6632__A1 net34 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_224_263 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5038_ core_0.execute.rf.reg_outputs\[5\]\[13\] _1486_ _1487_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_181_2687 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input11_I i_core_int_sreg[4] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_197_627 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_169_318 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_79_132 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_839 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7188__A2 _3372_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_196_159 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_24_801 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5199__A1 _0782_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4246__I0 net66 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6989_ _3198_ _3206_ _3175_ _3207_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__6935__A2 _1689_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_105_1770 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_216_3101 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4946__A1 _1195_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_48_563 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_63_500 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_75_360 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_94_179 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_192_354 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_522 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6148__B1 _2534_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_91_842 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_235 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_192_387 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6123__B _1456_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_118_473 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5518__I net104 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_180_527 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_63_566 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_408 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6699__A1 _2994_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_35_279 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_23_419 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_134_2122 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_63_599 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_16_471 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7360__A2 _2521_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_133_476 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_189 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_160_295 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3921__A2 _0530_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_102_863 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_56_1179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
Xoutput76 net76 dbg_pc[13] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
Xoutput87 net87 dbg_pc[9] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XTAP_TAPCELL_ROW_227_3241 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_235_528 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5674__A2 _1501_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4477__A3 _1069_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput98 net98 dbg_r0[4] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_228_580 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6285__S _2102_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_215_252 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4229__A3 _0844_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6623__A1 core_0.execute.rf.reg_outputs\[7\]\[5\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5426__A2 _1811_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_145_2251 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_215_263 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_188_605 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_199_2904 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_188_616 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_208_97 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_187_115 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3988__A2 core_0.execute.rf.reg_outputs\[4\]\[9\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_86_614 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_98_474 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6226__I1 _2611_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_85_113 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_196_660 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_230_299 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_184_811 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_224_74 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6926__A2 _3130_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_73_308 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6812__I _1963_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_183_321 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_238_3370 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_128_259 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_393 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_80_1475 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_171_516 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_171_527 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_59_Right_59 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_109_484 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_54_566 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_352 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_152_730 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_54_588 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_119_1939 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_156_2380 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_41_216 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_81_385 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__7351__A2 _3502_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_124_454 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_112_605 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_124_465 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5362__A1 core_0.execute.alu_mul_div.comp vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4165__A2 _0782_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_124_476 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_111_104 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4340_ core_0.fetch.prev_request_pc\[15\] _0957_ _0958_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_238_311 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1_346 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5114__A1 _0789_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4271_ core_0.fetch.prev_request_pc\[8\] _0889_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__inv_1
X_6010_ net81 _2268_ _2399_ _2245_ _2400_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XANTENNA_input3_I i_core_int_sreg[11] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_68_Right_68 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_182_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_219_591 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_118_31 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6614__A1 _2929_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_222_734 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7961_ _0139_ clknet_leaf_17_i_clk core_0.execute.hold_valid vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_206_296 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_179_638 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_221_244 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6090__A2 _2477_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_77_603 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_89_463 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6912_ _2981_ _3129_ _3141_ _0341_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_7892_ _0083_ clknet_leaf_71_i_clk core_0.decode.i_imm_pass\[1\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_178_159 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_159_340 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_49_338 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_76_124 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_77_647 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4640__A3 net183 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6843_ _2988_ _3087_ _3101_ _0312_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_49_349 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_77_658 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_413 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6917__A2 _3135_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_43_72 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_76_157 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_186_181 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_174_321 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4928__A1 core_0.execute.prev_sys vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6774_ _2994_ _3043_ _3061_ _0283_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_3986_ core_0.execute.rf.reg_outputs\[1\]\[9\] _0616_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XPHY_EDGE_ROW_77_Right_77 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_91_127 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_73_842 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_190_825 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5725_ _2091_ _2092_ _2126_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_162_527 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_174_387 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_115_432 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_150_73 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_279 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5656_ _1789_ _1576_ _2057_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_143_752 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_32_227 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_142_240 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_547 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4607_ core_0.decode.i_flush core_0.fetch.flush_event_invalidate _1168_ vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_2
XTAP_TAPCELL_ROW_211_3042 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_4_162 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_102_104 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5587_ _1987_ _1549_ _1988_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_142_295 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_41_772 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7326_ _2565_ _2606_ _3499_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4538_ core_0.decode.oc_alu_mode\[12\] _1123_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XANTENNA__4398__B _0970_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_13_485 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_130_457 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_7_72 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_159_60 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input59_I i_req_data[29] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_111_660 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7257_ _3433_ _3434_ _3438_ _0389_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_159_82 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4469_ _1052_ _1062_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XPHY_EDGE_ROW_86_Right_86 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_111_693 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5656__A2 _1576_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_183_2705 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6208_ _1550_ _1700_ _2594_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_110_181 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_245_848 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7188_ _3367_ _3372_ core_0.execute.alu_mul_div.div_res\[13\] _3379_ vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_6139_ _2360_ _2526_ _2527_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_99_216 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6605__A1 _2936_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7221__C _1736_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_213_734 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_212_222 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_222_3171 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_222_3182 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_212_244 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_67_102 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_95_422 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_240_597 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_68_658 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_166_811 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_184_107 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_191_80 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_669 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_95_Right_95 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_138_524 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_166_833 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_184_129 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7030__A1 _1908_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_83_617 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_138_535 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_140_2192 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6464__S0 _2294_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4919__A1 net185 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_177_181 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_194_2845 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5041__B1 _1435_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_193_674 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_382 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_138_579 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5592__A1 _1713_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_165_387 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_63_341 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_63_352 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4152__I _0770_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_91_683 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7920__CLK clknet_leaf_8_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_106_454 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_23_238 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_58_1208 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_15_Left_262 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__7097__A1 core_0.execute.alu_mul_div.mul_res\[10\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_121_479 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7097__B2 core_0.execute.alu_mul_div.mul_res\[11\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_102_671 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_236_804 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_101_181 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_223_509 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_204_712 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_216_594 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_69_1337 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_207_2999 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6998__I2 _1929_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_24_Left_271 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_99_772 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_204_778 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_188_457 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_35_929 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_80_26 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_80_37 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_clkbuf_leaf_13_i_clk_I clknet_4_9__leaf_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_74_617 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_105 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_184_663 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7572__A2 _3672_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_842 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_27_544 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_183_162 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_156_387 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_15_697 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_13_86 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_801 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_82_661 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5510_ _1811_ _1942_ _1943_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_125_741 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_89_35 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6490_ _2360_ _2859_ _2868_ _2869_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_125_763 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6698__B _3016_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_81_182 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_124_240 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_33_Left_280 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__5335__A1 core_0.execute.alu_mul_div.div_cur\[8\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
X_5441_ _1794_ _1878_ _1879_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_112_424 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_772 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_112_446 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8160_ _0336_ clknet_leaf_88_i_clk net97 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_4
XANTENNA__5886__A2 _2209_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5372_ core_0.execute.alu_mul_div.div_cur\[0\] _1819_ _1820_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_93_1633 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_112_457 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6210__C _1765_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7088__A1 _1224_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7111_ _2778_ _3313_ _3319_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_112_479 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_196_47 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4323_ _0867_ _0940_ _0941_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_8091_ _0267_ clknet_leaf_98_i_clk core_0.execute.rf.reg_outputs\[5\]\[14\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__6835__A1 core_0.execute.rf.reg_outputs\[2\]\[8\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_227_837 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_226_314 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7042_ _3240_ _3255_ _3189_ _3256_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4254_ _0869_ _0870_ _0872_ _0873_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_242_818 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4185_ _0802_ _0803_ _0804_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_0_241_317 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6063__A2 _2268_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7944_ _0122_ clknet_leaf_14_i_clk net72 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_4
XANTENNA__4074__A1 _0567_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_54_82 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_89_282 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_222_597 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_210_737 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_166_107 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7875_ _0066_ clknet_leaf_83_i_clk core_0.decode.i_instr_l\[0\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_194_449 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6826_ _3085_ _3092_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_147_343 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_102_1740 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_161_72 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_147_376 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_162_302 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5574__A1 _1980_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4377__A2 _0947_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6757_ _2972_ _3042_ _3052_ _0275_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_163_836 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3969_ _0517_ _0524_ _0527_ core_0.execute.rf.reg_outputs\[2\]\[11\] _0601_ vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_0_45_352 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_163_858 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5708_ _2107_ _2108_ _1819_ _2109_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_60_300 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6688_ _2983_ _2999_ _3012_ _0246_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_61_834 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_190_677 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7315__A2 _3393_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_116_774 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_150_519 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5326__A1 core_0.execute.alu_mul_div.div_cur\[3\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
X_5639_ _1756_ _1591_ _2040_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_0_13_282 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7309_ net77 _3398_ _3399_ _3483_ _3484_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_218_804 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8289_ _0465_ clknet_leaf_45_i_clk core_0.dec_mem_width vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5629__A2 _2019_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_229_174 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_53_1149 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_224_3200 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_218_859 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_217_336 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_245_656 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_244_133 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_129_2065 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_232_317 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_142_2221 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7251__A1 _2611_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_198_744 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_240_361 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_201_726 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4065__B2 net97 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_198_788 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_200_214 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_200_225 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_444 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3986__I core_0.execute.rf.reg_outputs\[1\]\[9\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_200_247 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_138_310 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_403 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_83_414 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_138_332 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_64_1278 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_126_505 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_842 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_165_162 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_138_387 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_138_398 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_153_324 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_64_661 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_165_195 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_12_656 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_107_752 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_153_368 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_40_987 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_40_998 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_51_333 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5317__A1 _1461_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_116_1909 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_153_2350 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_181_699 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_134_571 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_122_722 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_122_733 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_208 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_161_390 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4610__I _1170_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5868__A2 _1385_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4540__A2 _1056_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_184_Right_184 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_209_826 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_37 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_246_3480 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_236_667 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_216_391 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6045__A2 _2434_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5990_ _2123_ _2109_ _2301_ _1721_ _2381_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_0_59_422 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7793__A2 _3786_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_204_597 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_148_107 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_87_753 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4941_ _1301_ _1402_ _0109_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_188_287 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3896__I core_0.dec_r_reg_sel\[2\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_4_0__f_i_clk_I clknet_3_0_0_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_145_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_115_76 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7660_ _3765_ _0465_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_4872_ core_0.decode.i_imm_pass\[11\] _1341_ _1350_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_24_85 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7545__A2 _1742_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_46_138 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6611_ _2936_ _2956_ _2957_ _0224_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__5556__A1 _0982_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7591_ _3682_ _3709_ _3710_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_62_609 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_145_836 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_157_696 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_27_352 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_rebuffer1_I _0548_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_661 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_145_858 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_43_812 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6542_ net128 _2611_ _2906_ _2912_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_131_53 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_144_379 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_131_86 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_160_839 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6473_ _1993_ _2178_ _1457_ _2852_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_8212_ _0388_ clknet_leaf_35_i_clk net84 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_2
XANTENNA__5859__A2 _1197_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_112_232 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5424_ core_0.execute.alu_mul_div.div_cur\[8\] _1812_ _1841_ _1865_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xoutput200 net200 sr_bus_data_o[15] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_140_552 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_8143_ _0319_ clknet_leaf_119_i_clk core_0.execute.rf.reg_outputs\[1\]\[2\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_10_230 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5355_ _1526_ _1527_ _1803_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_2
XANTENNA__4531__A2 _1053_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_10_241 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_167_2519 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_151_Right_151 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_226_100 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4306_ _0888_ _0895_ _0891_ _0924_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or3_1
X_8074_ _0250_ clknet_leaf_100_i_clk core_0.execute.rf.reg_outputs\[6\]\[13\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_2
X_5286_ _0810_ _1734_ _1735_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_4
X_7025_ _2567_ _3181_ _3182_ _3239_ _3209_ _1613_ _0356_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai222_1
X_4237_ _0824_ _0855_ _0856_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4295__A1 core_0.fetch.out_buffer_valid vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_241_103 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_226_177 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4168_ core_0.ew_reg_ie\[7\] _0774_ _0777_ core_0.ew_reg_ie\[6\] _0787_ vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_223_851 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_92 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_241_158 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6036__A2 _2009_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_222_350 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4047__B2 core_0.execute.rf.reg_outputs\[5\]\[4\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
X_4099_ _0713_ _0718_ _0719_ _0720_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_4
XFILLER_0_179_254 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_78_731 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_222_383 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7927_ _0105_ clknet_leaf_0_i_clk core_0.execute.alu_mul_div.cbit\[2\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_2
XANTENNA__5795__A1 _2187_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_65_403 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_77_263 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_178_2648 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_65_414 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7858_ _0050_ clknet_leaf_62_i_clk core_0.fetch.prev_request_pc\[1\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_194_268 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_148_663 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_842 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_93_756 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_175_460 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_191_2804 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6809_ _2992_ _3065_ _3081_ _0298_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_108_516 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_147_162 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5547__A1 net85 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8121__CLK clknet_leaf_99_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_108_527 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_163_622 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_18_341 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_92_255 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7789_ core_0.decode.i_instr_l\[13\] _3786_ _3802_ core_0.decode.i_instr_l\[10\]
+ _1133_ _3856_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_0_18_352 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_190_441 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_135_346 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_135_368 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_151_839 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4770__A2 _1285_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_104_733 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4430__I _0735_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_230_3270 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_33_388 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_591 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7839__CLK clknet_leaf_67_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5970__B _1061_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_103_276 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4522__A2 _1095_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_189_2777 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_218_601 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_103_298 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_111_1839 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_218_645 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_218_667 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_206_807 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__7472__A1 _0553_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_205_317 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7224__A1 net81 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6027__A2 _2414_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4038__A1 core_0.execute.rf.reg_outputs\[6\]\[5\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_204_2958 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_66_1307 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_213_372 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_17_715 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_216_97 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_201_556 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5250__A3 _1452_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_56_403 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_84_723 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_96_594 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7527__A2 _3646_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_122_1979 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_56_447 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_173_419 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_127_836 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_127_858 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_83_277 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_153_121 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_153_132 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4210__A1 _0723_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_4_717 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_142_839 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_52_664 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_141_338 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_77_1436 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_51_185 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_110_725 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5710__A1 _1596_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4513__A2 core_0.decode.i_instr_l\[2\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5140_ core_0.execute.rf.reg_outputs\[1\]\[8\] net218 _1486_ core_0.execute.rf.reg_outputs\[5\]\[8\]
+ core_0.execute.rf.reg_outputs\[6\]\[8\] _1435_ _1589_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_0_20_594 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_244_3439 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_5071_ _1507_ _1512_ _1517_ _1519_ _1520_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_4
XANTENNA__4277__A1 _0892_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_208_166 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_236_486 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_208_177 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4022_ core_0.execute.rf.reg_outputs\[1\]\[6\] _0649_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_0_224_648 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_223_136 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_223_147 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6018__A2 _2300_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_126_53 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_88_1565 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_59_230 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5973_ _1601_ _2361_ _2363_ _1686_ _2364_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_177_758 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_75_712 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7712_ _1382_ _0514_ _3807_ _0475_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4924_ _1195_ _1387_ _1388_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__7518__A2 _3640_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_74_211 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_192_728 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7643_ net206 _3733_ _3752_ _3753_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_145_611 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4855_ _0857_ _1306_ _1340_ _0085_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_191_249 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_801 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_51_72 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_145_644 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_220_Right_220 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
X_7574_ core_0.execute.pc_high_out\[3\] _3688_ _3695_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_2
X_4786_ _1290_ _1297_ _0059_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__4201__A1 _0816_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_145_699 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_173_2589 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6525_ core_0.ew_data\[15\] _1985_ _2903_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4752__A2 _1241_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_70_461 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6456_ _2360_ _2825_ _2833_ _2835_ _2836_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_113_552 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_185 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_30_325 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_3_772 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6886__B _3124_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5407_ core_0.execute.alu_mul_div.div_cur\[6\] _1761_ _1849_ _1850_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_113_585 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4504__A2 _1068_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_246_206 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6387_ _2090_ _2459_ _2767_ _2626_ _2768_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai211_4
XTAP_TAPCELL_ROW_208_3003 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_8126_ _0302_ clknet_leaf_93_i_clk core_0.execute.rf.reg_outputs\[2\]\[1\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_101_769 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_208_3014 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_5338_ _1782_ _1784_ _1785_ _1786_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or3_1
XANTENNA_input41_I i_req_data[12] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7454__A1 _0592_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_50_1108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6257__A2 _1765_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_8057_ _0233_ clknet_leaf_99_i_clk core_0.execute.rf.reg_outputs\[7\]\[12\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__4268__A1 _0723_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5269_ core_0.decode.oc_alu_mode\[12\] _1707_ _1709_ _1717_ _1718_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XFILLER_0_242_412 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_227_486 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7008_ _3214_ _3218_ _3223_ _3224_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_242_434 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_126_2024 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_98_804 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_199_349 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7510__B _1217_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_230_629 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4815__I0 _0865_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_210_375 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4440__A1 core_0.decode.i_instr_l\[6\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_219_3143 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_66_745 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_155_419 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_167_279 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_26_609 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_836 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_182_227 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_661 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_61_1248 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_109_858 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_148_493 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_417 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_277 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_748 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_191_772 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_22_773 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_137_2153 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_80_247 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_34_642 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_18_193 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_124_839 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_190_271 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_123_327 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_34_664 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_34_675 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4160__I _0778_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_174 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6796__B _3072_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_238_718 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_21_369 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7693__B2 _1037_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_237_206 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5192__S _1461_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8017__CLK clknet_leaf_48_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_246_740 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_218_453 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_72_1377 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_206_626 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_148_2293 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_206_659 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_199_861 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_202_865 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4026__A4 core_0.execute.rf.reg_outputs\[6\]\[6\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5223__A3 _0776_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6420__A2 _1501_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_159_769 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_69_583 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_201_375 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_139_460 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_158_279 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_173_216 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_174_739 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_56_244 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_56_255 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_127_622 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_56_277 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_72_737 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_84_597 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_112_33 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4640_ net181 net184 net183 _1199_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or3_2
XANTENNA__6184__A1 _2569_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_72_759 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_7_Left_254 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_25_653 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4571_ _1150_ net157 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__5931__A1 _1689_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_126_187 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_181_282 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5166__I _1608_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_601 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_152 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_547 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_114_349 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6310_ _2576_ _2692_ _2693_ _0187_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_25_686 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_188_37 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_12_314 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7290_ net75 net74 _3454_ _3467_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and3_2
XANTENNA__7133__B1 net214 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_185 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_4_14__f_i_clk clknet_3_7_0_i_clk clknet_4_14__leaf_i_clk vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_97_46 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_667 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6241_ _1693_ _1698_ _1452_ _2626_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_4
XANTENNA__7684__A1 _1044_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_228_228 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6172_ _1559_ net223 _1555_ _2559_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or3_2
XANTENNA__7436__A1 _0626_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5123_ core_0.execute.rf.reg_outputs\[2\]\[10\] _1438_ _1572_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_243_209 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_224_401 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5054_ _1466_ net192 _1503_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4005_ _0517_ _0535_ _0527_ core_0.execute.rf.reg_outputs\[2\]\[8\] _0634_ vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_0_177_500 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_211_139 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_149_202 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_67_509 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_149_235 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4017__A4 core_0.execute.rf.reg_outputs\[2\]\[7\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_94_317 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_47_200 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_165_706 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5956_ core_0.execute.sreg_irq_pc.o_d\[2\] _2264_ _2265_ core_0.execute.alu_flag_reg.o_d\[2\]
+ _2258_ net105 _2347_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_0_177_566 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4422__A1 _0959_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_48_745 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_137_419 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_175_2607 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_48_756 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_62_93 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_175_2618 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_61_i_clk_I clknet_4_14__leaf_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_47_1081 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_47_244 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4907_ _1371_ _1372_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_164_216 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_48_778 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_48_789 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5887_ _0800_ _2279_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_164_238 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4973__A2 _1393_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_164_249 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_47_277 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_35_417 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7626_ _0735_ _3729_ _3740_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6175__A1 _1480_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_145_452 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4838_ _1280_ net42 _1170_ _1329_ _1330_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_7_352 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_62_225 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_145_463 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_173_772 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_62_247 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_117_165 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4725__A2 _1237_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5922__A1 _1553_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_90_578 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_145_496 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7557_ _3673_ _3679_ _3680_ _0447_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_4769_ _1284_ _1288_ _0051_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_133_647 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_31_601 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_675 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_214_3084 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6508_ _1457_ _2873_ _2875_ _1458_ _2885_ _2886_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai221_4
XFILLER_0_132_146 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7488_ core_0.execute.trap_flag _3633_ _3635_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_113_360 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_101_511 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6439_ _1059_ _2814_ _2516_ _2815_ _2818_ _2819_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_0_219_217 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_166 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4489__A1 _1041_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_30_177 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_132_2094 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_101_566 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_186_2747 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5150__A2 net202 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_101_588 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8109_ _0285_ clknet_leaf_96_i_clk core_0.execute.rf.reg_outputs\[3\]\[0\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_228_784 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_242_220 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_227_294 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_199_113 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_242_231 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_199_135 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_98_601 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6650__A2 _2962_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_97_133 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_86_807 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_211_640 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_201_2928 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_27_832 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6938__B1 _1601_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_85_317 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_97_177 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_39_723 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_97_188 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6402__A2 _2279_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_195_352 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4413__A1 net81 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_745 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_531 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_197_2876 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_66_553 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_149_791 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_255 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_715 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_277 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_136_430 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_737 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_597 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_214 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_81_556 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5913__A1 _1554_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_53_269 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_151_422 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_163_282 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4716__A2 _1253_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_601 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_198 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_123_135 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_472 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_124_669 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_151_477 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_74_1406 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_21_133 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_10_807 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_22_667 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7666__A1 _1414_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_104_382 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7666__B2 _3767_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7418__A1 net215 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_246_570 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_241_3409 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_206_401 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_233_231 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_83_37 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6641__A2 _2981_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4652__A1 _1197_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_50_i_clk clknet_4_12__leaf_i_clk clknet_leaf_50_i_clk vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_16_53 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_85_1535 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_187_842 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_186_330 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_76_317 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_88_177 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_202_662 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5810_ _2201_ _2209_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_201_150 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6790_ _2961_ _3064_ _3071_ _0289_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__4404__A1 _0836_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_9_628 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5741_ _1471_ _1475_ _2141_ _2142_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XANTENNA__4955__A2 _0637_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_45_704 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_29_255 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xclkbuf_leaf_65_i_clk clknet_4_15__leaf_i_clk clknet_leaf_65_i_clk vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_225_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__7376__I _3542_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_45_726 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_737 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6157__A1 _2244_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_32_85 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5672_ _1702_ _1491_ _2073_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_155_772 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7411_ _1357_ _1008_ _3546_ _3572_ _3573_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_44_247 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_115_636 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4623_ _1175_ core_0.execute.alu_flag_reg.o_d\[2\] _1180_ _1176_ _1182_ vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai22_1
XANTENNA__5904__A1 _2294_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_72_578 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_142_422 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_170_731 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_182_591 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_115_669 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_170_2548 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_7342_ _3510_ _3512_ _3513_ _0399_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_4554_ _1131_ _1134_ _1135_ _1136_ _0006_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_0_52_291 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_96_1664 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_142_488 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_13_656 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_130_639 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_111_820 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7273_ _3447_ _3448_ _3452_ _0391_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_13_678 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_111_842 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4485_ core_0.decode.i_instr_l\[6\] _1047_ core_0.decode.i_instr_l\[5\] _1078_ vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_0_229_537 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_486 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_177 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6224_ core_0.execute.alu_mul_div.div_cur\[7\] _1117_ _2610_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5132__A2 core_0.execute.rf.reg_outputs\[4\]\[9\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_244_507 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7409__A1 _3543_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6155_ _2403_ _2456_ _2495_ _2541_ _2542_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or4_1
XANTENNA__6880__A2 _3108_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4891__A1 _0726_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5106_ _1542_ _1550_ _1554_ _1555_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_6086_ core_0.decode.oc_alu_mode\[11\] _2466_ _2467_ _2471_ _2474_ _2475_ vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_0_32_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5037_ _0782_ _0767_ _0775_ _1486_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_4
Xclkbuf_leaf_18_i_clk clknet_4_8__leaf_i_clk clknet_leaf_18_i_clk vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__4643__A1 _1196_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_181_2688 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_224_286 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_224_297 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_68_807 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_196_127 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_73_92 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_24_802 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5199__A2 _0768_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_177_352 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6988_ _3203_ _3205_ _3206_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_138_728 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_105_1771 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_165_525 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_216_3102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4946__A2 net205 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5939_ core_0.execute.alu_mul_div.div_res\[1\] _2331_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_0_35_203 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6190__I _2201_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_737 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6148__A1 core_0.execute.pc_high_buff_out\[6\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_35_225 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6148__B2 net13 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_90_331 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_35_247 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_63_556 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_192_399 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_7_160 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output195_I net195 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7609_ _3676_ _3724_ _3725_ _3726_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__6699__A2 _3000_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_145_282 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_134_2123 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_90_375 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_105_146 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_121_617 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_43_291 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_133_488 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7235__B _1395_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7648__A1 core_0.execute.pc_high_buff_out\[7\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_31_486 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5123__A2 _1438_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6320__A1 _2287_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_79_Left_326 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_101_352 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_output72_I net72 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6320__B2 _1690_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_101_363 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_227_3231 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_101_374 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput77 net77 dbg_pc[14] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XTAP_TAPCELL_ROW_227_3242 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
Xoutput88 net88 dbg_r0[0] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_207_209 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6566__S _2201_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput99 net99 dbg_r0[5] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA__6871__A2 _3114_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_228_592 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_216_754 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_231_702 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_145_2252 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4229__A4 _0847_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6623__A2 _2962_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_4_560 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_208_87 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_203_415 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_199_2905 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_188_628 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_98_431 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_169_831 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_169_842 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_230_256 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_58_317 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_129_706 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6387__A1 _2090_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8205__CLK clknet_leaf_2_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_88_Left_335 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_129_739 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_224_86 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_211_492 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_224_97 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_238_3371 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_144_709 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_39_597 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6139__A1 _2360_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_109_452 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_80_1476 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_137_772 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_26_247 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_82_865 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_156_2381 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_41_206 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_152_742 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_112_617 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5362__A2 _0801_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_78_37 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7639__A1 net227 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_97_Left_344 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_111_138 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_637 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4270_ core_0.fetch.prev_request_pc\[12\] _0823_ _0854_ core_0.fetch.prev_request_pc\[11\]
+ _0888_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai22_1
XANTENNA__4173__I0 core_0.ew_reg_ie\[4\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6862__A2 _3108_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_207_710 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4873__A1 _0854_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_118_43 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3899__I _0523_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_118_54 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_175_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__7811__A1 _1034_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_74 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7960_ _0138_ clknet_leaf_1_i_clk core_0.execute.alu_mul_div.div_cur\[0\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_221_212 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_85 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_179_628 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6911_ net102 _3135_ _3139_ _3141_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_178_138 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3979__A3 _0549_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7891_ _0082_ clknet_leaf_82_i_clk core_0.decode.i_imm_pass\[0\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_175_801 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_221_289 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6842_ core_0.execute.rf.reg_outputs\[2\]\[11\] _3092_ _3098_ _3101_ vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_159_352 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_76_136 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_147_514 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_175_823 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_202_492 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_187_694 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_134_97 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_76_169 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6773_ core_0.execute.rf.reg_outputs\[4\]\[14\] _3041_ _3057_ _3061_ vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3985_ _0615_ net195 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_186_193 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_190_804 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_44_1040 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_18_737 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5724_ _1819_ _2124_ _2125_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_45_556 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_127_260 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_17_258 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_353 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_198_Right_198 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_45_578 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5655_ _1508_ _1509_ _2053_ _2056_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_4
XFILLER_0_115_422 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_515 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_642 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4606_ net17 net160 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_32_239 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5586_ _1521_ _1522_ _1987_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_2
XTAP_TAPCELL_ROW_211_3043 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_7325_ _2711_ _2734_ _2746_ _3498_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_142_285 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4561__B1 _1064_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4537_ _1034_ _1120_ _1122_ _0001_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_159_50 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7256_ _3384_ _3437_ _3438_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6302__A1 _2281_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4468_ core_0.decode.oc_alu_mode\[7\] _1061_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_40_294 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6207_ core_0.decode.oc_alu_mode\[11\] _2592_ _2593_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_183_2706 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_7187_ _1748_ _3378_ _0379_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_244_326 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4399_ _1004_ _0966_ _1006_ _1007_ _0877_ net173 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_0_244_337 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4864__A1 _0833_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6138_ _1117_ _2524_ _2525_ _2526_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_4
XFILLER_0_99_206 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_225_562 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_213_702 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6605__A2 _2951_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6069_ _2244_ _2455_ _2457_ _2458_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
XTAP_TAPCELL_ROW_107_1800 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_222_3172 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_1_530 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_169_127 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4092__A2 _0594_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_37_960 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output208_I net208 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6369__A1 core_0.execute.alu_mul_div.div_cur\[11\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_95_456 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7030__A2 _1637_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_140_2193 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6464__S1 _2123_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_194_2835 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_83_629 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_95_489 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4919__A2 _1382_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5529__I _1955_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_194_2846 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4433__I _0745_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_76_692 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_119_750 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_82_139 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_181_815 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_192_163 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5592__A2 net214 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_64_865 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_118_271 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_181_859 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_134_731 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_180_336 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_EDGE_ROW_165_Right_165 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_90_172 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_51_537 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_51_548 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_58_1209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_210_77 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7097__A2 _3285_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_208_518 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6844__A2 _3092_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_101_193 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4855__A1 _0857_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6057__B1 _2260_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5213__B _1483_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_188_403 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_203_212 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4607__A1 core_0.decode.i_flush vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_69_1338 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6998__I3 _1665_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_86_401 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4083__A2 _0529_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_626 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5280__A1 _1432_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_157_812 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_58_158 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_156_311 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_157_834 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_168_171 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_46_309 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_86_478 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_158_2410 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_129_558 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_156_333 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_168_193 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_156_344 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_172_804 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_73_139 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_156_366 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_172_815 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7309__B1 _3399_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_15_687 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6780__A1 core_0.execute.rf.reg_outputs\[3\]\[0\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_15_698 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_144_539 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_156_399 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_172_859 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_109_282 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_EDGE_ROW_132_Right_132 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_89_47 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5440_ _1790_ _1788_ _1878_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_120_33 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_89_69 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5335__A2 _1756_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_23_751 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_124_285 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xclkbuf_4_2__f_i_clk clknet_3_1_0_i_clk clknet_4_2__leaf_i_clk vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_5371_ _1554_ _1819_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XTAP_TAPCELL_ROW_93_1623 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_50_570 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_93_1634 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_120_99 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_239_632 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7110_ _2778_ _3181_ _3318_ _0362_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_2_667 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4322_ _0868_ _0940_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__inv_1
X_8090_ _0266_ clknet_leaf_100_i_clk core_0.execute.rf.reg_outputs\[5\]\[13\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_196_59 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7041_ _3149_ _3253_ _3254_ _3255_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_4253_ _0820_ _0871_ _0872_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__6835__A2 _3092_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5902__I _2293_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4846__A1 _1280_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_226_348 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_129_86 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4184_ core_0.decode.o_submit core_0.execute.alu_mul_div.i_mul _0803_ vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_38_95 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_207_562 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6599__A1 _2936_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_222_521 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_234_381 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7943_ _0121_ clknet_leaf_42_i_clk core_0.execute.sreg_priv_control.o_d\[15\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_77_401 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5271__A1 core_0.decode.oc_alu_mode\[12\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_103 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_194_417 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_210_749 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7874_ _0065_ clknet_leaf_71_i_clk core_0.fetch.out_buffer_data_pred vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_166_119 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_200 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6825_ _2956_ _3086_ _3091_ _0304_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_147_322 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_77_489 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_102_1741 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_58_681 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_175_664 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_175_675 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_320 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5574__A2 _0745_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6756_ core_0.execute.rf.reg_outputs\[4\]\[6\] _3049_ _3045_ _3052_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_9_277 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3968_ _0533_ _0541_ _0543_ core_0.execute.rf.reg_outputs\[5\]\[11\] _0600_ vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_0_161_84 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_865 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_70_82 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_162_314 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_45_364 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5707_ _1123_ _1652_ net211 _2092_ _2108_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_0_128_591 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6687_ core_0.execute.rf.reg_outputs\[6\]\[9\] _3006_ _3004_ _3012_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3899_ _0523_ _0535_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_45_386 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_312 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_559 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5638_ _2036_ _2038_ _2039_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__5326__A2 _1765_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_103_403 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_115_263 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input71_I i_rst vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_60_367 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4534__B1 _1094_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_170_391 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5569_ _1419_ _0735_ _0160_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_130_244 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7308_ net77 net76 _3467_ _3483_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_2
X_8288_ _0464_ clknet_leaf_48_i_clk core_0.dec_mem_long vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_229_142 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_218_827 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__7513__B _3651_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6908__I _0722_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_113_1870 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output158_I net158 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7239_ net83 _3422_ _3423_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_224_3201 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4837__A1 _1280_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_217_348 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_129_2055 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_129_2066 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4428__I _0739_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_244_189 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_142_2211 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7787__B1 _3827_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_198_734 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_142_2222 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7251__A2 _3391_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_87_209 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_197_233 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_96_710 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_234_Right_234 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__6643__I _1963_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_185_417 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_200_237 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_95_242 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_178_491 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_205_88 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_489 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_96_798 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5014__A1 _0568_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_165_130 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_64_1279 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_235_3330 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_193_472 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6762__A1 core_0.execute.rf.reg_outputs\[4\]\[9\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5565__A2 _1955_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_48_191 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_153_314 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_107_720 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4773__B1 _0881_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_107_731 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_150 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_181_656 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_12_657 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_51_301 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_40_988 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_3_409 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_180_155 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_91_492 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_181_689 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5317__A2 net187 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6514__A1 _2891_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_153_2351 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_180_177 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_180_188 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_134_583 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_121_244 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_32_581 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_732 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7423__B _3553_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_209_838 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5722__I _2102_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4828__A1 core_0.decode.i_instr_l\[11\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_246_3470 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_246_3481 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_246_40 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_217_860 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_164_2480 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7242__A2 _3421_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_188_233 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4056__A2 _0530_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5253__A1 _1528_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_188_244 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_188_255 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_201_Right_201 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
X_4940_ core_0.execute.sreg_long_ptr_en _1394_ _1401_ _1391_ _1402_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_176_417 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87_765 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_188_299 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_47_618 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_129_333 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4871_ _1348_ _1321_ _1349_ _0092_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_59_489 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5005__A1 core_0.decode.oc_alu_mode\[1\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_138_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6610_ core_0.execute.rf.reg_outputs\[7\]\[3\] _2941_ _1978_ _2957_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_200_793 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7590_ core_0.execute.pc_high_out\[5\] _3702_ _3709_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_28_843 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5556__A2 _1956_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6753__A1 _2961_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_41_1010 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_28_865 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_144_314 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_156_174 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5800__I0 net132 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_156_185 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6541_ _2911_ _0200_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4764__B1 _0881_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_42_301 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_160_807 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_54_172 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4801__I _1305_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6505__A1 _2133_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6472_ _2841_ _2844_ _2849_ _2850_ _2851_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XFILLER_0_40_85 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8211_ _0387_ clknet_leaf_31_i_clk net83 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_2
X_5423_ core_0.execute.alu_mul_div.div_cur\[7\] _1814_ _1863_ _1864_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_140_531 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput201 net201 sr_bus_data_o[1] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_23_570 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_112_244 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_2_453 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8073__CLK clknet_leaf_99_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_112_255 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_11_743 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8142_ _0318_ clknet_leaf_117_i_clk core_0.execute.rf.reg_outputs\[1\]\[1\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5354_ _1797_ _1799_ _1801_ _1802_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_140_597 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_497 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_100_439 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4305_ core_0.fetch.prev_request_pc\[7\] _0833_ _0923_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__6808__A2 _3070_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_8073_ _0249_ clknet_leaf_99_i_clk core_0.execute.rf.reg_outputs\[6\]\[12\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5285_ _1195_ _1203_ _1733_ _1734_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_4
XFILLER_0_10_286 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7024_ _2567_ _3237_ _3238_ _3239_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_4236_ core_0.fetch.out_buffer_data_instr\[19\] _0855_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__7481__A2 _1398_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_241_115 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_65_60 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4167_ _0772_ _0780_ _0784_ _0785_ _0786_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XFILLER_0_223_830 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_207_381 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7769__B1 _3833_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_97_518 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_223_863 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4098_ net88 _0521_ _0719_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or2_2
XFILLER_0_179_233 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7559__I _3681_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4047__A2 _0661_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7926_ _0104_ clknet_leaf_0_i_clk core_0.execute.alu_mul_div.cbit\[1\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_77_220 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_179_277 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5795__A2 _2194_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_194_214 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6992__A1 _1665_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_77_242 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_167_439 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_194_236 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_178_2649 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_7857_ _0049_ clknet_leaf_61_i_clk core_0.fetch.prev_request_pc\[0\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_4
XFILLER_0_194_247 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_77_275 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_147_130 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_92_223 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_148_675 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_37_139 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6808_ core_0.execute.rf.reg_outputs\[3\]\[13\] _3070_ _3072_ _3081_ vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_191_2805 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_93_768 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5547__A2 _1953_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7788_ _1136_ _3855_ _0503_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_80_407 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_147_196 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6739_ core_0.ew_reg_ie\[4\] _2934_ _3041_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_0_190_453 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_162_155 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_61_632 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_492 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_150_317 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_162_177 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6131__C _2412_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_356 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_153 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_61_676 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_230_3271 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_60_186 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_197_80 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_189_2778 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_218_613 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_52_Left_299 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA_clkbuf_leaf_56_i_clk_I clknet_4_11__leaf_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_245_443 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7472__A2 _3546_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5483__A1 _1909_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_232_104 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_232_115 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6574__S _2201_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3997__I _0626_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4038__A2 _0661_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_66_1308 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_204_2959 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_216_76 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_17_716 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_198_586 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_240_181 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_198_597 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_186_737 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6983__A1 _3183_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_242 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_787 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_629 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_185_269 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_28_117 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_83_212 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_166_450 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_139_675 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_166_461 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_232_53 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_153_100 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_138_185 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_166_494 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7418__B _3545_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_193_291 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5943__C1 _2258_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_52_610 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_142_807 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_154_667 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_92_790 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8096__CLK clknet_leaf_94_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_181_486 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_24_345 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_356 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_51_142 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_52_676 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_134_380 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_77_1437 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7160__A1 _1369_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_51_197 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5710__A2 _1481_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_110_737 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_122_597 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_86_37 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_208_101 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_20_584 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_208_134 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5070_ _1461_ net205 _1518_ _1519_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_0_224_616 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4277__A2 _0837_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4021_ net216 net207 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_223_115 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_205_830 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_189_531 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6018__A3 _1624_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_518 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4029__A2 _0523_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_88_1566 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7379__I _3540_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_220_811 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_149_406 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_189_586 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5972_ _1059_ _2362_ _2000_ _2363_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_87_540 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_75_702 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_87_562 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7711_ core_0.decode.i_imm_pass\[0\] _1064_ _3807_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_176_247 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4923_ _1209_ core_0.execute.sreg_priv_control.o_d\[0\] _1386_ _1387_ vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_118_804 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4732__S _1246_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_145_601 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7642_ _0745_ _3729_ _3752_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_74_234 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6726__A1 _2983_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4854_ core_0.decode.i_imm_pass\[3\] _1307_ _1340_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_145_623 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_191_239 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_74_267 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4588__I0 core_0.ew_data\[0\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_117_347 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4785_ core_0.fetch.prev_request_pc\[10\] net225 _0880_ net162 _1297_ vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_0_7_556 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7573_ _3673_ _3693_ _3694_ _1950_ _0449_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_172_453 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_790 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_55_492 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_132_317 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6524_ _0553_ _2901_ _2241_ _2902_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_144_177 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_43_676 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_142 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_144_199 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_153 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_99_1695 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_125_380 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_3_740 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6455_ _2356_ _2834_ _2835_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__7151__A1 _1838_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5406_ _1777_ _1778_ _1849_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_6386_ _2089_ _2766_ _2767_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_30_359 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_113_597 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_294 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_208_3004 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_8125_ _0301_ clknet_leaf_92_i_clk core_0.execute.rf.reg_outputs\[2\]\[0\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_2
X_5337_ core_0.execute.alu_mul_div.div_cur\[9\] _1754_ _1785_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_100_247 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_11_595 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_50_1109 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_167_72 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__7454__A2 _3546_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_8056_ _0232_ clknet_leaf_104_i_clk core_0.execute.rf.reg_outputs\[7\]\[11\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5268_ _1710_ _1711_ _1713_ _1716_ _1717_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_4
XANTENNA_input34_I i_mem_data[7] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4268__A2 net61 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5465__A1 _1232_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_215_627 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4219_ net52 core_0.fetch.out_buffer_data_instr\[22\] _0724_ _0838_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_214_104 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_199_306 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7007_ core_0.execute.alu_mul_div.mul_res\[4\] _3217_ _3223_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_126_2025 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_5199_ _0782_ _0768_ _1646_ _1647_ _1648_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai31_2
XANTENNA__7206__A2 _1195_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_211_800 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5217__A1 _0771_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6193__I _2254_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6965__A1 _3183_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4815__I1 core_0.decode.i_instr_l\[6\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7909_ _0100_ clknet_leaf_52_i_clk core_0.fetch.pc_flush_override vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_195_578 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4440__A2 core_0.decode.i_instr_l\[4\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_155_409 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_183_718 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_219_3144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_210_387 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_38_448 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6717__A1 _2967_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_65_245 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_256 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6568__I1 core_0.ew_reg_ie\[4\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_232_3300 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_61_1249 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_93_576 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_136_645 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_202_34 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_19_684 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_18_150 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_738 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_108_358 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_124_807 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__7390__A1 _1357_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_137_2154 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_22_774 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_80_237 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_151_615 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_163_475 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_202_89 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_33_142 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_150_2310 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_21_315 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_131_361 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_60_Left_307 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_131_383 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_218_421 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_72_1378 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_246_774 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_245_262 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_148_2283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_148_2294 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_221_619 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5208__A1 _0782_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_161_2450 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_220_107 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5221__B _0769_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_243_41 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6036__C _1059_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_551 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_702 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_69_562 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_159_759 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_158_247 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_84_510 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_69_595 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6708__A1 _2946_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_139_472 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_72_705 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_37_492 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_25_632 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_126_155 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4570_ _1149_ _1150_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_114_317 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_182_795 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6987__B _2436_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5931__A2 _1652_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_52_451 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_21_98 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_97_14 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_141_136 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_52_473 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_25_698 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7133__A1 _3149_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7133__B2 _3209_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_12_326 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6240_ _2356_ _2624_ _2625_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_97_58 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_97_69 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_228_207 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6171_ _1613_ _2555_ _2557_ _2558_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5122_ _1569_ _1570_ _1571_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__7436__A2 _3544_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8111__CLK clknet_leaf_109_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5447__A1 core_0.execute.alu_mul_div.div_cur\[11\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_224_424 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5053_ _1482_ _1501_ _1502_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_46_51 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_224_457 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4004_ _0565_ _0541_ _0543_ core_0.execute.rf.reg_outputs\[5\]\[8\] _0633_ vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_4
XPHY_EDGE_ROW_108_Left_355 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_137_97 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_79_315 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_79_337 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4526__I _0798_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6947__A1 _1231_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_153_52 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5955_ core_0.dec_mem_access _2346_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_47_212 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_175_2608 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_87_392 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6741__I _3041_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_153_96 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_47_1071 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_4906_ _1222_ _1371_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_0_75_543 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_47_1082 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_5886_ core_0.ew_data\[1\] _2209_ _2278_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7625_ _3732_ _3738_ _3739_ _0456_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_7_342 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_865 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_106_807 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4837_ _1280_ _1257_ _1329_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_EDGE_ROW_117_Left_364 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
X_7556_ core_0.execute.pc_high_out\[0\] _3673_ _1216_ _3680_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4768_ core_0.fetch.prev_request_pc\[2\] _1285_ _0881_ net169 _1288_ vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai22_1
XANTENNA__5922__A2 _2019_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6897__B _3124_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_15_142 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_214_3085 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_43_473 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6507_ _2877_ _2878_ _2884_ _2885_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and3_1
XANTENNA__7124__A1 _3175_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4699_ _1247_ _0022_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7487_ _1217_ _1207_ _3634_ _0423_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_15_197 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_31_668 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6438_ _1994_ _2816_ _2817_ _2818_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA__7675__A2 _3766_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5686__A1 _1711_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4489__A2 _1056_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_132_2095 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5092__I net214 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_186_2748 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6369_ core_0.execute.alu_mul_div.div_cur\[11\] _1117_ _2751_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_8108_ _0284_ clknet_leaf_96_i_clk core_0.execute.rf.reg_outputs\[4\]\[15\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5438__A1 core_0.execute.alu_mul_div.div_cur\[10\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7521__B _3651_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_126_Left_373 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
X_8039_ _0216_ clknet_leaf_81_i_clk core_0.ew_reg_ie\[6\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_215_457 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_199_125 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_194_81 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7240__C _1735_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_98_613 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_202_107 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6938__A1 _1231_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_201_2929 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_27_833 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6938__B2 _1926_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_85_307 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_702 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4413__A2 _0883_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_195_364 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5610__A1 _1695_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_197_2877 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_39_757 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_543 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_94_863 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_623 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_155_228 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_213_66 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_183_559 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_135_Left_382 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_19_481 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_492 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_151_401 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_259 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_177 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5913__A2 _1501_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3924__A1 _0539_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7115__A1 _1364_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_635 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_111_309 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_292 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_151_489 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7666__A2 _3766_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_238_527 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_120_865 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_219_741 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_219_752 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_219_763 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7418__A2 _3544_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_144_Left_391 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__5429__A1 _1232_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_234_733 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_206_424 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_7_591 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8284__CLK clknet_leaf_29_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_233_265 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6047__B _0798_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_88_101 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_221_416 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4652__A2 _1199_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_202_630 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_199_692 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_16_65 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6929__A1 _1915_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_85_1536 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_88_156 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_EDGE_ROW_179_Right_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_16_98 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4404__A2 _0947_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_29_212 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5601__A1 _2001_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5740_ _1551_ _1552_ _2140_ _1449_ _2141_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_0_57_554 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_146_228 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7729__I0 net193 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_32_53 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_123_66 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_84_373 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5671_ _1528_ _1529_ _1994_ _2072_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_0_120_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_161_209 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_218_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_44_237 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7410_ _1357_ core_0.execute.mem_stage_pc\[5\] _3572_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4168__A1 core_0.ew_reg_ie\[7\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_142_401 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4168__B2 core_0.ew_reg_ie\[6\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4622_ core_0.dec_jump_cond_code\[1\] core_0.dec_jump_cond_code\[0\] _1181_ vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_154_272 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_127_497 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_451 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5904__A2 _2295_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_115_648 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3915__A1 _0534_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_170_2549 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_7341_ core_0.execute.alu_flag_reg.o_d\[1\] _3510_ _3139_ _3513_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4553_ _1051_ _1136_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_4_356 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_12_101 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_114_158 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_80_590 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_96_1665 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_7272_ _3384_ _3451_ _3452_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_40_454 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4484_ _1070_ _1076_ _1077_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_6223_ core_0.execute.alu_mul_div.div_res\[7\] _2332_ _2279_ _2609_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_40_498 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_690 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4340__A1 core_0.fetch.prev_request_pc\[15\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6154_ _2540_ _2541_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_57_72 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7341__B _3139_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5105_ _1553_ _1554_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
X_6085_ _1690_ _2013_ _2472_ _1929_ _2473_ _2474_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_0_224_221 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_225_766 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6093__A1 _1117_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5036_ core_0.execute.rf.reg_outputs\[2\]\[13\] _1438_ _1443_ core_0.execute.rf.reg_outputs\[3\]\[13\]
+ net218 core_0.execute.rf.reg_outputs\[1\]\[13\] _1485_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_0_225_788 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_25_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_197_629 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_49_1100 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5840__A1 net137 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_181_2689 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_212_449 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_240_769 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_95_627 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_177_331 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_146_Right_146 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__7593__A1 net205 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6987_ _1222_ _3204_ _2436_ _3205_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_24_803 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6396__A2 _2768_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_88_690 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_105_1772 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_192_312 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_543 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5938_ _2281_ _2328_ _2329_ _2330_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_76_863 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_137_228 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_216_3103 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_192_323 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6148__A2 _2249_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_118_453 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5869_ _2251_ _1382_ _1197_ _2262_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_0_8_662 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4159__A1 core_0.dec_l_reg_sel\[1\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7608_ core_0.execute.pc_high_buff_out\[7\] _3676_ _3725_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_90_343 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_32_891 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_63_568 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_44_760 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_50_207 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_134_2124 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_145_294 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_659 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_387 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output188_I net188 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7539_ core_0.execute.sreg_irq_flags.o_d\[2\] _1398_ core_0.execute.sreg_irq_flags.i_d\[2\]
+ _3666_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_161_787 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_432 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_121_629 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5108__B1 _0703_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7648__A2 _3732_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_114_681 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_113_180 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_102_865 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput78 net78 dbg_pc[15] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XTAP_TAPCELL_ROW_227_3232 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
Xoutput89 net89 dbg_r0[10] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA__4882__A2 _1136_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_243_541 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6084__A1 _1061_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6084__B2 _1109_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_4_561 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_145_2253 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_231_714 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7820__A2 _1032_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_231_725 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_199_2906 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_187_139 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_58_329 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_830 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_113_Right_113 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_85_137 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_195_150 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_39_532 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4398__A1 _0838_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_195_172 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_340 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_183_323 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_238_3372 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_183_334 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_109_431 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_66_384 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6139__A2 _2526_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_54_535 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_80_1477 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_26_237 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_82_855 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_109_497 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_156_2382 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5898__A1 _2286_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_81_376 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5898__B2 _1686_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3954__B _0520_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_151_253 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_169_18 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_590 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_670 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_681 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_239_836 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_239_858 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_10_649 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4173__I1 core_0.ew_reg_ie\[5\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_94_37 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4873__A2 _1321_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7161__B _3357_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_246_390 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6075__A1 core_0.decode.oc_alu_mode\[4\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_206_243 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_168_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_206_298 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6910_ _2977_ _3129_ _3140_ _0340_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_7890_ _0081_ clknet_leaf_77_i_clk core_0.decode.i_instr_l\[15\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_77_627 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_89_487 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_159_331 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_221_279 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6841_ _2986_ _3087_ _3100_ _0311_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_187_662 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7575__A1 core_0.execute.pc_high_out\[3\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7387__I _3540_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_119_206 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4389__A1 _0996_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_186_172 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_863 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6772_ _2992_ _3043_ _3060_ _0282_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_119_228 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3984_ _0608_ _0613_ _0614_ _0615_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_0_147_559 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_44_1041 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_5723_ _1124_ _1491_ _2091_ _2092_ _2124_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai211_2
XANTENNA__7327__A1 _2477_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_395 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_134_209 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4740__S _1246_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5654_ _2052_ _2054_ _2055_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_5_632 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_150_75 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_60_527 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_387 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4605_ _1167_ core_0.ew_mem_width net158 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_142_242 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_60_549 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5585_ _1986_ _0168_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_211_3044 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_103_629 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_130_404 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_5_698 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_130_415 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7324_ _2821_ _3497_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__4561__A1 _1137_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_4_186 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4536_ _1121_ _1053_ _1122_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_40_251 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_111_640 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_229_335 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7255_ net85 _3435_ _3436_ _3437_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_7_74 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6302__A2 _2684_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4467_ _1034_ _1058_ _1060_ _0009_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_111_662 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_111_673 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4313__A1 core_0.fetch.prev_request_pc\[0\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6206_ _2031_ _2021_ _2553_ _2592_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
XTAP_TAPCELL_ROW_183_2707 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_4398_ _0838_ _0947_ _0970_ _1007_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XTAP_TAPCELL_ROW_55_1170 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_7186_ _3365_ _3372_ core_0.execute.alu_mul_div.div_res\[12\] _3378_ vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XPHY_EDGE_ROW_215_Right_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__4864__A2 _1321_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6137_ core_0.execute.alu_mul_div.div_cur\[5\] _1432_ _2525_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_175_72 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_240_500 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6068_ _2403_ _2456_ _2457_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_175_83 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_240_522 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_107_1801 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_197_415 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_1_520 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_240_533 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_222_3173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_5019_ net88 _0521_ _1468_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_169_139 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_200_419 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_68_638 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_37_961 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_95_424 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7566__A1 core_0.execute.pc_high_out\[2\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6369__A2 _1117_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_138_504 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_166_813 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output103_I net103 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_140_2194 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_193_632 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4919__A3 _1197_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_194_2836 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_82_107 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_192_131 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_193_665 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_36_513 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_193_676 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7318__A1 _3409_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_48_395 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_119_762 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_125_209 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_193_687 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_64_855 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_106_401 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5973__C _1686_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_146_581 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_118_283 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_133_220 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_134_765 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_118_1930 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_133_242 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_161_551 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_210_34 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_161_562 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_44_590 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4552__A1 _1037_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_9_620 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_126_i_clk_I clknet_4_1__leaf_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_102_695 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_236_839 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xclkbuf_leaf_64_i_clk clknet_4_15__leaf_i_clk clknet_leaf_64_i_clk vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__4855__A2 _1306_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6057__A1 core_0.execute.sreg_irq_flags.o_d\[4\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6057__B2 net11 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5804__A1 _1987_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_69_1339 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4825__S _1305_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_763 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5280__A2 core_0.execute.alu_mul_div.div_cur\[0\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_79_i_clk clknet_4_13__leaf_i_clk clknet_leaf_79_i_clk vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_58_104 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8322__CLK clknet_leaf_83_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7557__A1 _3673_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_196_470 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_86_457 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_158_2411 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_169_695 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_157_846 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5032__A2 _1469_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_384 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_54_310 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_156_356 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_183_142 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7309__A1 net77 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_13_66 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6780__A2 _3065_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_156_378 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_15_688 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_82_641 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_13_88 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4791__A1 core_0.fetch.prev_request_pc\[13\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_137_592 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_89_26 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_42_527 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_218 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_54_387 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_124_242 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_124_253 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_152_573 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_613 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_112_415 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_17_i_clk clknet_4_8__leaf_i_clk clknet_leaf_17_i_clk vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_112_426 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4543__A1 _1037_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5370_ core_0.execute.alu_mul_div.div_cur\[1\] _1603_ _1769_ _1818_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_22_251 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_93_1624 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_10_413 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4321_ _0935_ _0936_ _0937_ _0938_ _0939_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor4_4
XTAP_TAPCELL_ROW_169_2540 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6296__A1 _1109_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4252_ _0869_ _0870_ _0871_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7040_ _3243_ _3252_ _3254_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__6296__B2 core_0.decode.oc_alu_mode\[6\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_227_839 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4846__A2 net44 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5404__B _1816_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4183_ core_0.decode.o_submit _0801_ _0802_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_38_85 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6048__A1 core_0.execute.alu_mul_div.div_res\[3\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6599__A2 _2946_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_222_533 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7942_ _0120_ clknet_leaf_43_i_clk core_0.execute.sreg_priv_control.o_d\[14\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5271__A2 _1719_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4074__A3 _0548_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_89_262 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_210_728 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7548__A1 _1955_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_148_802 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7873_ core_0.fetch.submitable clknet_leaf_50_i_clk core_0.decode.i_submit vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_194_429 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_49_137 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_187_470 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_34_920 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6824_ core_0.execute.rf.reg_outputs\[2\]\[3\] _3087_ _3083_ _3091_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_187_492 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_65_619 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_175_632 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_92_405 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6220__A1 _1107_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_64_107 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_102_1731 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_102_1742 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6755_ _2967_ _3042_ _3051_ _0274_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_3967_ _0517_ core_0.execute.rf.reg_outputs\[3\]\[11\] net231 _0599_ vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_0_18_535 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_181 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_175_687 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_46_855 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6771__A2 _3049_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_175_698 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4782__A1 _1290_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5706_ _1123_ _1676_ net211 _1720_ _2107_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_0_174_197 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6686_ _2981_ _2999_ _3011_ _0245_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_61_814 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_92_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_3898_ _0533_ _0534_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_45_398 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5637_ _2037_ _1592_ _2038_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_131_702 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_60_335 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_61_858 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_115_275 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_116_798 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_130_201 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_484 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4534__A1 _1084_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4534__B2 _1039_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5568_ _1419_ _0736_ _0159_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_131_757 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_input64_I i_req_data[4] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7307_ net76 _3467_ _3482_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_41_582 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4519_ _1034_ _1106_ _1108_ _0007_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_8287_ _0463_ clknet_leaf_47_i_clk core_0.decode.input_valid vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__dffq_2
X_5499_ _1908_ _1931_ _1932_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6287__A1 _2090_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_130_289 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7238_ _1742_ _3413_ _3422_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_113_1871 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4298__B1 _0860_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_224_3202 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_229_198 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4709__I _1236_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_233_809 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7169_ _3358_ _3367_ core_0.execute.alu_mul_div.div_res\[5\] _3368_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_129_2056 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_226_861 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_232_308 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_213_500 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_142_2212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_198_724 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_241_842 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_197_212 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_240_352 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_206_2990 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5262__A2 _1522_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_205_34 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_68_457 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_138_312 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6211__A1 _1831_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5014__A2 core_0.execute.rf.reg_outputs\[3\]\[0\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_52_i_clk_I clknet_4_14__leaf_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_235_3331 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_83_438 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_165_142 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_166_676 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6762__A2 _3049_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_138_378 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_165_164 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_193_484 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_107_710 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_165_175 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_180_101 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_52_803 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4773__B2 net171 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_365 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_180_123 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_12_658 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_221_66 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_24_527 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_40_989 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_63_184 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_134_551 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_153_2352 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6514__A2 _0798_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7711__A1 core_0.decode.i_imm_pass\[0\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_18 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4525__A1 core_0.decode.i_instr_l\[3\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_121_212 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_106_297 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_593 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7704__B _3799_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6278__A1 _1379_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_246_3460 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_208_327 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4828__A2 _1321_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_246_3471 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_246_3482 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_235_157 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_246_74 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_244_691 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_216_382 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_204_522 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_188_201 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_164_2481 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_231_352 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6450__A1 net76 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5253__A2 _1529_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6450__B2 _2537_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_582 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_231_374 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_115_34 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_86_243 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87_777 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_405 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_157_632 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_169_492 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4870_ core_0.decode.i_imm_pass\[10\] _1341_ _1349_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_46_107 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_200_761 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_28_811 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_24_87 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6202__A1 _1088_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5005__A2 core_0.decode.oc_alu_mode\[6\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_129_356 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_184_440 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_200_783 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_156_142 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6753__A2 _3042_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_41_1000 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5800__I1 _2199_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6540_ net127 _2571_ _2906_ _2911_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__4764__A1 core_0.fetch.prev_request_pc\[0\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4764__B2 net161 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_54_151 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_144_348 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_172_657 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6502__C _2123_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_43_836 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_42_313 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_200_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_43_858 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6471_ _2559_ _2642_ _2850_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_82_493 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_113_702 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_125_562 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_335 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6505__A2 _2604_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7702__A1 _1085_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_8210_ _0386_ clknet_leaf_31_i_clk net82 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_2
X_5422_ _1375_ _1861_ _1862_ _1838_ _1863_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_112_212 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput202 net202 sr_bus_data_o[2] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_70_699 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_11_733 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8141_ _0317_ clknet_leaf_90_i_clk core_0.execute.rf.reg_outputs\[1\]\[0\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_2_465 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5353_ _1800_ _1801_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__6269__A1 _2346_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4304_ _0902_ _0921_ _0922_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
X_8072_ _0248_ clknet_leaf_103_i_clk core_0.execute.rf.reg_outputs\[6\]\[11\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_227_625 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5284_ core_0.dec_jump_cond_code\[4\] _1193_ _1733_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_226_102 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4819__A2 core_0.fetch.submitable vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7023_ _1372_ _1939_ _3238_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4235_ _0824_ net57 _0853_ _0854_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_4
XTAP_TAPCELL_ROW_52_1140 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_226_157 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5492__A2 _1924_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4166_ core_0.dec_mem_long core_0.execute.sreg_long_ptr_en _0785_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_0_65_72 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6744__I _1963_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_97_508 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_179_212 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4097_ _0714_ _0715_ _0716_ _0717_ _0718_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_0_78_711 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7925_ _0003_ clknet_leaf_9_i_clk core_0.decode.oc_alu_mode\[13\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_139_109 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6992__A2 _3209_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_148_621 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7856_ core_0.fetch.current_req_branch_pred clknet_leaf_71_i_clk core_0.fetch.prev_req_branch_pred
+ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_148_643 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_147_120 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_175_440 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_37_129 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_438 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6807_ _2990_ _3065_ _3080_ _0297_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_147_142 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_3_6_0_i_clk clknet_0_i_clk clknet_3_6_0_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XTAP_TAPCELL_ROW_191_2806 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_7787_ core_0.dec_rf_ie\[7\] _1133_ _3827_ _3850_ _3855_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_4999_ _0769_ _1442_ _1443_ core_0.execute.rf.reg_outputs\[3\]\[0\] _1447_ _1448_
+ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_0_162_101 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_34_803 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6738_ _2996_ _3022_ _3040_ _0268_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_151_808 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_33_313 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_387 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_482 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6669_ core_0.execute.rf.reg_outputs\[6\]\[1\] _3000_ _2984_ _3002_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_61_644 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_116_562 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_116_584 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_103_212 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5028__C _1476_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_230_3272 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_131_554 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output170_I net170 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5180__A1 _0776_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_189_2779 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_245_422 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_217_124 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_217_146 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6680__A1 _2967_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5483__A2 net214 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_232_127 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_214_831 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5235__A2 _1683_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_66_1309 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_69_722 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_213_363 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_17_717 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6983__A2 _3184_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_766 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_29_619 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4994__A1 _0770_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_185_248 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_107 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_56_427 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_232_65 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6735__A2 _3020_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_139_698 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4746__A1 net57 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_37_663 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_279 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5943__B1 _2265_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_153_123 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_37_685 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_836 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_24_302 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_4_708 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_858 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_107_562 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6499__A1 _1109_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_134_370 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_34 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_12_508 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6499__B2 _1987_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_150_830 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_77_1438 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_40_839 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7160__A2 _3358_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_177_18 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_110_749 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_209_614 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_208_113 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_166_2510 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4349__I _0965_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4020_ _0641_ _0646_ _0647_ _0648_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_0_205_842 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6018__A4 _1549_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_189_554 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4029__A3 _0526_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_88_1567 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_5971_ _1458_ _2007_ _2144_ _1457_ _2362_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_0_150_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_149_418 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_126_99 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7710_ _2242_ _1134_ _3758_ _3806_ _1283_ _0474_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi221_2
X_4922_ _1385_ _1386_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_59_265 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_47_416 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_192_708 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_736 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7641_ _3732_ _3750_ _3751_ _0460_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_129_142 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_191_207 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_758 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_157_462 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4853_ _0860_ _1306_ _1339_ _0084_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__6726__A2 _3021_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_191_229 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5908__I _1641_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_28_652 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8040__CLK clknet_leaf_81_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4588__I1 core_0.ew_data\[8\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_62_419 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7572_ core_0.execute.pc_high_out\[2\] _3672_ _3694_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_4784_ _1290_ _1296_ _0058_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_28_685 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_780 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_145_679 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6523_ _2893_ _2900_ _2244_ _2901_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_43_644 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_132_307 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_82_290 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_42_132 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_15_346 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_132_329 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6454_ _2826_ _2832_ _2834_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_99_1696 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_42_165 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_30_305 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_485 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5162__A1 _0776_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5405_ _1747_ _1843_ _1848_ _0127_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_6385_ _2122_ _2103_ _2113_ _2766_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_2_273 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_101_749 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8124_ _0300_ clknet_leaf_96_i_clk core_0.execute.rf.reg_outputs\[3\]\[15\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_140_395 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_100_237 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5336_ _1783_ _1784_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_208_3005 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_55_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_239_282 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_227_422 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_167_51 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_110_1830 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_8055_ _0231_ clknet_leaf_104_i_clk core_0.execute.rf.reg_outputs\[7\]\[10\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5267_ _1714_ _1715_ _1705_ _1716_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_227_466 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_242_403 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7006_ core_0.execute.alu_mul_div.mul_res\[5\] _3222_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_4218_ net56 core_0.fetch.out_buffer_data_instr\[26\] _0824_ _0837_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_4
X_5198_ _0770_ _0767_ core_0.execute.rf.reg_outputs\[7\]\[1\] _1647_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_2
XTAP_TAPCELL_ROW_126_2026 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input27_I i_mem_data[15] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_242_436 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_214_127 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_242_447 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4149_ _0767_ _0768_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_98_839 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_223_661 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6414__A1 _2346_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5217__A2 _0773_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_223_683 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_211_834 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6965__A2 _3184_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7908_ _0099_ clknet_leaf_83_i_clk core_0.fetch.flush_event_invalidate vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__4976__A1 core_0.execute.sreg_priv_control.o_d\[14\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_195_557 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4976__B2 _1390_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_427 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_219_3145 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_66_747 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7519__B _3651_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7839_ _0032_ clknet_leaf_67_i_clk core_0.fetch.out_buffer_data_instr\[16\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_176_771 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6717__A2 _3021_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_121_1970 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_61_1239 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4728__A1 net47 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_65_268 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_232_3301 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_53_419 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_65_279 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_136_657 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_696 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7390__A2 net79 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_202_57 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5039__B _0779_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_137_2155 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_22_775 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_199_Left_446 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_61_430 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_151_627 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_150_2311 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3951__A2 _0528_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output95_I net95 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_839 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_61_485 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_132_863 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_150_159 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7254__B _3409_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6102__B1 _2249_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_72_1379 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_243_3430 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_148_2284 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_245_296 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_214_650 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_88_305 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_161_2440 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_199_863 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5208__A2 _0767_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_88_349 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_243_20 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_186_524 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8063__CLK clknet_leaf_109_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_158_237 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4967__B2 _1391_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_174_708 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_139_440 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_438 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_84_522 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_174_719 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7429__B _3553_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_173_207 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_201_399 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6708__A2 _3021_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_139_484 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_173_229 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_194_590 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_577 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4719__A1 net43 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_37_460 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_166_292 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_154_454 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_4_516 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5392__A1 _1233_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_126_167 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_655 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_21_66 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_154_498 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_25_666 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_88 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_172_2580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_80_794 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_97_37 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5144__A1 _1481_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7164__B _3357_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_110_513 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_122_384 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6170_ core_0.decode.oc_alu_mode\[7\] _2156_ _2022_ core_0.decode.oc_alu_mode\[6\]
+ _2556_ _2557_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_0_209_422 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_20_371 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_198_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_237_742 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_209_433 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5121_ core_0.execute.rf.reg_outputs\[6\]\[10\] _1435_ net218 core_0.execute.rf.reg_outputs\[1\]\[10\]
+ _1570_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_237_764 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5447__A2 _1812_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7611__C _3673_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5052_ _1500_ _1501_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XPHY_EDGE_ROW_127_Right_127 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
X_4003_ _0517_ core_0.execute.rf.reg_outputs\[3\]\[8\] _0549_ _0632_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_0_211_119 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_EDGE_ROW_212_Left_459 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__6947__A2 _1711_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_220_664 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5954_ _2278_ _2345_ _0179_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_48_725 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_220_675 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_165_708 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4905_ _1363_ _1368_ _1370_ _0105_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_175_2609 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_47_1072 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_192_527 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_75_555 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5885_ _2277_ _0178_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_7_310 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7624_ core_0.execute.pc_high_buff_out\[1\] _3732_ _1216_ _3739_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_35_419 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_8_855 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_90_514 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_123 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4836_ core_0.decode.i_instr_l\[13\] _1307_ _1328_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_118_657 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_99_i_clk_I clknet_4_7__leaf_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_16_633 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5383__A1 _1748_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7555_ net194 _3675_ _3678_ _3679_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_4767_ _1284_ _1287_ _0050_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_145_487 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_761 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_214_3075 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_31_603 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_15_154 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6506_ _2881_ _2882_ _2883_ _2626_ _2884_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai211_4
XFILLER_0_71_772 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_214_3086 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_7486_ net106 _3633_ _3634_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_160_457 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4698_ core_0.fetch.out_buffer_data_instr\[6\] net66 _1246_ _1247_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_30_102 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_221_Left_468 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
X_6437_ _1061_ _1702_ _2072_ _1109_ _2741_ _2817_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_0_3_582 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5686__A2 _1549_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_132_2096 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_30_179 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6368_ core_0.execute.alu_mul_div.div_res\[11\] _2332_ _2279_ _2750_ vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_2
XTAP_TAPCELL_ROW_186_2749 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_87_92 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8107_ _0283_ clknet_leaf_96_i_clk core_0.execute.rf.reg_outputs\[4\]\[14\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5319_ core_0.execute.alu_mul_div.div_cur\[2\] _1600_ _1767_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__xor2_2
X_6299_ _2673_ _2675_ _2682_ _2683_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA__6635__A1 core_0.execute.rf.reg_outputs\[7\]\[7\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5438__A2 _1812_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_8038_ _0215_ clknet_leaf_78_i_clk core_0.ew_reg_ie\[5\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__dffq_2
XANTENNA_output133_I net133 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8336__D _0512_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_230_Left_477 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_97_113 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_230_439 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4249__I0 net64 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_201_2919 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6938__A2 _1831_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_195_310 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_27_834 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7060__A1 _2648_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4949__A1 _1381_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_725 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5610__A2 _1637_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_210_174 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_197_2878 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_78_393 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_155_207 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_195_387 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_39_769 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_93_352 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4452__I core_0.decode.i_instr_l\[4\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_26_419 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_123 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_19_471 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_780 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_668 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_136_454 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_124_605 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4177__A2 _0795_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_191_582 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_123_104 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_151_413 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_124_649 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_22_603 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_229_Right_229 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_22_614 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_151_457 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_34_496 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_61_282 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_21_146 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6874__A1 _2981_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_120_855 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7712__B _3807_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_238_53 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6626__A1 net33 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_218_263 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_238_86 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_218_285 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_7_592 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5232__B _1480_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_233_244 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_233_277 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_89_647 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4652__A3 _1200_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_88_124 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6929__A2 _1221_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_85_1537 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7051__A1 _1224_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_202_664 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_186_332 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_186_343 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_186_354 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_522 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5601__A2 _1599_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_201_174 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_29_224 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_85_842 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_201_185 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_107 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_186_387 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_129 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_139_270 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4362__I net75 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_32_65 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_29_279 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5670_ _2069_ _2070_ _2071_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_2
XANTENNA__5365__A1 core_0.execute.alu_mul_div.div_cur\[1\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
X_4621_ core_0.execute.alu_flag_reg.o_d\[2\] core_0.execute.alu_flag_reg.o_d\[0\]
+ _1180_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_127_476 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_154_251 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_290 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_836 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_113_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_4_313 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_858 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7340_ net201 _3502_ _3511_ _3512_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_13_614 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3915__A2 _0542_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4552_ _1037_ _1095_ _1132_ _1135_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_142_457 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_130_619 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_96_1666 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_7271_ net87 _3449_ _3450_ _1735_ _3451_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_40_444 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_123_682 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4483_ _1068_ _1075_ _1076_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_40_466 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_12_157 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6222_ _2588_ _2607_ _1114_ _2608_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_0_110_365 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6153_ _1378_ _2538_ _2539_ _2540_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_237_550 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_110_387 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6617__A1 core_0.execute.rf.reg_outputs\[7\]\[4\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
X_5104_ _1551_ _1552_ _1553_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_0_209_274 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6084_ _1061_ _1683_ _2462_ _1109_ _2473_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__7290__A1 net75 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5142__B _1590_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5035_ _0770_ _0767_ _0775_ _1484_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_4
XTAP_TAPCELL_ROW_181_2679 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_224_277 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_240_737 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_196_107 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_49_1101 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5840__A2 _2209_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_18_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_73_72 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_94 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6986_ _1366_ _3202_ _3204_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_177_343 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_24_804 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_48_522 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5937_ _2281_ core_0.execute.alu_mul_div.mul_res\[1\] _0799_ _2329_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_105_1773 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_177_376 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_193_836 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_48_555 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_341 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4272__I core_0.fetch.prev_request_pc\[9\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_216_3104 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_193_858 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_192_335 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_75_352 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_63_525 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_300 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5868_ core_0.execute.sreg_priv_control.o_d\[0\] _1385_ _2260_ net1 _2261_ vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_2
X_7607_ core_0.execute.pc_high_out\[7\] _3723_ _3724_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_63_547 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4159__A2 core_0.dec_l_reg_sel\[0\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5356__A1 core_0.execute.alu_mul_div.div_cur\[12\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_133_402 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4819_ _1315_ core_0.fetch.submitable _1316_ _0073_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_28_290 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_162 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_105_104 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_32_892 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_5799_ _2197_ _2198_ _2199_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_16_463 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_134_2125 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_7538_ _3663_ _3665_ _0443_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_44_794 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_133_468 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_282 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_31_422 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5108__A1 net95 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_114_660 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_114_671 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_120_107 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5108__B2 _0708_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_160_287 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7469_ core_0.execute.mem_stage_pc\[15\] _3621_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_31_466 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6856__A1 _2940_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_102_855 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_101_343 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput79 net79 dbg_pc[1] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XTAP_TAPCELL_ROW_227_3233 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_228_550 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6608__A1 _2929_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_215_200 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7805__B1 _3866_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4882__A3 _0727_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_228_594 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_216_745 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_208_34 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_215_244 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6084__A2 _1683_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_145_2254 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_4_562 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4095__A1 _0565_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_231_737 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_169_811 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_230_247 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7033__A1 _1226_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_308 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_85_105 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_19_Right_19 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_67_842 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4398__A2 _0947_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_195_162 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_78_190 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_156_527 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_168_387 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_183_313 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_555 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_566 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_238_3373 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_80_1467 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_171_508 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_54_547 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_80_1478 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8101__CLK clknet_leaf_107_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_152_722 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_156_2383 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4910__I _1374_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_35_772 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5898__A2 _1603_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_124_446 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_260 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_720 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_580 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6330__C _2332_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_152_777 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_22_422 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_2_839 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_111_118 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_28_Right_28 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_105_693 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6847__A1 _2992_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_120_663 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7442__B _3545_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6837__I _0722_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4173__I2 core_0.ew_reg_ie\[6\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_47_i_clk_I clknet_4_12__leaf_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_206_200 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_207_745 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7272__A1 _3384_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_206_255 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_89_422 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_222_737 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5897__B _1652_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_178_107 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_37_Right_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_221_247 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__7024__A1 _2567_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6840_ core_0.execute.rf.reg_outputs\[2\]\[10\] _3092_ _3098_ _3100_ vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__4389__A2 _0966_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_9_416 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6771_ core_0.execute.rf.reg_outputs\[4\]\[13\] _3049_ _3057_ _3060_ vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_230_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_3983_ net89 _0578_ _0614_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_9_438 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_147_538 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_159_398 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_175_858 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_18_728 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5722_ _2102_ _2123_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XTAP_TAPCELL_ROW_44_1042 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_84_160 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_683 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_91_119 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7327__A2 _2521_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_162_508 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5653_ _1789_ _2053_ _2054_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_115_402 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4820__I core_0.decode.i_instr_l\[8\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4604_ core_0.ew_addr\[0\] _1167_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__7336__C _1950_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_46_Right_46 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_26_794 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_4_132 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5584_ core_0.dec_mem_we net159 _1985_ _1986_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_41_720 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_411 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_25_282 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_115_479 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_211_3045 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_102_107 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7323_ core_0.dec_alu_flags_ie _3495_ _1955_ _3496_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4535_ core_0.decode.oc_alu_mode\[11\] _1121_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XANTENNA__4561__A2 _1062_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_229_303 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_7254_ net85 _3435_ _3409_ _3436_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_4466_ _1059_ _1053_ _1060_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_229_347 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_110_140 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6205_ _2031_ _2553_ _2021_ _2591_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XANTENNA__4313__A2 _0851_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5510__A1 _1811_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7185_ _1748_ _3377_ _0378_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_111_696 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_183_2708 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_4397_ _0959_ _1005_ _1006_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_244_317 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_55_1171 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6136_ core_0.execute.alu_mul_div.div_res\[5\] _2332_ _2523_ _2524_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_225_542 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7263__A1 _1400_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7263__B2 _1430_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6067_ _2454_ _2456_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XPHY_EDGE_ROW_55_Right_55 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_213_726 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_212_203 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_107_1802 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_1_521 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_5018_ _1466_ _1467_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XTAP_TAPCELL_ROW_222_3174 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_212_247 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_68_617 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_37_951 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_240_589 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_191_50 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7566__A2 core_0.execute.pc_high_out\[1\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_37_962 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_166_803 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_842 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_67_138 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_177_173 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_220_291 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6969_ _3180_ _3181_ _3182_ _3187_ _3188_ _0351_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai221_1
XTAP_TAPCELL_ROW_140_2195 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_194_2837 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_76_661 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_48_374 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_76_683 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_165_346 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_193_699 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_118_251 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7527__B _3651_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5329__A1 core_0.execute.alu_mul_div.div_cur\[5\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_64_Right_64 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_51_506 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_17_772 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_51_517 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_173_390 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_106_457 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_118_1931 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_63_399 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_121_416 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4552__A2 _1095_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_31_252 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_9_621 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_236_807 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_7_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_219_66 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_73_Right_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__6057__A2 _2250_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7254__A1 net85 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_720 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_0_i_clk i_clk clknet_0_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_203_203 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_216_597 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5804__A2 _2183_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_235_54 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_188_438 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_235_65 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_235_76 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_169_663 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6325__C _2294_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_80_18 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5568__A1 _1419_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_158_2412 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_168_195 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4240__A1 core_0.fetch.out_buffer_valid vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7309__A2 _3398_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_82_Right_82 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_104_69 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_183_154 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_15_689 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_109_262 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_172_839 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_183_187 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6517__B1 _2577_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_125_755 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_152_541 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_81_174 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4543__A2 _1092_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_2_647 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_93_1625 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_4320_ net68 core_0.fetch.out_buffer_data_instr\[8\] _0725_ _0938_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__7172__B core_0.execute.alu_mul_div.div_res\[6\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7493__A1 _3637_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_169_2541 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_4251_ net63 core_0.fetch.out_buffer_data_instr\[3\] _0724_ _0870_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_227_829 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_91_Right_91 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_120_493 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_238_177 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_226_317 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_129_66 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4182_ _0799_ _0800_ _0801_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_4
XANTENNA_input1_I i_core_int_sreg[0] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_180_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6048__A2 _1114_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_54_30 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7941_ _0119_ clknet_leaf_42_i_clk core_0.execute.sreg_priv_control.o_d\[13\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_7872_ _0064_ clknet_leaf_63_i_clk core_0.fetch.prev_request_pc\[15\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_222_589 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_49_116 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_54_85 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_203_792 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_34_921 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6823_ _2951_ _3086_ _3090_ _0303_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_58_650 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_224 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_92_417 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_102_1732 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_147_335 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6220__A2 _2590_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_45_300 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6754_ core_0.execute.rf.reg_outputs\[4\]\[5\] _3049_ _3045_ _3051_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__4231__A1 core_0.fetch.out_buffer_valid vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3966_ _0565_ _0524_ _0527_ core_0.execute.rf.reg_outputs\[6\]\[11\] _0598_ vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_0_147_368 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_116_700 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5705_ _2104_ _2105_ _1819_ _2106_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_9_279 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_190_636 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6685_ core_0.execute.rf.reg_outputs\[6\]\[8\] _3006_ _3004_ _3011_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3897_ _0532_ _0533_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_45_366 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4550__I _1132_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_162_349 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_60_314 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5636_ _1503_ _1504_ _2037_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_EDGE_ROW_162_Left_409 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_60_325 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_85_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_14_731 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_170_360 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_143_585 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5567_ _1419_ _0739_ _0158_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_57_1200 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_41_550 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_496 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_103_438 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7306_ _2864_ _3479_ _3480_ _3481_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_131_769 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_13_274 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4518_ _1107_ _1053_ _1108_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_8286_ _0462_ clknet_leaf_32_i_clk core_0.execute.pc_high_buff_out\[7\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5498_ _1930_ _1483_ _1658_ _1663_ _1931_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XANTENNA_input57_I i_req_data[27] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7237_ _1414_ core_0.execute.sreg_irq_pc.o_d\[5\] _1406_ _1431_ _1736_ _3421_ vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XANTENNA__7484__A1 _3514_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_245_604 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4449_ _1038_ _1043_ _1044_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_4
XANTENNA__4298__A1 core_0.fetch.prev_request_pc\[3\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1_691 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_3_2_0_i_clk clknet_0_i_clk clknet_3_2_0_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XTAP_TAPCELL_ROW_113_1872 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_224_3203 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_7168_ _1369_ _1915_ _1230_ _3367_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_0_244_147 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_95_81 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7236__A1 _2526_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_95_92 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_129_2057 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6119_ _1999_ _2009_ _2507_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XPHY_EDGE_ROW_171_Left_418 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
X_7099_ _1230_ _1920_ _3308_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_213_512 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7787__A2 _1133_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_142_2213 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5798__A1 _1987_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_213_556 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_206_2980 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_201_718 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_95_200 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_197_257 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_96_734 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_96_745 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7539__A2 _1398_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_197_279 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_185_419 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_95_222 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_95_244 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_138_302 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_469 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_139_836 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_139_858 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_193_430 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6211__A2 _2594_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5014__A3 _0549_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5984__C _1603_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_235_3332 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4222__A1 _0726_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_311 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_180_Left_427 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__4773__A2 _1285_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5970__A1 _1137_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_63_130 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_153_327 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_733 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_63_152 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_153_349 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_12_659 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_63_163 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_36_399 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_106_243 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_196 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7711__A2 _1064_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_134_563 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_153_2353 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_122_714 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_122_725 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_161_371 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4525__A2 core_0.decode.i_instr_l\[2\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_712 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_122_769 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_734 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_208_317 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_246_3461 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_246_3472 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_246_3483 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_246_20 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_235_136 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_164_2482 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_231_331 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_188_224 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6450__A2 _2531_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4461__A1 core_0.decode.i_instr_l\[0\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_231_386 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_176_419 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_197_780 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87_767 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_86_266 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6202__A2 _2587_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5005__A3 core_0.decode.oc_alu_mode\[7\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_156_121 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_157_644 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_119 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_74_428 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4213__A1 _0724_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_322 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_41_1001 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_55_653 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4764__A2 _1285_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5961__A1 net80 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5961__B2 _2245_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_54_163 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_125_541 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_171_146 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_54_174 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6470_ _2845_ _2848_ _2849_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_131_78 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_42_347 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_113_714 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7702__A2 _1098_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5421_ _1374_ _1856_ _1862_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_140_511 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_70_667 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_30_509 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput203 net203 sr_bus_data_o[3] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_113_758 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_140_544 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8140_ _0316_ clknet_leaf_98_i_clk core_0.execute.rf.reg_outputs\[2\]\[15\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5352_ core_0.execute.alu_mul_div.div_cur\[12\] _1701_ _1800_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_100_419 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4303_ _0905_ _0920_ _0921_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__7010__S0 _1226_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_140_599 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7466__A1 _0563_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_767 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8071_ _0247_ clknet_leaf_100_i_clk core_0.execute.rf.reg_outputs\[6\]\[10\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_10_255 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5283_ core_0.execute.sreg_irq_pc.o_d\[0\] _1732_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_239_486 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7022_ _3224_ _3230_ _3236_ _3237_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_4234_ core_0.fetch.out_buffer_valid _0852_ _0853_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_52_1141 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7218__A1 _3384_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_226_169 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4165_ _0783_ _0782_ _0784_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_4
XANTENNA__7769__A2 _3766_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6977__B1 _3181_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4096_ _0568_ _0535_ _0536_ core_0.execute.rf.reg_outputs\[2\]\[0\] _0717_ vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_0_223_865 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7924_ _0002_ clknet_leaf_121_i_clk core_0.decode.oc_alu_mode\[12\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_4
XFILLER_0_195_728 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_179_279 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7855_ _0048_ clknet_leaf_69_i_clk core_0.fetch.out_buffer_valid vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_81_72 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_187_290 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_37_119 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6806_ core_0.execute.rf.reg_outputs\[3\]\[12\] _3070_ _3072_ _3080_ vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__4204__A1 _0723_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4998_ _0710_ _1444_ _1446_ _1447_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_7786_ _1136_ _3854_ _0502_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_191_2807 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_163_614 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_18_333 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_63_1270 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_92_247 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_136_839 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4755__A2 _1238_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_46_664 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3949_ _0534_ _0542_ _0544_ core_0.execute.rf.reg_outputs\[5\]\[12\] _0582_ vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_4
X_6737_ core_0.execute.rf.reg_outputs\[5\]\[15\] _3020_ _3031_ _3040_ vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__5952__A1 _2244_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_63_i_clk clknet_4_15__leaf_i_clk clknet_leaf_63_i_clk vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_6668_ _2940_ _2999_ _3001_ _0237_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__5165__C1 _1606_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5619_ _1761_ _2019_ _2020_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__5704__A1 _1123_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_5_282 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6599_ _2936_ _2946_ _2947_ _0222_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_103_224 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_143_393 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_230_3273 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_60_166 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_60_177 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8338_ _0514_ clknet_leaf_16_i_clk core_0.decode.o_submit vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__dffq_4
Xclkbuf_leaf_78_i_clk clknet_4_13__leaf_i_clk clknet_leaf_78_i_clk vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_103_268 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output163_I net163 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8312__CLK clknet_leaf_76_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_8269_ _0445_ clknet_leaf_23_i_clk core_0.execute.sreg_irq_flags.o_d\[3\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_218_615 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7209__A1 _2390_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_245_467 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_217_158 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6680__A2 _2999_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_233_629 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_226_681 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_213_320 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_241_640 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_216_34 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6156__B _2541_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_213_342 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_16_i_clk clknet_4_8__leaf_i_clk clknet_leaf_16_i_clk vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_TAPCELL_ROW_17_718 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_240_183 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_96_542 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_244 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_68_255 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_wire212_I net213 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_56_406 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_715 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_56_439 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_37_620 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_480 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_759 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_153_102 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4746__A2 _1241_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_193_282 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_269 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_126_327 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5943__A1 core_0.execute.sreg_irq_pc.o_d\[1\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_181_422 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4404__B _0970_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5943__B2 core_0.execute.alu_flag_reg.o_d\[1\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_52_601 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_461 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_37_697 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_314 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_36_185 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_51_111 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_153_168 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_40_807 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_52_667 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_77_1439 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6111__S _2102_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_108_Right_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_110_717 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7448__A1 _0604_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_103_780 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_209_626 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7006__I core_0.execute.alu_mul_div.mul_res\[5\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_166_2500 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_20_597 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6120__A1 _2014_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_66 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6671__A2 _3000_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_223_106 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_189_511 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_126_34 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_88_1568 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7620__A1 core_0.execute.pc_high_buff_out\[0\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4029__A4 core_0.execute.rf.reg_outputs\[2\]\[6\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_200 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5970_ _1137_ _1676_ _1061_ _2361_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_126_78 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_126_89 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4921_ _1384_ _1385_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_59_255 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4985__A2 _0773_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_143_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_59_277 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7640_ core_0.execute.pc_high_buff_out\[5\] _3731_ _1216_ _3751_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__6187__A1 _2346_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4852_ core_0.decode.i_imm_pass\[2\] _1307_ _1339_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_177_2640 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_185_772 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5234__I0 net188 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_28_642 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_247 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_118_839 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_200_592 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_144_102 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_157_496 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7571_ net221 _3675_ _3692_ _3693_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_4783_ core_0.fetch.prev_request_pc\[9\] net225 _0880_ net176 _1296_ vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai22_1
XANTENNA__5934__A1 _1831_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_28_664 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_145_647 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_349 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_55_472 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6522_ _2866_ _2899_ _2900_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_43_623 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_100 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_174 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5129__C _1531_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_144_157 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_111 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_420 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_132_319 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7687__A1 _1038_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6453_ _2826_ _2832_ _2833_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_42_144 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_99_1697 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_141_842 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_30_317 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5404_ core_0.execute.alu_mul_div.div_cur\[4\] _1838_ _1816_ _1847_ _1848_ vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_3_764 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_113_566 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6384_ _1501_ _1455_ _2765_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or2_1
X_8123_ _0299_ clknet_leaf_97_i_clk core_0.execute.rf.reg_outputs\[3\]\[14\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5335_ core_0.execute.alu_mul_div.div_cur\[8\] _1756_ _1783_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_208_3006 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_8054_ _0230_ clknet_leaf_103_i_clk core_0.execute.rf.reg_outputs\[7\]\[9\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_227_434 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5266_ _1519_ _1715_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XTAP_TAPCELL_ROW_110_1831 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_48_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_7005_ _3212_ _3177_ _3221_ _0354_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_4217_ net51 core_0.fetch.out_buffer_data_instr\[21\] _0723_ _0836_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA_clkbuf_leaf_95_i_clk_I clknet_4_7__leaf_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6662__A2 _2935_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_215_629 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5197_ core_0.execute.rf.reg_outputs\[5\]\[1\] _1646_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_126_2027 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_98_807 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_4148_ core_0.dec_l_reg_sel\[1\] _0767_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_207_191 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7611__A1 _3675_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6414__A2 net197 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_168_706 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4079_ _0533_ _0541_ _0543_ core_0.execute.rf.reg_outputs\[5\]\[1\] _0701_ vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_0_183_84 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_223_695 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_203_2950 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_7907_ _0098_ clknet_leaf_51_i_clk core_0.fetch.dbg_out vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_78_564 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4976__A2 _1393_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_66_737 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_219_3135 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6178__A1 _2295_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_219_3146 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_38_439 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_19_620 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_225 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7838_ _0031_ clknet_leaf_73_i_clk core_0.fetch.out_buffer_data_instr\[15\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_121_1960 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4728__A2 _1253_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5925__A1 _1596_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_163_422 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_175_282 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_232_3302 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_18_141 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7769_ core_0.dec_rf_ie\[0\] _3766_ _3833_ _3843_ _3844_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_202_47 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_151_606 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_34_634 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_22_776 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_137_2156 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_190_263 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_135_168 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_190_274 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_667 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_22_807 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_150_2312 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_21_306 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_33_166 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6350__A1 _2090_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_104_577 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output88_I net88 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5055__B _1460_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_246_710 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_245_220 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6102__B2 core_0.execute.pc_high_buff_out\[5\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_243_3431 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7852__CLK clknet_leaf_67_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6665__I _2998_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6653__A2 _2962_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_233_415 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4664__A1 core_0.decode.i_flush vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_148_2285 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_227_66 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_205_139 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_199_842 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_199_853 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_88_317 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_161_2441 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_214_662 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7602__A1 net215 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5208__A3 core_0.execute.rf.reg_outputs\[3\]\[3\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8208__CLK clknet_leaf_32_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_202_824 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_243_10 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_241_492 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_159_739 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_243_43 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4967__A2 _1393_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_201_356 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_186_558 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_56_214 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6169__A1 _1761_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_167_761 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_56_247 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_166_260 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5916__A1 _1819_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_127_636 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4719__A2 _1253_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_71_206 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_181_241 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_645 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_64_291 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_133 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7669__A1 _0514_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_123_842 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_172_2581 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_80_784 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_97_16 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_40_637 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_150_661 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5144__A2 _1592_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_117_i_clk_I clknet_4_4__leaf_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5120_ core_0.execute.rf.reg_outputs\[5\]\[10\] _1486_ _1569_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_236_231 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6644__A2 _2962_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5051_ net91 _1492_ _1495_ _1499_ _1500_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai22_4
XFILLER_0_209_489 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4655__A1 net106 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4002_ _0565_ _0524_ _0527_ core_0.execute.rf.reg_outputs\[6\]\[8\] _0631_ vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_0_224_448 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_137_66 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_189_352 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_204_183 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_149_227 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_66 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_149_238 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_153_54 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5953_ _2242_ net201 _2190_ _2344_ _2345_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_177_547 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_737 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_153_76 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4904_ _1369_ _1221_ _1370_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_8_801 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_62_85 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5884_ core_0.ew_data\[0\] _2276_ _2190_ _2277_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_47_1073 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_164_219 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_118_625 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7623_ net201 _3733_ _3737_ _3738_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_35_409 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_145_422 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4835_ _1325_ _1327_ _0078_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_157_282 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_16_601 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_62_217 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_344 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_145_455 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4766_ core_0.fetch.prev_request_pc\[1\] _1285_ _0881_ net168 _1287_ vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_7554_ core_0.execute.pc_high_out\[0\] _3676_ _3677_ _3678_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_173_786 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6505_ _2133_ _2604_ _2883_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_214_3076 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_7485_ _1392_ _1206_ _3633_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_4697_ _1236_ _1246_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_15_177 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_113_330 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_rebuffer12_I net232 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6436_ _1137_ _1702_ _2740_ _2816_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__6332__A1 _2714_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_113_352 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_113_385 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_140_171 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7875__CLK clknet_leaf_83_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6367_ _2281_ _2747_ _2748_ _1114_ _2749_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XTAP_TAPCELL_ROW_132_2097 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_186_2739 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4894__A1 _1321_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_228_743 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8106_ _0282_ clknet_leaf_94_i_clk core_0.execute.rf.reg_outputs\[4\]\[13\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5318_ core_0.execute.alu_mul_div.div_cur\[3\] _1765_ _1766_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_6298_ _1107_ _2677_ _2681_ _2682_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_227_253 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6635__A2 _2962_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5249_ _1695_ _1697_ _1698_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_2
X_8037_ _0214_ clknet_leaf_80_i_clk core_0.ew_reg_ie\[4\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_242_212 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4646__A1 core_0.dec_jump_cond_code\[4\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_230_407 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_3_Left_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__6399__A1 _1088_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_97_125 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_196_812 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_223_492 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_211_632 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_27_835 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7060__A2 _3181_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4949__A2 net215 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_704 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_195_344 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_39_737 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_211_687 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_195_366 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_211_698 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_197_2879 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_38_247 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_556 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_94_865 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_136_400 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_195_399 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_450 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_164_731 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_53_206 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_148_293 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_109_658 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_163_252 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_191_572 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_136_477 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_431 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_193_Right_193 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_49_Left_296 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_105_842 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5564__I _1963_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_62_784 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_114 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_22_659 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6874__A2 _3107_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_131_193 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4885__A1 _1279_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_219_743 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_246_540 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_219_776 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_218_275 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_233_212 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_7_593 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_199_650 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_16_34 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_199_661 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_85_1527 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_107_69 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_16_67 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_85_1538 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_198_171 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7051__A2 _3215_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_16_78 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_186_322 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_201_131 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_201_142 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5062__A1 _1460_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_159_558 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_394 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_96_191 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_201_197 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_707 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_578 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_139_282 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA_clkbuf_leaf_43_i_clk_I clknet_4_9__leaf_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_32_55 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_84_364 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_217 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4620_ _1174_ _1177_ _1178_ _1179_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_0_72_559 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5365__A2 _1812_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4412__I1 _0857_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_25_453 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_4_325 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4551_ _1133_ _1134_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XPHY_EDGE_ROW_160_Right_160 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__3915__A3 _0544_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_106_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_13_626 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_190 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7270_ net87 _3449_ _3450_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_13_648 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_12_125 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_96_1667 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_4482_ _1042_ _1072_ _1074_ _1075_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_6221_ _2281_ _2606_ _2607_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_123_694 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6865__A2 _3114_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_122_193 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4876__A1 core_0.decode.i_imm_pass\[13\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6152_ _1378_ core_0.execute.sreg_irq_pc.o_d\[6\] _2539_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_110_377 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_237_562 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_225_702 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5103_ _0713_ _0718_ _1460_ _0719_ _1552_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai211_4
XANTENNA__6617__A2 _2962_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6083_ _1137_ _1683_ _1456_ _2472_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_209_286 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_224_223 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5034_ core_0.dec_l_reg_sel\[2\] core_0.dec_l_reg_sel\[1\] core_0.dec_l_reg_sel\[0\]
+ _1483_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_4
XANTENNA__7290__A2 net74 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_224_256 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_224_267 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_49_1102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_196_119 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_79_136 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_178_823 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_205_492 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_79_158 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_95_607 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_189_182 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_95_629 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6985_ _1372_ _1367_ core_0.execute.alu_mul_div.mul_res\[3\] _3202_ _3203_ vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_1
XANTENNA__5053__A1 _1482_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6254__B _2638_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_24_805 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4553__I _1051_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5936_ _2292_ _2299_ _2327_ _2328_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_0_137_208 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_105_1774 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_192_314 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_76_865 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_118_400 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_216_3105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_118_422 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_146_731 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5867_ _1196_ _1383_ _2247_ _2260_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and3_2
XFILLER_0_91_846 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7606_ core_0.execute.pc_high_out\[6\] core_0.execute.pc_high_out\[5\] core_0.execute.pc_high_out\[4\]
+ _3695_ _3723_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_0_8_664 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4818_ _0935_ core_0.fetch.submitable _1316_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_35_239 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5356__A2 _1803_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6553__A1 _2209_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5798_ _1987_ _2187_ _2183_ _2198_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_32_893 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_16_442 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_134_2115 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_173_594 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_367 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_134_2126 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_145_296 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_160_222 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7537_ core_0.execute.sreg_irq_flags.o_d\[1\] _3664_ core_0.execute.prev_sys _3665_
+ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_4749_ _0821_ _1238_ _1275_ _0044_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_90_389 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_160_244 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_160_255 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_189_72 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5108__A2 _0521_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6305__A1 core_0.execute.alu_mul_div.div_cur\[9\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
X_7468_ _3581_ _3620_ _0418_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_98_92 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_160_299 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_101_311 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6419_ _2051_ _2058_ _2695_ _2173_ _2171_ _2799_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai32_1
XANTENNA__6856__A2 _3107_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7399_ net37 _3563_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XTAP_TAPCELL_ROW_227_3234 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4331__A3 core_0.fetch.prev_request_pc\[0\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7805__A1 core_0.decode.i_instr_l\[14\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7805__B2 core_0.decode.i_instr_l\[11\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_215_212 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_4_563 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_145_2255 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_208_79 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4095__A2 _0541_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5292__A1 _1739_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_98_423 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5987__C _1480_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_187_119 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7033__A2 _1613_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_98_478 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_224_34 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_196_664 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_85_139 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_224_78 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_183_303 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_238_3363 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_94_651 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_238_3374 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_184_859 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_109_422 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_93_150 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_26_217 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_80_1468 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_66_397 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_57_Left_304 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_54_559 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_124_403 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_35_740 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_488 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_164_583 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_152_734 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_156_2384 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_151_244 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_807 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_112_609 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_592 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_34_294 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_105_672 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7344__I0 _3514_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_151_277 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4307__B1 _0886_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6847__A2 _3087_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_10_629 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7442__C _3598_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4173__I3 core_0.ew_reg_ie\[7\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_207_702 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_207_713 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XPHY_EDGE_ROW_66_Left_313 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_246_370 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_234_532 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_234_554 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_27_66 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_27_77 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_221_204 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6853__I _3106_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_178_119 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_77_629 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_134_34 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5035__A1 _0770_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_134_45 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6232__B1 _2534_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_76_128 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6783__A1 _2946_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3982_ _0609_ _0610_ _0611_ _0612_ _0613_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_4
X_6770_ _2990_ _3043_ _3059_ _0281_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__5586__A2 _1522_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_174_303 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_186_174 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_58_865 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5721_ _2118_ _2121_ _2102_ _2122_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XPHY_EDGE_ROW_75_Left_322 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_44_1043 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_223_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_190_807 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6802__B _3072_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_190_829 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_73_846 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_5_601 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5652_ _1576_ _2053_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__inv_3
XFILLER_0_26_762 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_4603_ _1166_ net145 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5418__B _1816_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4546__B1 _1064_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5583_ _1984_ _1985_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_41_732 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_211_3046 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_4534_ _1084_ _1090_ _1094_ _1039_ _1119_ _1120_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi221_4
X_7322_ _1209_ _2265_ _3495_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_0_4_166 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_4_177 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_40_242 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_170_597 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6838__A2 _3092_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7253_ _1742_ _3426_ _3435_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4465_ core_0.decode.oc_alu_mode\[6\] _1059_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_13_489 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4849__A1 _0851_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6204_ _2018_ _2589_ _2590_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_0_159_86 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7184_ _1362_ _3373_ core_0.execute.alu_mul_div.div_res\[11\] _3377_ vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XPHY_EDGE_ROW_84_Left_331 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
X_4396_ _0904_ _0950_ _1005_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_110_174 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_183_2709 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_55_1172 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_110_185 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6135_ _1433_ _2521_ _2522_ _0799_ _2523_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai211_2
XANTENNA__6066__A3 _2454_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6066_ _2357_ _2405_ _2454_ _2455_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_0_30_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5017_ core_0.dec_r_bus_imm _1466_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_240_524 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_1_522 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_222_3175 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_206_790 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_240_557 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_37_952 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_67_106 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4283__I _0838_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7566__A3 core_0.execute.pc_high_out\[0\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_93_Left_340 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_191_84 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6968_ _1652_ _3178_ _3188_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6774__A1 _2994_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_166_837 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_138_539 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_140_2196 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_64_802 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_194_2838 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_5919_ _2300_ _2304_ _2310_ _2311_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_0_76_673 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_119_742 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_192_133 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_75_161 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_91_610 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_118_230 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6899_ net97 _3130_ _3124_ _3134_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_91_632 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_192_177 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6526__A1 _2576_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5329__A2 _1715_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_180_317 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_36_559 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_146_572 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_180_328 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_436 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_134_745 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_output193_I net193 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_91_687 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_63_389 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4001__A2 _0594_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_118_1932 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_210_69 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6829__A2 _3092_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_9_622 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_101_130 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_101_174 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_101_185 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_228_381 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_244_863 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_204_716 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4068__A2 _0541_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_243_362 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_204_727 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6673__I _1963_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_243_373 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_188_406 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_231_524 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_59_618 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_86_404 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_58_139 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5568__A2 _0736_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6765__A1 _2986_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_67_640 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_168_163 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_158_2413 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_183_100 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_104_37 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_156_336 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_364 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7718__B _3810_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_54_301 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_172_807 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_184_667 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_54_312 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_109_241 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_120 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_137_572 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6517__B2 core_0.execute.sreg_irq_pc.o_d\[15\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_54_356 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_81_142 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_125_734 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_152_531 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_164_391 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_570 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_125_767 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_120_47 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_152_575 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_22_231 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5740__A2 _1552_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_140_737 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_22_242 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7453__B _3553_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_253 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_50_562 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_93_1626 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_1_136 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1_158 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4250_ net60 core_0.fetch.out_buffer_data_instr\[2\] _0724_ _0869_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_120_461 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_169_2542 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6540__I1 _2571_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4368__I net74 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4181_ core_0.execute.alu_mul_div.i_mod _0800_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_3
XFILLER_0_129_89 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5256__A1 _1513_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4059__A2 _0594_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_173_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_234_362 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_207_576 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_234_373 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_89_220 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7940_ _0118_ clknet_leaf_43_i_clk core_0.execute.sreg_priv_control.o_d\[12\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_179_417 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_222_557 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_7871_ _0063_ clknet_leaf_63_i_clk core_0.fetch.prev_request_pc\[14\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_89_286 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_148_804 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6822_ core_0.execute.rf.reg_outputs\[2\]\[2\] _3087_ _3083_ _3090_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_77_448 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5559__A2 _1955_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6756__A1 core_0.execute.rf.reg_outputs\[4\]\[6\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_34_922 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_147_314 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_147_325 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_148_848 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_58_662 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_174_111 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7628__B _1216_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_102_1733 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_159_196 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6753_ _2961_ _3042_ _3050_ _0273_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_147_347 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3965_ _0593_ _0594_ _0595_ _0596_ _0597_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai211_4
XFILLER_0_9_258 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_73_632 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5704_ _1123_ _1931_ net211 _1720_ _2105_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai211_2
XANTENNA__6024__S _1596_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6508__A1 _1457_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_162_317 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_174_177 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3896_ core_0.dec_r_reg_sel\[2\] _0532_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_6684_ _2977_ _2999_ _3010_ _0244_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__6508__B2 _1458_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_190_648 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_174_199 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3990__A1 _0565_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_60_304 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_838 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5635_ _1754_ _2035_ _2036_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_2
XANTENNA__7181__A1 _1748_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_143_553 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_103_406 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_130_203 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5566_ _1977_ _1957_ _1979_ _0157_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_57_1201 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_78_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_79_72 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_7305_ _1431_ _1426_ _3480_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_41_562 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4517_ core_0.decode.oc_alu_mode\[4\] _1107_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_8285_ _0461_ clknet_leaf_29_i_clk core_0.execute.pc_high_buff_out\[6\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5497_ net97 _1930_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_13_286 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7236_ _2526_ _3391_ _3420_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_218_819 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4448_ core_0.decode.i_instr_l\[1\] _1043_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_4
XANTENNA__4298__A2 _0857_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_113_1873 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_4379_ net87 _0991_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XTAP_TAPCELL_ROW_224_3204 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_186_73 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7167_ _3357_ _3366_ _0371_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__7236__A2 _3391_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6118_ _2012_ _2506_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_129_2058 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_7098_ _3286_ _3288_ _3306_ _3307_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__6707__B _3016_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5247__A1 _1479_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_142_2214 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_225_384 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6049_ core_0.execute.alu_mul_div.div_cur\[3\] _2279_ _2439_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_198_737 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5798__A2 _2187_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_206_2981 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_68_1330 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_240_365 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_95_212 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_200_218 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_178_450 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_output206_I net206 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_200_229 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_459 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_95_234 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_205_58 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_640 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8241__CLK clknet_4_9__leaf_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_166_623 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_418 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_138_336 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_154_807 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_166_667 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4222__A2 net46 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_126_509 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_235_3333 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_48_172 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_119_550 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_181_626 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5970__A2 _1676_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_367 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_63_142 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_181_648 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_24_518 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3981__A1 _0568_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7172__A1 _3358_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_153_2343 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_106_255 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_17_592 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_134_575 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_153_2354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4525__A3 _1078_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_134_597 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_161_394 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7475__A2 _1398_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5486__A1 _1226_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_246_3462 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_246_3473 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_217_830 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7227__A2 _3407_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_217_852 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_246_54 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_216_351 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_232_811 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6617__B _1978_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4916__I _1379_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_216_384 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_204_524 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_164_2483 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_216_395 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_99_540 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_189_759 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_87_702 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_99_562 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_188_247 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_188_258 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_59_426 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4461__A2 _1039_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_34 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_87_757 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_115_58 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6738__A1 _2996_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_157_623 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_129_325 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7448__B _3545_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5005__A4 core_0.decode.oc_alu_mode\[4\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_184_453 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5410__A1 core_0.execute.alu_mul_div.div_cur\[5\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_632 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_492 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_41_1002 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_144_317 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5961__A2 _2268_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_125_520 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3972__A1 _0597_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_171_136 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7163__A1 _1369_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_125_553 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_495 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_113_704 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_125_564 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5420_ _1782_ _1783_ _1861_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_152_361 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_112_203 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6910__A1 _2977_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_140_523 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_562 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7183__B _3357_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput204 net204 sr_bus_data_o[4] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
X_5351_ _1798_ _1702_ _1799_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_112_247 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5482__I _1909_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50_381 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_42 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4302_ _0908_ _0919_ _0920_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_8070_ _0246_ clknet_leaf_106_i_clk core_0.execute.rf.reg_outputs\[6\]\[9\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_2
X_5282_ _1431_ _1729_ _1730_ _1195_ _1731_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__7466__A2 _3546_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5477__A1 _1908_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8114__CLK clknet_leaf_107_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4233_ core_0.fetch.out_buffer_data_instr\[27\] _0852_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_7021_ _3235_ _3236_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_52_1131 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_52_1142 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_65_30 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4164_ _0767_ _0769_ _0783_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_241_107 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5229__A1 _1625_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5431__B _1816_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6019__S _1559_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4095_ _0565_ _0541_ _0544_ core_0.execute.rf.reg_outputs\[5\]\[0\] _0716_ vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_0_234_181 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6977__A1 _3175_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_223_855 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6977__B2 _2386_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7923_ _0001_ clknet_leaf_120_i_clk core_0.decode.oc_alu_mode\[11\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_4
XFILLER_0_222_387 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_210_527 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_194_206 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_172_53 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7854_ _0047_ clknet_leaf_66_i_clk core_0.fetch.out_buffer_data_instr\[31\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_194_239 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_65_407 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_77_267 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6805_ _2988_ _3065_ _3079_ _0296_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_65_418 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_136_807 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_148_667 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7785_ core_0.dec_rf_ie\[6\] _1133_ _3827_ _3848_ _3854_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__4204__A2 net58 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_18_312 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4997_ _1445_ _1446_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XANTENNA__5401__A1 core_0.execute.alu_mul_div.div_cur\[5\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_105_80 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_191_2808 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_63_1271 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_92_259 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6736_ _2994_ _3022_ _3039_ _0267_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_163_626 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_345 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3948_ core_0.execute.rf.reg_outputs\[2\]\[12\] _0581_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA_clkbuf_leaf_91_i_clk_I clknet_4_6__leaf_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_45_142 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_18_356 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5952__A2 _2334_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_18_378 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_116_531 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_484 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6667_ core_0.execute.rf.reg_outputs\[6\]\[0\] _3000_ _2984_ _3001_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3879_ core_0.dec_r_reg_sel\[2\] _0515_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__inv_4
XFILLER_0_60_123 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_12_Left_259 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__5165__B1 _1605_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5618_ net100 _1611_ _1492_ _2019_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__5704__A2 _1931_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_104_737 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_116_597 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7805__C _1132_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6598_ core_0.execute.rf.reg_outputs\[7\]\[1\] _2941_ _1978_ _2947_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_230_3274 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_103_247 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8337_ _0513_ clknet_leaf_11_i_clk core_0.dec_pc_inc vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5549_ core_0.execute.mem_stage_pc\[8\] _1957_ _1964_ _1970_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_197_72 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8268_ _0444_ clknet_leaf_21_i_clk core_0.execute.sreg_irq_flags.o_d\[2\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_output156_I net156 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7219_ _3405_ _0384_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_217_115 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8199_ _0375_ clknet_leaf_1_i_clk core_0.execute.alu_mul_div.div_res\[8\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__4140__A1 core_0.ew_reg_ie\[4\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7209__A2 _3391_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4140__B2 core_0.ew_reg_ie\[5\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_232_107 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_226_671 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_21_Left_268 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_198_523 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6968__A1 _1652_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_702 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_713 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_216_68 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_198_567 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_186_729 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_17_719 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5640__A1 _1758_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_240_173 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_185_206 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7268__B _1736_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_56_418 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_56_429 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_232_34 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7393__A1 _1980_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4471__I _1063_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_138_177 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_232_78 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5943__A2 _2264_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_153 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3954__A1 _0539_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_153_136 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_30_Left_277 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_92_782 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_646 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_51_123 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_24_348 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_156 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8137__CLK clknet_leaf_99_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_51_189 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_20_521 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7448__A2 _3546_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_543 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_103_792 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_166_2501 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_205_822 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_189_534 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_220_803 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7620__A2 _3732_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_88_1569 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_35_66 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_59_212 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_189_578 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5631__A1 _1761_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_204_387 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6861__I _0722_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4920_ _1196_ _1201_ _1383_ _1384_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and3_1
XANTENNA__4985__A3 core_0.dec_l_reg_sel\[0\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_129_111 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_185_740 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_clkbuf_leaf_113_i_clk_I clknet_4_4__leaf_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_118_807 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_142_34 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4851_ _0914_ _1306_ _1338_ _0083_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__6187__A2 net206 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7384__A1 _0720_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_177_2641 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_191_209 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5234__I1 net204 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_136_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_145_615 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_184_261 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_157_486 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7570_ _3675_ _3691_ _3692_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_4782_ _1290_ _1295_ _0057_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_27_131 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_27_142 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_117_339 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3945__A1 _0576_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_172_445 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6521_ _1381_ core_0.execute.sreg_irq_pc.o_d\[15\] _2898_ _2899_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__6810__B _3072_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_144_169 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_43_646 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_160_629 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_125_361 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6452_ _1380_ core_0.execute.sreg_irq_pc.o_d\[13\] _2831_ _2832_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_70_465 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_99_1698 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_5403_ _1375_ _1845_ _1846_ _1822_ _1847_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_42_189 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_30_329 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_113_556 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6383_ _2764_ _0189_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_113_589 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4370__A1 core_0.fetch.prev_request_pc\[11\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_8122_ _0298_ clknet_4_7__leaf_i_clk core_0.execute.rf.reg_outputs\[3\]\[13\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_2_275 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5145__C _1531_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5334_ _1759_ _1780_ _1781_ _1782_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_140_397 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_208_3007 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_188_2770 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_8053_ _0229_ clknet_leaf_106_i_clk core_0.execute.rf.reg_outputs\[7\]\[8\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5265_ core_0.decode.oc_alu_mode\[12\] _1714_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__inv_2
XANTENNA__5940__I _0799_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_110_1832 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_38_i_clk_I clknet_4_11__leaf_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_76_62 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4122__A1 core_0.execute.pc_high_out\[7\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7004_ _1637_ _3178_ _3220_ _3177_ _3221_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_4216_ net50 core_0.fetch.out_buffer_data_instr\[20\] _0723_ _0835_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__5170__I0 net101 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_242_405 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5196_ core_0.execute.rf.reg_outputs\[6\]\[1\] _1435_ _1436_ core_0.execute.rf.reg_outputs\[4\]\[1\]
+ core_0.execute.rf.reg_outputs\[3\]\[1\] _1443_ _1645_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi222_2
XFILLER_0_214_107 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_208_660 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_126_2028 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5870__A1 _1196_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4147_ core_0.dec_used_operands\[0\] _0766_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_211_814 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4078_ core_0.execute.rf.reg_outputs\[1\]\[1\] _0700_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XANTENNA__5622__A1 _1715_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_78_521 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_222_173 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_167_206 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_203_2951 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_7906_ _0097_ clknet_leaf_68_i_clk core_0.decode.i_imm_pass\[15\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_211_858 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_195_526 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_195_559 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_174_Right_174 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_219_3136 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_210_379 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7837_ _0030_ clknet_leaf_72_i_clk core_0.fetch.out_buffer_data_instr\[14\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_176_751 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6178__A2 _2547_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_121_1961 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4189__A1 core_0.execute.alu_mul_div.comp vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_108_317 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7768_ core_0.decode.i_instr_l\[8\] core_0.decode.i_instr_l\[7\] _3842_ _3843_ vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_0_148_497 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_451 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_19_665 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_93_579 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_191_743 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_190_220 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_135_136 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6719_ _2972_ _3021_ _3030_ _0259_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__7127__A1 _2797_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_135_158 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_137_2157 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_22_777 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_7699_ _1135_ _3792_ _3793_ _3798_ _3799_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_0_18_197 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_151_629 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7678__A2 _1092_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_6_581 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_34_679 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_116_383 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_150_139 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_150_2313 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_33_178 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_132_865 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_131_342 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_131_375 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4361__A1 _0972_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_30_863 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_218_413 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_246_744 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6102__A2 _2254_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_218_457 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4113__A1 core_0.execute.pc_high_out\[3\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_243_3432 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6167__B _1458_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4664__A2 _1051_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_148_2286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_199_832 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_161_2442 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5613__A1 _1479_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_243_22 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_69_587 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_141_Right_141 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_201_379 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6169__A2 _1613_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_173_209 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_139_464 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_126_103 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5916__A2 _1585_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_154_434 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_181_220 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_112_37 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_484 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7118__A1 _1372_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_181_253 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_181_275 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_52_443 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_107_361 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7669__A2 _1084_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_156 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_172_2571 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_172_2582 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_24_167 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_24_189 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_97_39 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_110_504 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_236_243 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5050_ _1496_ _1497_ _1498_ _1499_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_0_224_405 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_224_416 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4001_ _0627_ _0594_ _0628_ _0629_ _0630_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai211_4
Xclkbuf_leaf_62_i_clk clknet_4_14__leaf_i_clk clknet_leaf_62_i_clk vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_205_685 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_204_162 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6591__I _2935_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_88_863 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5952_ _2244_ _2334_ _2343_ _2242_ _2344_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai211_1
Xclkbuf_leaf_77_i_clk clknet_4_13__leaf_i_clk clknet_leaf_77_i_clk vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_4903_ _1225_ _1369_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_220_688 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87_384 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_153_88 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_749 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7357__A1 _2711_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8302__CLK clknet_leaf_12_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5883_ _2242_ _0720_ _2275_ _2276_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_47_1074 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_7622_ _0736_ _3733_ _3737_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_185_570 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4834_ _1280_ net41 _1170_ _1326_ _1327_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_0_185_592 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_451 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_60_1230 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7636__B _1216_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_28_473 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7553_ core_0.execute.pc_high_buff_out\[0\] _3676_ _3670_ _3677_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__7109__A1 _3189_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4765_ _1284_ _1286_ _0049_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_55_270 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_145_467 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_117_169 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_145_489 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_16_657 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6504_ _2294_ _2730_ _2090_ _2882_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_43_454 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_126_681 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_214_3077 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_16_679 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_70_240 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7484_ _3514_ _3628_ _3632_ _0422_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_4696_ _1245_ _0021_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_70_251 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_167 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_30_104 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_125_191 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_540 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6435_ _1684_ _1480_ _2815_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_114_865 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_3_562 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6332__A2 _1114_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_15_i_clk clknet_4_8__leaf_i_clk clknet_leaf_15_i_clk vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__4343__A1 _0947_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_12_863 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6366_ _1433_ core_0.execute.alu_mul_div.mul_res\[11\] _2748_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_TAPCELL_ROW_132_2098 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_87_72 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_101_559 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8105_ _0281_ clknet_leaf_95_i_clk core_0.execute.rf.reg_outputs\[4\]\[12\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5317_ _1461_ net187 _1764_ _1765_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_4
XANTENNA__6766__I _1963_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_227_221 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6297_ _2311_ _2642_ _2680_ _2681_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__6096__A1 _2346_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_8036_ _0213_ clknet_leaf_82_i_clk core_0.ew_reg_ie\[3\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__dffq_2
XPHY_EDGE_ROW_243_Right_243 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
X_5248_ _1124_ _1696_ _1697_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_input32_I i_mem_data[5] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_71_1370 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4286__I core_0.fetch.prev_request_pc\[6\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_215_438 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_215_449 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_194_84 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5179_ core_0.execute.rf.reg_outputs\[4\]\[5\] _1436_ _1437_ core_0.execute.rf.reg_outputs\[2\]\[5\]
+ _1628_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_0_199_139 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_223_460 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7596__A1 _3663_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6399__A2 _2777_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_223_471 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_97_137 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output119_I net119 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_27_836 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_97_159 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_195_334 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5111__S _1559_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_66_524 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_78_384 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7348__A1 _1719_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_183_507 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_535 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_155_209 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_94_855 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_109_615 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_38_259 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_136_412 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_149_795 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_54_719 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6020__A1 _2300_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3909__A1 _0539_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_47_782 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_191_562 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4582__A1 core_0.ew_data\[5\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_163_286 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_105_832 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_123_139 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_22_616 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_22_627 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_104_Left_351 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_120_802 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7520__A1 _0626_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_131_150 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4334__A1 core_0.fetch.prev_request_pc\[9\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7281__B _1395_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_219_722 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4885__A2 _1285_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6676__I _2998_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_218_232 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_219_788 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_206_405 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_246_574 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_210_Right_210 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_7_594 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5834__A1 _2202_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_233_257 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_221_408 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_113_Left_360 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_233_279 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7587__A1 net204 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_202_622 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_85_1528 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_199_684 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_186_301 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_340 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5062__A2 net180 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_85_822 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7339__A1 _2183_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4270__B1 _0854_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_202_699 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_546 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_32_34 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_174_2600 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_45_719 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_72_505 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6011__A1 core_0.dec_sreg_irt vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_72_527 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_32_89 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_154_242 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_154_253 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_25_443 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_681 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_4550_ _1132_ _1133_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_52_251 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_571 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_424 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_115 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6314__A2 _2695_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4481_ _1066_ _1073_ _1074_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_52_295 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_96_1668 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4325__A1 _0725_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6220_ _1107_ _2590_ _2601_ _2605_ _2606_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XFILLER_0_40_457 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_110_301 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_4_5__f_i_clk clknet_3_2_0_i_clk clknet_4_5__leaf_i_clk vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__4876__A2 _1341_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5704__B net211 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_682 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6586__I _2935_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6151_ net84 _2531_ _2536_ _2537_ _2538_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_20_170 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6078__A1 _2300_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_209_243 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5102_ _1467_ net178 _1551_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_6082_ _1831_ _2470_ _1684_ _2471_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_225_736 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4628__A2 core_0.execute.alu_flag_reg.o_d\[0\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5033_ _1481_ _1482_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_225_758 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_240_706 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_240_717 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_212_408 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_79_104 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_224_279 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_49_1103 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_178_802 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7578__A1 _3675_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6984_ core_0.execute.alu_mul_div.cbit\[1\] _3199_ _3200_ _3201_ _3202_ vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai31_2
XFILLER_0_76_800 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_200_2910 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_189_194 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_94_107 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_220_452 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_502 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5053__A2 _1501_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_24_806 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_48_524 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5935_ _1480_ _2311_ _2326_ _1684_ _2327_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XFILLER_0_48_535 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_192_304 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_76_855 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_105_1775 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_87_192 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_165_529 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_216_3106 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_5866_ core_0.execute.pc_high_out\[0\] _2257_ _2258_ net106 _2259_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_35_207 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_63_516 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6002__A1 _2346_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_118_445 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7605_ core_0.execute.pc_high_out\[7\] _3722_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_90_313 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_173_540 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4817_ core_0.decode.i_instr_l\[7\] _1315_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__inv_1
XANTENNA__7842__CLK clknet_leaf_67_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_7_142 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_63_549 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_161_702 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_173_562 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_44_730 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5797_ _2195_ _2196_ _2197_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6553__A2 _2783_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_44_741 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_629 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7750__B2 _3827_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_32_894 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4564__A1 _0727_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_134_2116 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_7536_ _0730_ _3664_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_4748_ net58 _1241_ _1275_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_7_197 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_102_802 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7467_ core_0.execute.sreg_irq_pc.o_d\[14\] _3542_ _3619_ _3620_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_43_295 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_98_71 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6305__A2 _1117_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4679_ _1221_ _1234_ _0015_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__7502__A1 _3514_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_1_Right_1 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_113_150 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6418_ _1088_ _2797_ _2798_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_141_492 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7398_ _3543_ _3561_ _3562_ _0406_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_12_671 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_101_356 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6349_ _2294_ _2730_ _2731_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_101_367 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3913__I _0548_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_101_378 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_227_3235 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6069__A1 _2244_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5106__S _1554_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_216_703 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7805__A2 _3788_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4619__A2 core_0.execute.alu_flag_reg.o_d\[1\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_8019_ _0196_ clknet_leaf_31_i_clk net123 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_208_69 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_4_564 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4095__A3 _0544_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_145_2256 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_215_279 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_203_419 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7569__A1 core_0.execute.pc_high_buff_out\[2\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_98_435 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_98_446 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_98_457 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6241__A1 _1693_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_671 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5044__A2 _1438_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_195_142 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_85_129 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_168_367 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_78_181 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6792__A2 _3070_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_238_3364 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_7_i_clk_I clknet_4_2__leaf_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_183_326 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_137_732 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_376 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_81_313 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_80_1469 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_240_34 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_35_752 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_81_368 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_151_212 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_136_297 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_156_2385 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_50_711 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_640 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_722 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_50_733 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7344__I1 _2888_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4307__A1 core_0.fetch.prev_request_pc\[15\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_457 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4307__B2 core_0.fetch.prev_request_pc\[14\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_132_492 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4858__A2 _1306_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_206_213 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5807__A1 core_0.execute.rf.reg_outputs\[1\]\[2\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_207_769 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_118_58 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_89_413 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_222_728 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_221_216 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_215_780 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_180_2670 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_215_791 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_77_619 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_159_323 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_199_492 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_89_479 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_76_107 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5035__A2 _0767_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_202_452 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6232__B2 net15 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_186_142 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_175_805 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3981_ _0568_ _0535_ _0536_ core_0.execute.rf.reg_outputs\[2\]\[10\] _0612_ vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_0_147_518 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_175_827 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_66 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_58_855 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6783__A2 _3064_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_187_698 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5720_ _2119_ _2120_ _1554_ _2121_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__4794__A1 core_0.fetch.prev_request_pc\[14\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_44_1044 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_57_376 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_72_313 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7186__B core_0.execute.alu_mul_div.div_res\[12\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
X_5651_ _2051_ _2052_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_150_34 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_216_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_4602_ core_0.ew_data\[7\] core_0.ew_data\[15\] _1150_ _1166_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_4_101 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_72_357 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4546__A1 core_0.decode.oc_alu_mode\[13\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_115_426 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_170_521 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_5_646 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_519 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5582_ _1051_ _1953_ _1984_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_25_251 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_143_768 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7321_ core_0.execute.alu_flag_reg.o_d\[0\] _3494_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_4533_ _1056_ _1068_ _1069_ _1119_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_4
XTAP_TAPCELL_ROW_211_3047 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_7252_ _1414_ core_0.execute.sreg_irq_pc.o_d\[7\] _1410_ _1431_ _1736_ _3434_ vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_0_111_621 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4464_ _1055_ _1049_ _1057_ _1058_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_111_632 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_123_492 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_7_66 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4849__A2 _1306_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6203_ _2157_ _2550_ _2589_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_40_298 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_111_665 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7183_ _2714_ _3376_ _3357_ _0377_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_4395_ net84 _1004_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XTAP_TAPCELL_ROW_55_1173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6134_ core_0.execute.alu_mul_div.i_mul core_0.execute.alu_mul_div.mul_res\[5\] _2522_
+ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_EDGE_ROW_209_Left_456 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
X_6065_ _1378_ _2452_ _2453_ _2454_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_84_51 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5016_ _0714_ _0715_ _0716_ _0717_ _1465_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_0_225_588 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_1_523 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_222_3176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_212_238 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_205_290 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_68_619 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_177_120 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_221_761 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_37_953 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6223__A1 core_0.execute.alu_mul_div.div_res\[7\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5026__A2 core_0.execute.alu_flag_reg.o_d\[1\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_822 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_177_131 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_177_142 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6967_ _3180_ _3154_ _3186_ _3187_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor3_1
XANTENNA__6774__A2 _3043_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_48_332 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_140_2197 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_5918_ net224 _2309_ _2310_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__4785__B2 net162 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_194_2839 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7808__C _1279_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_177_197 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_193_657 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6898_ _2951_ _3129_ _3133_ _0335_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XPHY_EDGE_ROW_218_Left_465 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_193_679 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_527 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_48_387 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_76_696 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_324 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_192_167 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_180_307 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5849_ _2241_ _2242_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XANTENNA__3908__I _0543_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_90_121 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_106_404 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_118_275 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4537__A1 _1034_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_133_212 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_16_240 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_91_699 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_210_37 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_44_582 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_118_1933 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_7519_ core_0.execute.sreg_scratch.o_d\[9\] _3646_ _3651_ _3655_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA_output186_I net186 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_133_278 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_114_470 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_114_492 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_9_623 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_101_142 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_102_687 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_227_Left_474 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA_clkbuf_leaf_86_i_clk_I clknet_4_12__leaf_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_244_853 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4068__A3 _0543_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6462__A1 _2090_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_235_34 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7888__CLK clknet_leaf_83_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_235_78 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_169_632 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6214__A1 _1059_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_107 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6214__B2 _1620_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_211_282 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6765__A2 _3043_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_157_838 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_158_2403 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_236_Left_483 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_67_652 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_158_2414 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_104_27 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4776__A1 _1290_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_156_348 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_836 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_39_398 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_55_858 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_82_633 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_125_702 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4423__B _0970_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6517__A2 _1386_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_109_264 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_109_275 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_89_18 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4528__A1 _1034_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_70_839 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7190__A2 _3372_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4142__C _0539_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_120_26 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_120_37 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_152_587 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_93_1627 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_10_405 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_50_574 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_492 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_238_102 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_416 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_245_Left_492 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__4649__I _1206_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_169_2543 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_226_308 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4161__C1 core_0.ew_reg_ie\[1\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4180_ _0798_ _0799_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__inv_4
XFILLER_0_235_842 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6864__I _3106_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_207_555 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_207_566 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_207_599 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_145_34 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_54_32 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_166_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_7870_ _0062_ clknet_leaf_63_i_clk core_0.fetch.prev_request_pc\[13\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_145_78 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_203_772 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6821_ _2946_ _3086_ _3089_ _0302_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_159_142 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_148_816 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_202_271 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_34_923 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6756__A2 _3049_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_9_204 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6813__B _3083_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4767__A1 _1284_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_46_803 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6752_ core_0.execute.rf.reg_outputs\[4\]\[4\] _3049_ _3045_ _3050_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_9_226 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3964_ _0533_ core_0.execute.rf.reg_outputs\[4\]\[11\] net230 _0596_ vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_0_85_460 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_92_419 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_102_1734 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_161_66 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5703_ _1123_ _1637_ net211 _1720_ _2104_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_0_175_679 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6683_ core_0.execute.rf.reg_outputs\[6\]\[7\] _3006_ _3004_ _3010_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_73_644 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_161_88 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_45_346 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_70_86 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3895_ core_0.execute.rf.reg_outputs\[7\]\[15\] _0530_ _0531_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_14_680 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4519__A1 _1034_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_508 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5634_ _1579_ _1584_ _2035_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_115_212 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3990__A2 _0524_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_5_432 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_699 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8193__CLK clknet_leaf_2_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7644__B _1216_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_115_267 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_143_576 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5565_ core_0.execute.mem_stage_pc\[15\] _1955_ _1978_ _1979_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_103_418 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_57_1202 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_170_384 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7304_ _2859_ _3391_ _3479_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_5_498 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_124_790 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4516_ _1097_ _1100_ _1102_ _1105_ _1106_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor4_4
X_8284_ _0460_ clknet_leaf_29_i_clk core_0.execute.pc_high_buff_out\[5\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5496_ _1632_ _1636_ _1929_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_0_111_440 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7235_ _3416_ _3419_ _1395_ _0386_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_4447_ _1038_ _1039_ _1041_ _1042_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_0_111_473 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_108_i_clk_I clknet_4_5__leaf_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6692__A1 _2988_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_113_1863 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_113_1874 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_7166_ _3358_ _3365_ core_0.execute.alu_mul_div.div_res\[4\] _3366_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_224_3205 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_4378_ _0987_ _0966_ _0989_ _0990_ _0963_ net162 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_0_95_72 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6117_ _2502_ _2504_ _2505_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_129_2059 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_7097_ core_0.execute.alu_mul_div.mul_res\[10\] _3285_ _3300_ core_0.execute.alu_mul_div.mul_res\[11\]
+ _3306_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_225_352 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5247__A2 _1558_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6444__A1 core_0.execute.alu_mul_div.div_res\[13\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
X_6048_ core_0.execute.alu_mul_div.div_res\[3\] _1114_ _2435_ _2437_ _1432_ _2438_
+ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_0_241_834 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_142_2215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4455__B1 _1044_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_197_226 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_68_1331 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_206_2982 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_96_714 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6747__A2 _3043_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6723__B _3031_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7999_ _0176_ clknet_leaf_119_i_clk net138 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_178_473 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output101_I net101 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_193_410 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_166_635 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4758__A1 _0727_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_178_495 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_95_279 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_235_3334 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_76_493 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_193_476 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_37_858 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_9_760 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_107_702 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_119_562 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_180_115 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_357 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3981__A2 _0535_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_106_223 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_52_839 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_64_699 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_134_543 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_176 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_768 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_187 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_91_496 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_153_2344 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_162_863 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5183__A1 net98 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_51_349 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_134_587 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5853__I net187 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_79_1460 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_161_373 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_121_248 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_32_585 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6683__A1 core_0.execute.rf.reg_outputs\[6\]\[7\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5486__A2 _1501_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_246_3463 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_246_3474 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_217_864 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_188_Right_188 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__5238__A2 _1469_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_204_514 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5521__C _1950_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_246_88 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_164_2484 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6986__A2 _3202_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_188_226 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_188_237 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_86_224 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_212_580 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6738__A2 _3022_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_156_101 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_200_753 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5946__B1 _2260_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_129_337 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_129_348 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_156_134 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_95_780 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5410__A2 _1814_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_41_1003 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4153__B _0771_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_54_132 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_156_189 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_40_34 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_43_828 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3972__A2 _0602_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_125_532 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7903__CLK clknet_leaf_68_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_54_165 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_131_69 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7163__A2 _1362_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_699 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_11_650 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5174__A1 _1531_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_42_349 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6910__A2 _3129_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5350_ core_0.execute.alu_mul_div.div_cur\[13\] _1798_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_2
Xoutput205 net205 sr_bus_data_o[5] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_2_457 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_239_422 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4379__I net87 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4301_ _0911_ _0918_ _0919_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_11_747 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_49_54 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5281_ _1430_ net194 _1730_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_11_769 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_227_617 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5477__A2 _1620_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_10_257 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7020_ _3222_ _3228_ _3235_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or2_1
X_4232_ _0824_ net45 _0850_ _0851_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_4
XTAP_TAPCELL_ROW_52_1132 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6808__B _3072_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_4_34 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_242_609 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4163_ _0781_ _0782_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XPHY_EDGE_ROW_155_Right_155 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__5229__A2 _1665_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_241_119 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_235_672 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_64 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_222_311 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4328__B _0945_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_207_385 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4094_ core_0.execute.rf.reg_outputs\[7\]\[0\] _0530_ _0715_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6977__A2 _2322_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_222_333 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4988__A1 _0770_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7922_ _0000_ clknet_leaf_8_i_clk core_0.execute.alu_mul_div.i_mod vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_179_237 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7853_ _0046_ clknet_leaf_64_i_clk core_0.fetch.out_buffer_data_instr\[30\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_81_41 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6729__A2 _3027_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_148_613 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_77_257 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6804_ core_0.execute.rf.reg_outputs\[3\]\[11\] _3070_ _3072_ _3079_ vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_77_279 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7784_ _1136_ _3853_ _0501_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_4996_ core_0.dec_l_reg_sel\[2\] core_0.dec_l_reg_sel\[1\] core_0.dec_l_reg_sel\[0\]
+ _1445_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_0_147_134 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_19_836 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5401__A2 _1715_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_92_227 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_148_679 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_191_2809 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6735_ core_0.execute.rf.reg_outputs\[5\]\[14\] _3020_ _3031_ _3039_ vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3947_ _0580_ net198 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA_clkbuf_leaf_34_i_clk_I clknet_4_11__leaf_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_858 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_63_1272 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_73_430 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_135_318 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3963__A2 _0530_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6666_ _2998_ _3000_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_190_457 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_46_699 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_34_839 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4998__B _1446_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_60_102 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_636 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_144_863 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_162_159 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_73_496 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7374__B _0731_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5617_ _2017_ _1619_ _2018_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_2
XANTENNA__5165__B2 core_0.execute.rf.reg_outputs\[7\]\[7\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
X_6597_ _2930_ core_0.ew_data\[1\] _2945_ _2946_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_4
XFILLER_0_131_513 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_230_3275 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4912__A1 _1223_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_8336_ _0512_ clknet_leaf_118_i_clk core_0.dec_r_bus_imm vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_170_181 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5548_ _1968_ _1172_ _1969_ _1950_ _0149_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA_clkbuf_3_3_0_i_clk_I clknet_0_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input62_I i_req_data[31] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4289__I _0836_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_112_771 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8267_ _0443_ clknet_leaf_21_i_clk core_0.execute.sreg_irq_flags.o_d\[1\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5479_ _1909_ _1585_ _1912_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_112_782 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5468__A2 _1817_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7218_ _3384_ _3404_ _3405_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
X_8198_ _0374_ clknet_leaf_3_i_clk core_0.execute.alu_mul_div.div_res\[7\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__6718__B _3016_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_10_791 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7149_ _3342_ _3177_ _3352_ _3354_ _0365_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__4140__A2 _0520_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output149_I net149 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8089__CLK clknet_leaf_99_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_122_Right_122 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_232_119 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_214_823 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_198_502 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6968__A2 _3178_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4979__B2 _1390_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_198_579 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_69_758 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5848__I core_0.dec_mem_access vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_178_281 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_37_600 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_68_279 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_205 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_166_454 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_139_679 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_166_465 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_138_189 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_193_284 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_193_295 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_37_677 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_147_690 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_52_614 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_37_699 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5156__A1 _0770_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_162_671 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_10_37 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_122_524 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_134_384 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_166_2502 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_20_588 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_236_436 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6628__B _2971_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4131__A2 _0748_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4927__I _1390_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_223_119 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_217_694 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_216_171 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_204_311 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7081__A1 _2053_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_87_500 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_220_815 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7459__B _3553_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5631__A2 _2019_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_206_91 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_185_730 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_408 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_59_279 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4850_ core_0.decode.i_imm_pass\[1\] _1307_ _1338_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_177_2631 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7384__A2 _3544_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_177_2642 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_184_240 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5395__A1 core_0.execute.alu_mul_div.div_cur\[3\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
X_4781_ core_0.fetch.prev_request_pc\[8\] _1285_ _0880_ net175 _1295_ vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_0_145_627 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_172_413 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_51_66 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_157_498 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_129_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6520_ _1380_ _2897_ _2898_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_145_649 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3945__A2 _0578_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_83_772 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_16_839 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_55_474 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_172_457 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_42_102 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_70_411 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_222_90 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_496 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_126_863 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6451_ _1380_ _2830_ _2831_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__5707__B net211 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_42_157 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_113_524 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5402_ _1374_ _1836_ _1846_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_99_1699 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6895__A1 net95 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_224_Right_224 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_152_181 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6382_ core_0.ew_data\[11\] _2763_ _2190_ _2764_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_2_243 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8121_ _0297_ clknet_leaf_99_i_clk core_0.execute.rf.reg_outputs\[3\]\[12\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_2_265 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5333_ core_0.execute.alu_mul_div.div_cur\[7\] _1758_ _1781_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_11_555 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_140_387 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_208_3008 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_188_2771 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_8052_ _0228_ clknet_leaf_115_i_clk core_0.execute.rf.reg_outputs\[7\]\[7\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_2
X_5264_ _1712_ _1713_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_11_599 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_227_436 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_110_1833 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_7003_ _3214_ _3218_ _3219_ _3220_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_4215_ _0823_ _0827_ _0830_ _0833_ _0834_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and4_1
X_5195_ _1558_ _1553_ _1644_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_76_96 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_242_439 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4146_ _0759_ _0761_ _0762_ _0763_ _0764_ _0765_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XTAP_TAPCELL_ROW_126_2029 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_223_620 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7072__A1 _1224_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_207_193 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_223_653 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_222_130 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4077_ _0699_ net202 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XANTENNA__5622__A2 _1934_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_92_73 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_203_2952 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_7905_ _0096_ clknet_leaf_69_i_clk core_0.decode.i_imm_pass\[14\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_222_185 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_92_95 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_222_196 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_195_549 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_159_Left_406 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
X_7836_ _0029_ clknet_leaf_82_i_clk core_0.fetch.out_buffer_data_instr\[13\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_219_3137 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_59_780 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_148_443 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_148_454 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_148_465 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_176_774 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5386__A1 core_0.execute.alu_mul_div.div_cur\[3\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_121_1962 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4189__A2 _0804_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7767_ _3783_ _3837_ _3838_ _3841_ _3842_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and4_2
X_4979_ core_0.execute.sreg_priv_control.o_d\[15\] _1393_ _1428_ _1390_ _1429_ vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_190_210 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_830 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_18_154 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6718_ core_0.execute.rf.reg_outputs\[5\]\[6\] _3027_ _3016_ _3030_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__3936__A2 _0528_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7127__A2 _3181_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7698_ _1055_ _1094_ _3796_ _3797_ _3798_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XTAP_TAPCELL_ROW_137_2158 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_22_778 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_151_619 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5138__A1 _0789_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_124 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_150_107 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6649_ _2979_ core_0.ew_data\[11\] _2980_ net23 _2988_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XANTENNA__6335__B1 _2577_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_658 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_33_146 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_144_693 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_6_593 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_466 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_150_2314 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_33_168 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_116_395 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_21_319 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_132_855 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_42_680 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_371 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_76_1430 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_104_579 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_131_365 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4361__A2 _0966_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_8319_ _0495_ clknet_leaf_11_i_clk core_0.dec_jump_cond_code\[4\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_2
XPHY_EDGE_ROW_168_Left_415 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__5310__A1 _1513_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_246_778 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_243_3433 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_245_266 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_205_108 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_205_119 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_148_2287 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7063__A1 _1909_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6962__I _3173_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_161_2443 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_214_664 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_202_815 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_186_505 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5613__A2 _1665_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_241_483 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_213_174 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_97_842 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_EDGE_ROW_177_Left_424 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_213_185 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_202_859 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_198_387 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_186_527 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_69_555 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_213_196 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_243_56 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_29_419 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_69_599 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_167_752 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7366__A2 _3533_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_56_238 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8104__CLK clknet_leaf_109_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5377__A1 _1748_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_194_582 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_290 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6911__B _3139_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_182_733 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_772 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_64_260 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_154_457 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7118__A2 _3324_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_108_863 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5129__A1 _1482_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7669__A3 _1072_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_172_2572 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_181_298 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_122_310 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_135_693 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8254__CLK clknet_leaf_24_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_52_477 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_186_Left_433 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_21_842 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_122_387 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6629__A1 core_0.execute.rf.reg_outputs\[7\]\[6\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_236_200 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_237_734 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5301__A1 core_0.execute.alu_mul_div.div_cur\[15\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_236_255 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_209_469 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4000_ _0565_ core_0.execute.rf.reg_outputs\[4\]\[8\] _0520_ _0629_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_0_46_55 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_88 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_204_130 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_195_Left_442 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_79_319 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6801__A1 _2983_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_204_174 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5951_ _2272_ _2271_ _2342_ _2343_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_204_196 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_246_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87_352 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_177_549 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_220_667 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4902_ _1367_ _1231_ _1368_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_5882_ _2241_ _2274_ _2275_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_47_1075 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_75_547 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7621_ _3732_ _3735_ _3736_ _0455_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__5368__A1 _1232_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_157_262 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4833_ _1280_ _1255_ _1326_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_118_649 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_172_221 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7552_ _0732_ _1206_ _3676_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_2
XTAP_TAPCELL_ROW_60_1231 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_145_446 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4764_ core_0.fetch.prev_request_pc\[0\] _1285_ _0881_ net161 _1286_ vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_0_173_766 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_71_720 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_43_422 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6503_ _2123_ _2808_ _2880_ _2113_ _2881_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XFILLER_0_55_282 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5437__B _1817_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_132_107 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_753 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7483_ core_0.execute.sreg_jtr_buff.o_d\[2\] _3628_ _3384_ _3632_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4695_ core_0.fetch.out_buffer_data_instr\[5\] net65 _1241_ _1245_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_172_287 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_214_3078 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_113_310 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_126_693 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_43_477 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6868__A1 _2967_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6434_ _2072_ _2073_ _2814_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_102_93 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_113_332 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7652__B _1217_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6365_ _2734_ _2746_ _2747_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_23_190 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_141_696 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_11_352 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8104_ _0280_ clknet_leaf_109_i_clk core_0.execute.rf.reg_outputs\[4\]\[11\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_132_2099 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_11_363 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5316_ _1461_ net213 _1764_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_53_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6296_ _1109_ _2163_ _2036_ core_0.decode.oc_alu_mode\[6\] _2679_ _2680_ vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XANTENNA__6096__A2 net204 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7293__A1 _1430_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_8035_ _0212_ clknet_leaf_82_i_clk core_0.ew_reg_ie\[2\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__dffq_4
X_5247_ _1479_ _1558_ _1553_ _1641_ _1696_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor4_4
XTAP_TAPCELL_ROW_71_1360 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5843__A2 _2231_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5178_ core_0.execute.rf.reg_outputs\[1\]\[5\] _1615_ _1434_ core_0.execute.rf.reg_outputs\[6\]\[5\]
+ _1627_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XANTENNA_input25_I i_mem_data[13] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_242_247 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7045__A1 _2587_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_230_409 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4129_ core_0.execute.pc_high_out\[5\] _0732_ _0748_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_79_820 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_223_483 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_79_842 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_168_527 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_27_837 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_211_667 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5071__A3 _1517_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_211_689 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_210_166 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7348__A2 _2888_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_210_177 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_66_547 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_38_249 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_109_627 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7819_ _1461_ _1134_ _3758_ _3877_ _1283_ _0512_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XANTENNA__6731__B _3031_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_108_104 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_136_424 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6020__A2 _2409_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_452 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8277__CLK clknet_leaf_26_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3909__A2 _0542_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_163_232 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4031__A1 net100 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_485 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_411 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_720 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_159 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_151_405 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4582__A2 net157 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_606 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6859__A1 core_0.execute.rf.reg_outputs\[1\]\[2\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_488 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output93_I net93 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_15_680 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_132_663 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7520__A2 _3640_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_61_296 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5531__A1 _1024_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_30_650 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4885__A3 _0883_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_238_34 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_3_i_clk_I clknet_4_2__leaf_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7284__A1 _1742_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_219_767 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_218_266 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4098__A1 net88 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_218_277 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_234_737 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_7_595 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6906__B _3124_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_233_269 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7587__A2 _3675_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_85_1529 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_199_696 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_187_836 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_201_133 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_187_858 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_186_335 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_352 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_202_667 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_97_672 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_186_346 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_216 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4270__A1 core_0.fetch.prev_request_pc\[12\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_201_166 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_97_694 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7339__A2 _3502_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4270__B2 core_0.fetch.prev_request_pc\[11\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_174_519 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_139_251 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_57_558 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_127_402 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_139_273 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_174_2601 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_84_355 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_366 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6011__A2 _2400_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_155_766 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_37_282 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_142_405 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_660 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_114_107 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_142_438 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_488 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_583 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4480_ _1040_ _1045_ _1073_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_0_80_594 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_96_1669 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7472__B _3541_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4588__S net157 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_110_313 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_111_836 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_122_173 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_111_858 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6150_ _2245_ _2537_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_21_694 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_148_34 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7275__A1 net73 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_196_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_185_2730 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6078__A2 _1560_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5101_ _1531_ _1549_ _1550_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_209_255 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6081_ _2468_ _2469_ _2470_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5032_ _1462_ _1469_ _1481_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_4
XANTENNA__6308__S _2242_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_240_729 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_49_1104 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_164_66 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6983_ _3183_ _3184_ core_0.execute.alu_mul_div.cbit\[1\] _3201_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_200_2911 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6250__A2 _2161_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_73_97 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_88_672 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5934_ _1831_ _2319_ _2325_ _2326_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and3_1
XANTENNA__5011__I _1459_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4261__A1 _0722_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_177_368 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_105_1776 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7647__B _3731_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_216_3107 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_192_327 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5865_ _1382_ _1196_ _1201_ _2252_ _2258_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and4_2
XTAP_TAPCELL_ROW_196_2870 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_192_338 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_8_622 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6002__A2 net221 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7604_ _3663_ _3721_ _0453_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_4816_ _1314_ _0072_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_29_772 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_145_232 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_260 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_118_457 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_63_539 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5796_ _2187_ _2194_ _2196_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__7750__A2 _3766_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_7_165 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_145_276 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4747_ _0852_ _1238_ _1274_ _0043_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_43_230 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_32_895 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_7535_ _1283_ _3663_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XTAP_TAPCELL_ROW_134_2117 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_173_596 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_161_769 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7466_ _0563_ _3546_ _3541_ _3618_ _3619_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_4678_ _0804_ _1233_ _1234_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_31_436 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7502__A2 _3640_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6417_ core_0.execute.alu_mul_div.mul_res\[13\] _2797_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__inv_2
XFILLER_0_98_83 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_458 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_98_94 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_141_471 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7397_ core_0.execute.sreg_irq_pc.o_d\[2\] _3542_ _3516_ _3562_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_113_184 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6348_ _2729_ _2668_ _2123_ _2730_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_12_694 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_171 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_227_3236 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6279_ _2661_ _2662_ _2624_ _2663_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_228_597 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_208_37 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_8018_ _0195_ clknet_leaf_24_i_clk net116 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__7018__A1 _3189_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output131_I net131 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5630__B _2022_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_98_403 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_145_2257 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_231_718 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_4_565 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6218__S _2293_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_231_729 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7569__A2 _3682_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_169_858 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4252__A1 _0869_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_66_311 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_195_154 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_536 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_211_486 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_39_547 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_168_379 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_238_3365 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_66_344 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_93_130 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_94_653 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_82_804 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_94_664 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_109_413 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7049__S core_0.execute.alu_mul_div.cbit\[1\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4004__A1 _0565_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_54_539 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_82_i_clk_I clknet_4_13__leaf_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_61_i_clk clknet_4_14__leaf_i_clk clknet_leaf_61_i_clk vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__5752__A1 _1715_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_156_2386 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_62_550 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_22_403 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_151_246 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_151_257 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_151_279 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_22_447 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4307__A2 _0827_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_105_685 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_160_791 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_238_317 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_104_195 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_76_i_clk clknet_4_13__leaf_i_clk clknet_leaf_76_i_clk vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_219_542 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_234_501 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_91_1599 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5807__A2 _1615_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_234_523 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_118_37 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_246_394 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7009__A1 _3183_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5540__B _1964_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6480__A2 _1117_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4935__I _0731_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_180_2671 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_214_280 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_159_335 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6232__A2 _2579_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_230_762 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xclkbuf_leaf_14_i_clk clknet_4_8__leaf_i_clk clknet_leaf_14_i_clk vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_3980_ _0534_ _0542_ _0544_ core_0.execute.rf.reg_outputs\[5\]\[10\] _0611_ vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_4
XANTENNA__4243__A1 _0816_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_171 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_159_368 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_57_322 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_175_839 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5991__A1 _2294_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_128_733 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_152 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_44_1045 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4670__I core_0.execute.alu_mul_div.cbit\[0\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5650_ _1752_ _1567_ _2051_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_0_85_697 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_720 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6090__C _0799_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4601_ _1165_ net144 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xclkbuf_leaf_29_i_clk clknet_4_10__leaf_i_clk clknet_leaf_29_i_clk vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_26_753 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_182_371 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4546__A2 _1062_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5581_ _1983_ _0167_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_25_241 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_111_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_209_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7320_ _3487_ _3492_ _3493_ _0397_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_41_712 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_658 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4532_ _1034_ _1116_ _1118_ _0000_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_211_3048 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_130_419 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_7251_ _2611_ _3391_ _3433_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_41_767 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_244 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4463_ _1041_ _1048_ _1056_ _1057_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_0_13_469 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_1_842 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6202_ _1088_ _2587_ _2588_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_111_644 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_15_Right_15 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
X_7182_ _3361_ _3373_ _3376_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4394_ _0883_ _1002_ _1003_ _0963_ net174 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_4
X_6133_ _2295_ _2501_ _2520_ _2521_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_0_110_187 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_55_1174 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6064_ _1378_ core_0.execute.sreg_irq_pc.o_d\[4\] _2453_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5015_ core_0.execute.rf.reg_outputs\[6\]\[0\] _0661_ _0692_ core_0.execute.rf.reg_outputs\[1\]\[0\]
+ _1463_ _1464_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_0_175_76 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_240_504 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_213_718 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6471__A2 _2642_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_175_87 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_197_419 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_1_524 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6265__C _1432_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_222_3177 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_16_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__7420__A1 _1980_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_37_954 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6223__A2 _2332_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_178_644 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_24_Right_24 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__4234__A1 core_0.fetch.out_buffer_valid vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6966_ _1223_ _3185_ _3186_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_138_508 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_140_2187 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_132_Left_379 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_140_2198 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_178_699 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5917_ _2306_ _2308_ _1603_ _2309_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA_clkbuf_leaf_104_i_clk_I clknet_4_5__leaf_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_76_653 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_64_804 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6897_ net96 _3130_ _3124_ _3133_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_63_303 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_181_809 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_193_669 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_430 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_119_766 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_111 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_118_243 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5848_ core_0.dec_mem_access _2241_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__inv_2
XFILLER_0_75_196 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_17_742 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_119_788 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_161_500 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_133_202 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_146_585 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4537__A2 _1120_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_90_166 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5779_ _1993_ _2178_ _2179_ _2180_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_133_224 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_118_1923 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_90_177 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_118_1934 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_133_246 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_134_769 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_7518_ _0637_ _3640_ _3654_ _0434_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_44_594 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_140_90 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7487__A1 _1217_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_31_244 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_output179_I net179 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7449_ core_0.execute.sreg_irq_pc.o_d\[11\] _3542_ _3604_ _3605_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XPHY_EDGE_ROW_33_Right_33 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_114_482 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_169_Right_169 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_9_624 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_31_277 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_141_290 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_31_288 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_141_Left_388 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_229_862 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7239__A1 net83 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_102_699 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_29_i_clk_I clknet_4_10__leaf_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_244_865 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6462__A2 _2547_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4473__A1 _1065_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_767 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_98_244 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_231_559 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_42_Right_42 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__4691__S _1241_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7411__A1 _1357_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6214__A2 _2018_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6970__I _3176_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_196_441 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_98_288 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_150_Left_397 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_212_784 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_39_322 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_196_474 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_158_2404 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_169_699 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5973__A1 _1601_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_168_198 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_66_174 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_94_494 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_137_552 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_109_254 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7714__A2 _0514_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_70_807 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_82_667 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4528__A2 _1113_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_137_596 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_164_382 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_125_747 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_164_393 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_125_769 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_51_Right_51 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_50_520 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_62_380 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_120_49 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_2_617 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_112_419 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7478__A1 net194 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_23_767 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_93_1628 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_136_Right_136 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_239_626 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_22_288 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_50_597 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_169_2544 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_38_34 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4161__C2 _0779_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_182_2700 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_207_512 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_38_67 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_207_523 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_234_353 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5256__A3 _1515_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7650__A1 _1279_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_60_Right_60 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__4464__A1 _1055_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_179_419 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_187_430 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_77_417 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7402__A1 net212 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_159_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_187_441 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6820_ core_0.execute.rf.reg_outputs\[2\]\[1\] _3087_ _3083_ _3089_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_159_132 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_225_90 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_187_474 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_230_592 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_202_283 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_34_924 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7197__B _3384_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3963_ core_0.execute.rf.reg_outputs\[7\]\[11\] _0530_ _0595_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_58_664 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6751_ _3041_ _3049_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XTAP_TAPCELL_ROW_102_1735 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_58_675 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_147_349 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_18_517 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5702_ _2096_ _2099_ _2102_ _2103_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_6682_ _2972_ _2999_ _3009_ _0243_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_156_861 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3894_ _0529_ _0530_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_57_185 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_70_76 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5177__C1 _1606_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_5_400 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_45_369 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5716__A1 _1124_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_14_681 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_5633_ _2025_ _2029_ _2033_ _2034_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_0_61_818 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4519__A2 _1106_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3990__A3 _0527_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_5_422 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_143_533 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_171_842 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_155_393 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_116_769 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_723 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5564_ _1963_ _1978_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_115_279 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_5_488 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7303_ _3473_ _3474_ _3478_ _0395_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__5445__B _1838_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4515_ _1101_ _1104_ _1105_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_8283_ _0459_ clknet_leaf_27_i_clk core_0.execute.pc_high_buff_out\[4\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_13_244 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5495_ _1925_ _1927_ _1928_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_41_586 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_103_Right_103 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_110_71 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_123_290 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_288 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7234_ _3409_ _3418_ _3419_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6141__A1 _2346_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4446_ _1040_ core_0.decode.i_instr_l\[2\] _1041_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_0_229_136 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_111_485 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_113_1864 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6692__A2 _3000_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7165_ _1369_ _1227_ _1230_ _3365_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_2
X_4377_ _0837_ _0947_ _0970_ _0990_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XANTENNA_clkbuf_leaf_30_i_clk_I clknet_4_10__leaf_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_226_821 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_224_3206 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6116_ _1457_ _2503_ _2504_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_186_97 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7096_ core_0.execute.alu_mul_div.mul_res\[11\] _3300_ _3305_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_226_865 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4575__I _1152_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_241_813 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7641__A1 _3732_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_213_504 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6047_ _1433_ _2436_ _0798_ _2437_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XANTENNA__5247__A3 _1553_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6444__A2 _2332_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_119_91 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_198_717 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4455__A1 _1037_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_198_728 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_142_2216 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_206_2983 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_68_1332 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_240_356 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_197_249 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_96_737 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4207__A1 _0824_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7819__C _1283_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7998_ _0175_ clknet_leaf_9_i_clk net137 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_95_247 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_178_485 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_193_422 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6949_ _1756_ _1754_ _1789_ _1752_ _1915_ _1364_ _3170_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux4_4
XPHY_EDGE_ROW_238_Right_238 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_154_809 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_193_455 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_166_669 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_235_3335 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_48_174 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_772 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_63_122 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_645 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_193_488 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_165_179 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_52_807 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_63_133 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_667 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5707__A1 _1123_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_63_155 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_146_382 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3981__A3 _0536_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_91_486 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_106_235 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_122_706 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_153_2345 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_32_520 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5183__A2 _1446_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_161_352 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6380__A1 _2244_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_32_531 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_79_1461 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_20_704 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6030__I _1456_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_737 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4143__B1 _0549_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_208_309 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6683__A2 _3006_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_5_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_236_629 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_246_3464 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_246_3475 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_216_331 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6186__B core_0.dec_mem_access vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7632__A1 core_0.execute.pc_high_buff_out\[3\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_216_353 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6435__A2 _1480_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5238__A3 _1451_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_232_813 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_188_205 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_164_2485 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_189_739 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_99_542 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_99_553 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6199__A1 _1379_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_231_389 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_86_236 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_86_247 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_169_474 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_130 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_169_496 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4749__A2 _1238_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5946__A1 core_0.execute.pc_high_buff_out\[1\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_69 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_74_409 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_200_765 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5946__B2 net8 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_205_Right_205 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_27_303 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_55_634 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_41_1004 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_28_859 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_55_645 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_144_308 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_94_291 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_144 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_55_667 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_70_604 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_153_842 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_11_640 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7163__A3 _3358_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_54_177 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_339 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_70_648 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_23_520 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_70_659 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_23_531 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_112_216 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xoutput206 net206 sr_bus_data_o[6] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
X_4300_ _0912_ _0915_ _0916_ _0917_ _0918_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_50_372 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6123__A1 _1137_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5280_ _1432_ core_0.execute.alu_mul_div.div_cur\[0\] _1726_ _1728_ _1729_ vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_0_121_772 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_66 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_10_247 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4231_ core_0.fetch.out_buffer_valid _0849_ _0850_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6674__A2 _3000_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_227_629 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_52_1133 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_207_320 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4162_ core_0.dec_l_reg_sel\[2\] _0781_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_156_34 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_235_651 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4395__I net84 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7623__A1 net201 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_65_43 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4093_ _0568_ core_0.execute.rf.reg_outputs\[4\]\[0\] _0520_ _0714_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_234_161 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4437__A1 _0812_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_234_172 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_234_183 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7921_ _0012_ clknet_leaf_121_i_clk core_0.decode.oc_alu_mode\[9\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_2
XANTENNA__4988__A2 _0773_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6824__B _3083_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_78_715 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_19_740 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_7852_ _0045_ clknet_leaf_67_i_clk core_0.fetch.out_buffer_data_instr\[29\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_81_31 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_77_236 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_148_625 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_175_400 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6803_ _2986_ _3065_ _3078_ _0295_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_187_282 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5937__A1 _2281_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8160__CLK clknet_leaf_88_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_172_88 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7783_ core_0.dec_rf_ie\[5\] _1133_ _3827_ _3845_ _3853_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_148_647 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_58_461 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4995_ _0770_ _0767_ _1444_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or2_4
XFILLER_0_46_612 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_314 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_58_483 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_147_146 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6734_ _2992_ _3022_ _3038_ _0266_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_163_606 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4070__C1 _0692_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3946_ _0570_ _0575_ _0579_ _0580_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_4
XTAP_TAPCELL_ROW_63_1273 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_46_667 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_34_807 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_116_511 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_6_731 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6665_ _2998_ _2999_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
X_5616_ _1513_ _1514_ _2017_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_116_566 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_143_352 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5165__A2 _1604_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_5_252 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6362__A1 _1059_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6596_ _2929_ _2943_ _2944_ _2945_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_0_83_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_60_158 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_103_216 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_143_385 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_171_694 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8335_ _0511_ clknet_leaf_9_i_clk core_0.dec_alu_flags_ie vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_230_3276 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4912__A2 _1221_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5547_ net85 _1953_ _1969_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_131_558 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_597 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6114__A1 _2010_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5478_ _1909_ _1592_ _1910_ _1911_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_8266_ _0442_ clknet_leaf_21_i_clk core_0.execute.sreg_irq_flags.o_d\[0\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_input55_I i_req_data[25] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_197_96 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7390__B _3553_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4429_ _0736_ net109 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_7217_ _1736_ _3396_ _3403_ _3404_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_111_282 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_3_7_0_i_clk_I clknet_0_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_8197_ _0373_ clknet_leaf_129_i_clk core_0.execute.alu_mul_div.div_res\[6\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__4676__A1 _1223_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_217_128 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5873__B1 _2265_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7148_ _3353_ _3354_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_226_651 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7614__A1 core_0.dec_sreg_jal_over vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7079_ _3286_ _3288_ _3290_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_225_172 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_214_835 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_213_312 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_241_632 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_213_334 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_213_345 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4979__A2 _1393_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_715 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_213_367 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6226__S _2356_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_241_698 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_179_772 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_68_247 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_138_102 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_194_731 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5928__A1 _1819_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_96_578 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_49_461 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_178_293 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_194_753 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_83_228 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_194_786 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_500 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_153_105 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_37_667 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_119_371 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_64_453 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_92_762 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_689 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_135_842 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_36_177 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_24_317 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5156__A2 core_0.dec_l_reg_sel\[1\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_51_136 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_134_374 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_150_834 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_161_182 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_161_193 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_681 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_110_709 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6105__A1 _1378_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_103_772 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6909__B _3139_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_209_618 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6656__A2 _2962_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6695__I _1963_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_166_2503 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_208_117 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_236_448 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4419__A1 _0883_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7081__A2 _3178_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_126_37 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6644__B _2984_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_231_142 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_189_558 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_99_372 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5631__A3 _2018_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_87_556 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_16_710 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5919__A1 _2300_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_157_422 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_169_282 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_200_540 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_28_601 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_177_2632 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_185_764 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4780_ _1290_ _1294_ _0056_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_200_584 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5395__A2 _1814_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_28_656 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_807 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_28_667 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_28_689 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6344__A1 core_0.ew_data\[10\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6450_ net76 _2531_ _2829_ _2537_ _2830_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__5707__C _2092_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_125_352 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_70_467 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5401_ core_0.execute.alu_mul_div.div_cur\[5\] _1715_ _1844_ _1845_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_30_309 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6895__A2 _3130_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6381_ _2242_ _0604_ _2762_ _2763_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_180_491 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_70_489 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_3_756 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_113_569 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8120_ _0296_ clknet_leaf_103_i_clk core_0.execute.rf.reg_outputs\[3\]\[11\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5332_ _1762_ _1777_ _1778_ _1779_ _1780_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai31_2
XFILLER_0_11_545 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8051_ _0227_ clknet_leaf_115_i_clk core_0.execute.rf.reg_outputs\[7\]\[6\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_2
XANTENNA__6647__A2 _2962_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5263_ _1523_ _1524_ _1712_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_TAPCELL_ROW_208_3009 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_188_2772 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_4214_ _0724_ net53 _0832_ _0833_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_4
X_7002_ _3214_ _3218_ _3175_ _3219_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_110_1834 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_5194_ _1481_ _1451_ _1643_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_2
XTAP_TAPCELL_ROW_126_2019 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_4145_ core_0.dec_used_operands\[1\] _0764_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_223_610 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_223_632 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_207_183 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4076_ _0690_ _0578_ _0693_ _0698_ _0699_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_0_223_665 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5083__A1 _1482_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_78_501 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_223_687 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_195_506 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7904_ _0095_ clknet_leaf_69_i_clk core_0.decode.i_imm_pass\[13\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_211_838 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_203_2953 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_210_326 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4830__A1 _1280_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_188_591 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7835_ _0028_ clknet_leaf_73_i_clk core_0.fetch.out_buffer_data_instr\[12\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_176_731 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_219_3138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_65_217 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_191_712 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5386__A2 _1831_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_121_1963 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_7766_ _3839_ _3840_ _3841_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__4189__A3 _0807_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6583__A1 _0785_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_163_414 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4978_ _1381_ _0553_ _1428_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_19_667 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6717_ _2967_ _3021_ _3029_ _0258_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_3929_ _0563_ net199 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_117_842 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_191_767 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_784 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7697_ _1038_ _1101_ _1041_ _3797_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_0_190_244 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_34_626 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_177 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_73_272 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_137_2159 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_22_779 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_18_199 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5138__A2 core_0.execute.rf.reg_outputs\[4\]\[8\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_61_434 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6648_ _2941_ _2986_ _2987_ _0231_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_144_672 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_150_2315 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6886__A2 _3106_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_143_182 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6579_ _2242_ _2202_ _2931_ _0218_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_61_489 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_76_1420 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8056__CLK clknet_leaf_104_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_14_383 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8318_ _0494_ clknet_leaf_11_i_clk core_0.dec_jump_cond_code\[3\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_30_865 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6729__B _3031_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output161_I net161 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6638__A2 core_0.ew_mem_width vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_8249_ _0425_ clknet_leaf_23_i_clk net105 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_4
XTAP_TAPCELL_ROW_243_3423 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_243_3434 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_148_2288 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_198_311 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7063__A2 _1592_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_214_654 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_161_2444 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_213_142 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5074__A1 _1467_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_241_462 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4763__I _0879_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_97_832 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_87_1560 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4821__A1 _0938_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_139_400 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_139_422 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6949__I0 _1756_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_56_206 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_139_444 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_127_606 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_166_252 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_154_403 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_182_712 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_139_488 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_194_594 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_65_762 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_182_745 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_52_401 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_330 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_24_103 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_423 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_92_592 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6326__A1 _2294_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5129__A2 _1568_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_123_812 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_172_2573 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6877__A2 _3114_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_150_631 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_122_333 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_122_344 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_110_517 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_237_702 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_110_539 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_209_404 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6629__A2 _2962_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4938__I _1381_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_209_426 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_20_375 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_209_437 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_237_768 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5301__A2 _1711_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_224_407 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_46_34 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_77_i_clk_I clknet_4_13__leaf_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_46_45 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_205_632 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_205_687 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6801__A2 _3064_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5950_ _1378_ core_0.execute.sreg_irq_pc.o_d\[1\] _2341_ _2342_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_0_88_865 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_87_342 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_158_720 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_177_539 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4901_ _1366_ _1367_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_153_57 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_220_679 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_48_729 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_141_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5881_ _1729_ _2244_ _2272_ _2273_ _2274_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_0_239_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7620_ core_0.execute.pc_high_buff_out\[0\] _3732_ _1216_ _3736_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_185_550 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_47_1076 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_4832_ core_0.decode.i_instr_l\[12\] _1321_ _1325_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_75_559 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7551_ _3674_ _3675_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XTAP_TAPCELL_ROW_60_1232 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_90_518 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4763_ _0879_ _1285_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_7_347 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_173_756 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4040__A2 _0523_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_172_244 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_15_103 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_272 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_172_255 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6502_ _1689_ _2130_ _2879_ _2123_ _2880_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_4
X_4694_ _1244_ _0020_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_70_220 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7482_ _3630_ _3628_ _3631_ _1950_ _0421_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_70_242 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_71_765 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_214_3079 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6868__A2 _3107_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6433_ _2090_ _2501_ _2626_ _2813_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_43_489 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4879__A1 _0886_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5009__I core_0.decode.oc_alu_mode\[11\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_113_366 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6364_ _1107_ _2736_ _2738_ _1121_ _2745_ _2746_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_0_140_163 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_3_586 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5540__A2 _1957_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_12_865 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8103_ _0279_ clknet_leaf_94_i_clk core_0.execute.rf.reg_outputs\[4\]\[10\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5453__B _1841_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5315_ core_0.execute.alu_mul_div.div_cur\[4\] _1695_ _1763_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__xor2_2
X_6295_ _2035_ _1455_ _2678_ _1754_ _2638_ _2679_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai221_2
X_8034_ _0211_ clknet_leaf_80_i_clk core_0.ew_reg_ie\[1\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_227_245 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5246_ _1461_ net204 _1694_ _1695_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_0_243_716 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_71_1361 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_89_Right_89 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_227_267 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5177_ core_0.execute.rf.reg_outputs\[5\]\[5\] _1604_ _1605_ core_0.execute.rf.reg_outputs\[7\]\[5\]
+ _1606_ core_0.execute.rf.reg_outputs\[3\]\[5\] _1626_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_0_236_790 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_208_481 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4128_ core_0.execute.prev_pc_high\[7\] _0742_ net112 _0744_ _0746_ _0747_ vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XANTENNA__5056__A1 _1466_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input18_I i_irq vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_196_804 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_127_80 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4059_ _0681_ _0594_ _0682_ _0683_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_97_139 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_210_101 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_27_838 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4803__A1 _1038_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_210_134 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_39_707 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_195_336 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6005__B1 _2265_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_195_369 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_183_509 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7818_ _3873_ _3875_ _3876_ _3877_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_0_148_263 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_93_345 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_98_Right_98 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_47_762 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_53_209 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_108_127 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3909__A3 _0544_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7749_ core_0.decode.i_instr_l\[9\] _1032_ _3827_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_0_46_261 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_191_553 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_124_609 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_62_732 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_661 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_191_586 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_151_417 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_445 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6859__A2 _3108_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_61_264 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_116_193 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_120_804 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_21_139 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_131_152 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5531__A2 _1956_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output86_I net86 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_219_702 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4590__I0 core_0.ew_data\[1\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_30_662 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_18_Left_265 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__7808__A1 _0789_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_218_212 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_218_234 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4098__A2 _0521_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_206_407 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_233_204 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_218_289 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_7_596 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_199_642 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_28 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_37 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_202_613 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_198_163 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6795__A1 _2972_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_186_314 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_69_342 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_198_196 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_27_Left_274 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__4270__A2 _0823_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_526 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_323 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_201_189 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_174_2602 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_167_594 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_154_233 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_154_244 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_142_417 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_317 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5770__A2 _1568_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_170_737 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_96_1659 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_52_297 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_36_Left_283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_40_459 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_123_686 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5522__A2 core_0.decode.o_submit vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_0_512 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6570__I1 core_0.ew_reg_ie\[5\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_150_483 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_209_212 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_185_2731 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_5100_ _1543_ _1548_ _1549_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_4
XANTENNA__7275__A2 net87 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6080_ _1603_ _1623_ _1640_ _1600_ _2469_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA_clkbuf_4_9__f_i_clk_I clknet_3_4_0_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_66 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5286__A1 _0810_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_209_278 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_189_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5031_ _1479_ _1480_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XANTENNA__6883__I _0722_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7027__A2 _1939_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_164_34 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_49_1105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_79_128 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_178_804 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_45_Left_292 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
X_6982_ _1908_ _1931_ _3200_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__6786__A1 core_0.execute.rf.reg_outputs\[3\]\[3\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_232_281 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_189_174 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_73_76 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_232_292 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_88_651 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_200_2912 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_220_454 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5933_ _1603_ _2321_ _2324_ _1624_ _2325_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_177_347 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_177_358 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4261__A2 _0879_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_105_1777 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_196_2860 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_48_559 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5864_ _2256_ _2257_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XTAP_TAPCELL_ROW_216_3108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_158_594 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7603_ core_0.execute.pc_high_out\[6\] _3673_ _3720_ _3721_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4815_ _0865_ core_0.decode.i_instr_l\[6\] _1305_ _1314_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_75_378 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_63_529 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4013__A2 _0594_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5210__A1 _0771_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5795_ _2187_ _2194_ _2195_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_8_667 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_133_406 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_743 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_28_294 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7534_ _3581_ _3662_ _0442_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_4746_ net57 _1241_ _1274_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_44_754 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_32_896 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_134_2118 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_43_242 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_467 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_562 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7465_ _3563_ net77 _3540_ _3617_ _3618_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_4677_ _1232_ _1233_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_102_804 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_43_297 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_114_664 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6416_ _2576_ _2795_ _2796_ _0190_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_114_675 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6710__A1 _2951_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_101_303 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7396_ net221 _3544_ _3560_ _3561_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_141_483 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_12_662 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6347_ _2119_ _2117_ _1625_ _2729_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_12_673 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_101_347 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_100_i_clk_I clknet_4_7__leaf_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_227_3237 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_11_183 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6278_ _1379_ core_0.execute.sreg_irq_pc.o_d\[9\] _2662_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_215_204 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8017_ _0194_ clknet_leaf_48_i_clk core_0.ew_addr\[0\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5229_ _1625_ _1665_ _1677_ _1559_ _1678_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_0_138_90 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_243_557 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_4_555 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_145_2247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_243_568 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_215_259 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_4_566 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_145_2258 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6077__I0 _2013_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5029__A1 _1467_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_169_815 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_98_448 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6777__A1 core_0.ew_reg_ie\[3\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_168_314 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_223_292 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_224_37 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_196_645 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6241__A3 _1452_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_85_109 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_196_656 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_196_667 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6742__B _3031_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_184_807 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4252__A2 _0870_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_695 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_559 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_183_317 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6529__A1 net116 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_238_3366 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_93_142 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_26_209 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_clkbuf_leaf_25_i_clk_I clknet_4_10__leaf_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4004__A2 _0541_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5201__A1 core_0.execute.rf.reg_outputs\[2\]\[1\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_117_Right_117 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_35_721 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_136_244 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5201__B2 _0769_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_164_575 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_34_231 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5752__A2 _1631_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_164_597 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_156_2387 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4689__S _1241_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_264 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_713 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_105_642 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_22_426 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_132_450 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_120_601 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_163 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_697 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6701__A1 _2996_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_219_554 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6917__B _3139_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_206_215 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_118_27 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7009__A2 _3184_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_89_415 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_89_426 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_180_2672 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_202_421 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_187_623 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6768__A1 _2988_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_230_741 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_202_432 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4779__B1 _0881_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_186_122 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_76_109 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_134_37 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_202_454 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_175_807 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_85_621 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_187_678 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_409 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_97_492 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_186_177 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_174_317 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_44_1035 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_44_1046 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7193__A1 _2891_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_127_244 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4600_ core_0.ew_data\[6\] core_0.ew_data\[14\] _1150_ _1165_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_38_592 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_732 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_127_266 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6940__A1 _1227_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5580_ core_0.dec_sys _0177_ _1983_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_150_69 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_182_383 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_143_748 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_702 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_562 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_142_236 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7483__B _3384_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_53_573 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4531_ _1117_ _1053_ _1118_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_41_724 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_142_247 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_41_735 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_80_370 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_104_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_211_3049 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_13_437 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_7250_ _3429_ _3432_ _1395_ _0388_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_40_234 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4462_ _1038_ _1043_ _1056_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_0_110_100 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_159_34 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_111_634 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6201_ core_0.execute.alu_mul_div.mul_res\[7\] _2587_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_2
X_4393_ net85 _0883_ _1003_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_7181_ _1748_ _3375_ _0376_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_111_656 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_0_342 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_21_492 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_111_689 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6132_ _2505_ _2510_ _2514_ _2519_ _2520_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_0_110_166 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_238_863 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_110_177 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_55_1175 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6827__B _3083_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5259__A1 _1701_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5731__B _2113_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6063_ net82 _2268_ _2451_ _2245_ _2452_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XPHY_EDGE_ROW_53_Left_300 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
X_5014_ _0568_ core_0.execute.rf.reg_outputs\[3\]\[0\] _0549_ _1463_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__and3_1
XPHY_EDGE_ROW_219_Right_219 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_175_99 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_240_527 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4482__A2 _1072_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_1_525 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_222_3178 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_240_549 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_221_730 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6759__A1 _2977_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_37_955 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_191_54 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6965_ _3183_ _3184_ _1366_ _1229_ _3185_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai211_4
XFILLER_0_48_301 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_166_807 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5431__A1 core_0.execute.alu_mul_div.div_cur\[8\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_178_667 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_166_829 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5916_ _1819_ _1585_ _2307_ _1624_ _2308_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai211_2
XTAP_TAPCELL_ROW_140_2188 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6054__S _2190_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_192_103 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_177_177 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_131 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6896_ _2946_ _3129_ _3132_ _0334_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_119_734 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_165_339 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_8_420 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3993__A1 _0517_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_48_378 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_75_164 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_76_687 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_146_531 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_17_710 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7184__A1 _1362_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5847_ _2202_ _2239_ _2240_ _0176_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_63_326 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_29_581 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_118_255 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_337 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5778_ _1713_ net214 _2179_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_134_737 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_173_394 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7517_ core_0.execute.sreg_scratch.o_d\[8\] _3646_ _3651_ _3654_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_118_1924 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_4729_ _0858_ _1238_ _1265_ _0034_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__4810__B _1311_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_31_212 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_114_450 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_102_601 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7448_ _0604_ _3546_ _3545_ _3603_ _3604_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__6534__I1 _2440_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7731__I0 net179 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_31_256 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_9_625 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_102_645 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_102_667 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7379_ _3540_ _3546_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XANTENNA__4101__I net71 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_101_177 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6737__B _3031_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6447__B1 _2534_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_101_199 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_228_373 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_216_513 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_max_cap218_I _1484_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_203_207 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4473__A2 _1039_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_231_527 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_99_746 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_235_69 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_224_590 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7411__A2 _1008_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_196_453 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6472__B _2849_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5422__A1 _1375_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_67_632 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_158_2405 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_104_18 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_168_177 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_clkbuf_4_15__f_i_clk_I clknet_3_7_0_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_94_440 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_137_520 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_184_659 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3984__A1 _0608_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5088__B _0779_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_94_473 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7175__A1 _3357_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_183_158 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_657 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_152_501 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5186__B1 _1437_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_109_277 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5725__A2 _2092_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_125_737 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6922__A1 _2992_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_35_562 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_702 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_125_759 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_124_247 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_180_865 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_22_234 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7478__A2 _1398_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_256 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_93_1629 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_50_576 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5489__A1 _1367_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_120_420 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_238_104 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_169_2545 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4161__A1 core_0.ew_reg_ie\[3\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4161__B2 core_0.ew_reg_ie\[2\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6647__B _2984_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_120_497 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5551__B _1964_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_182_2701 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_219_384 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_38_79 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7650__A2 _1945_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_89_212 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_234_387 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_222_527 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5661__A1 _2045_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_54_78 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_54_89 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7402__A2 _3544_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_148_807 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_225_80 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5413__A1 core_0.execute.alu_mul_div.div_cur\[7\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_34_925 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6750_ _2956_ _3042_ _3048_ _0272_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_174_103 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_202_295 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3962_ _0516_ _0540_ _0518_ _0594_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_4
XFILLER_0_58_654 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5964__A2 _2342_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_102_1736 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_5701_ _2101_ _2102_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_221_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_193_2830 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6681_ core_0.execute.rf.reg_outputs\[6\]\[6\] _3006_ _3004_ _3009_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__7166__A1 _3358_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3893_ core_0.dec_r_reg_sel\[2\] core_0.dec_r_reg_sel\[1\] _0518_ _0529_ vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and3_2
XFILLER_0_190_629 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_72_123 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5177__B1 _1605_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5632_ _2030_ _2031_ _2032_ _2033_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XANTENNA__5716__A2 _1568_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_14_682 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6913__A1 net103 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_115_214 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_128_597 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3990__A4 core_0.execute.rf.reg_outputs\[6\]\[9\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_170_331 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_584 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5563_ net78 _1977_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_53_370 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_13_212 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_170_364 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7302_ _3384_ _3477_ _3478_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4514_ _1055_ _1103_ _1104_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_8282_ _0458_ clknet_leaf_29_i_clk core_0.execute.pc_high_buff_out\[3\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_41_554 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_79_64 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5494_ _1451_ _1926_ _1927_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_110_61 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7233_ _2453_ _3417_ _3418_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_13_278 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_640 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_110_83 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4445_ core_0.decode.i_instr_l\[3\] _1040_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__inv_3
XANTENNA__6141__A2 net227 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7164_ _3363_ _3364_ _3357_ _0370_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_113_1865 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_4376_ _0892_ _0952_ _0988_ _0989_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_0_172 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_238_671 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5461__B _1816_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6115_ _2152_ _2463_ _2010_ _2503_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__4856__I _1305_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_95_74 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7095_ _3304_ _0361_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_95_85 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_95_96 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_119_81 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6046_ core_0.execute.alu_mul_div.mul_res\[3\] _2436_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XANTENNA__5247__A4 _1641_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_28_90 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_213_516 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_60_i_clk clknet_4_14__leaf_i_clk clknet_leaf_60_i_clk vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_TAPCELL_ROW_142_2217 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_197_206 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_241_858 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_206_2984 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_68_1333 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_95_204 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_178_442 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5404__A1 core_0.execute.alu_mul_div.div_cur\[4\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
X_7997_ _0174_ clknet_leaf_120_i_clk net136 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_221_571 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_49_632 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_138_306 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_138_317 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6948_ _1225_ _3167_ _3168_ _3169_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_0_138_328 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_165_114 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_193_434 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_75_i_clk clknet_4_13__leaf_i_clk clknet_leaf_75_i_clk vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__3966__A1 _0565_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_235_3336 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7157__A1 _2331_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6879_ core_0.execute.rf.reg_outputs\[1\]\[11\] _3114_ _3112_ _3122_ vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_63_101 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_91_410 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_165_158 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5168__B1 _1437_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_64_657 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5707__A2 _1652_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_17_540 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6904__A1 net99 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_107_748 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_562 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_167 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output191_I net191 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_106_247 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_153_2346 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_162_865 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_44_370 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_258 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4540__B _1101_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_134_567 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6380__A2 _2752_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_122_729 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_79_1462 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_121_206 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_60_863 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_13_i_clk clknet_4_9__leaf_i_clk clknet_leaf_13_i_clk vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__4143__A1 core_0.ew_reg_ie\[2\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4143__B2 core_0.ew_reg_ie\[3\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_102_497 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_246_3465 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_246_3476 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7632__A2 _3731_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_28_i_clk clknet_4_10__leaf_i_clk clknet_leaf_28_i_clk vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__4446__A2 core_0.decode.i_instr_l\[2\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_164_2475 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_216_387 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_204_527 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_164_2486 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_231_368 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_59_418 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_99_598 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6199__A2 core_0.execute.sreg_irq_pc.o_d\[7\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7396__A1 net221 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_37 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_200_733 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_197_784 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_169_486 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5946__A2 _2249_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_184_423 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_39_142 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_129_339 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_157_648 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_55_613 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_41_1005 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_55_657 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_137_361 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_184_489 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_43_808 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_125_534 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_125_545 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_69 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_11_641 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_180_651 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_54_189 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_113_718 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4382__A1 _0959_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_23_543 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_437 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput207 net207 sr_bus_data_o[7] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_23_576 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_140_548 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_239_413 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7761__B _1116_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_34 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6123__A2 _1693_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_10_226 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4230_ core_0.fetch.out_buffer_data_instr\[16\] _0849_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__4685__A2 _1237_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4161_ core_0.ew_reg_ie\[3\] _0774_ _0777_ core_0.ew_reg_ie\[2\] core_0.ew_reg_ie\[1\]
+ _0779_ _0780_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XTAP_TAPCELL_ROW_52_1134 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_4092_ _0710_ _0594_ _0711_ _0712_ _0713_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai211_4
XFILLER_0_223_814 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_128_2050 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_171_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_235_696 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_223_847 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7920_ _0011_ clknet_leaf_8_i_clk core_0.execute.alu_mul_div.i_mul vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_4
XANTENNA__5501__S _1492_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4988__A3 _0769_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_236_90 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_77_204 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7851_ _0044_ clknet_leaf_66_i_clk core_0.fetch.out_buffer_data_instr\[28\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_19_741 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_222_379 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_172_34 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6802_ core_0.execute.rf.reg_outputs\[3\]\[10\] _3070_ _3072_ _3078_ vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_81_65 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5300__I _1747_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7782_ _1136_ _3852_ _0500_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__5937__A2 core_0.execute.alu_mul_div.mul_res\[1\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
X_4994_ _0770_ _0783_ _1443_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_6733_ core_0.execute.rf.reg_outputs\[5\]\[13\] _3027_ _3031_ _3038_ vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_175_456 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7139__A1 _1915_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3945_ _0576_ _0578_ _0579_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__4070__B1 _0662_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6840__B _3098_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_63_1263 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4070__C2 core_0.execute.rf.reg_outputs\[1\]\[2\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_18_348 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_63_1274 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_45_134 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_18_359 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6664_ core_0.ew_reg_ie\[6\] _2934_ _2998_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_0_128_372 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_190_437 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_162_139 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5615_ _2012_ _2015_ _2016_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_60_104 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_144_865 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_171_640 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6595_ net28 _1150_ _2944_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_26_370 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_521 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_26_392 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_104_729 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4373__A1 _0982_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_8334_ _0510_ clknet_leaf_9_i_clk core_0.dec_alu_carry_en vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_42_863 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5546_ core_0.execute.mem_stage_pc\[7\] _1968_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_103_228 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_230_3277 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_76_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8265_ _0441_ clknet_leaf_33_i_clk core_0.execute.sreg_scratch.o_d\[15\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__7311__A1 _3409_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5477_ _1908_ _1620_ _1910_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7216_ net80 _3398_ _3399_ _3402_ _3403_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_4428_ _0739_ net108 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_8196_ _0372_ clknet_leaf_2_i_clk core_0.execute.alu_mul_div.div_res\[5\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_1_492 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_input48_I i_req_data[19] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4676__A2 _1225_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5873__B2 core_0.execute.alu_flag_reg.o_d\[0\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7147_ _1719_ _3209_ _3189_ _3353_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4359_ _0946_ _0956_ _0974_ _0975_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_0_226_663 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_214_803 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7078_ _3286_ _3288_ _3289_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_226_685 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_213_302 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5625__A1 _1999_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6029_ _1480_ _2411_ _2418_ _2419_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_241_644 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_240_132 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_198_559 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_96_502 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_96_546 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA_output204_I net204 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5928__A2 _1637_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_451 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_77_760 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6050__A1 _2438_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_193_220 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_232_37 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_49_473 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3939__A1 _0568_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_37_624 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_484 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_166_467 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_64_421 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_166_478 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_194_798 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_36_123 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_154_629 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7565__C _1950_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_51_104 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_150_802 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7550__A1 _1209_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_17_381 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6353__A2 _2695_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_150_813 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4364__A1 core_0.fetch.prev_request_pc\[12\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_513 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7302__A1 _3384_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_32_384 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_32_395 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4116__A1 core_0.execute.pc_high_out\[1\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_103_784 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_130_581 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_166_2504 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_208_107 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4496__I core_0.execute.alu_mul_div.i_mul vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8328__CLK clknet_leaf_89_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5616__A1 _1513_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6925__B _3139_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_189_515 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_244_493 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_205_858 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_126_49 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_87_502 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_59_204 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_16_700 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_129_103 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_129_114 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_200_552 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_68_771 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_207 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_177_2633 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_28_613 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_129_136 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_142_37 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6592__A2 _2941_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_157_478 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_145_629 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_185_798 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_55_454 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_73_i_clk_I clknet_4_13__leaf_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_43_627 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_413 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_82_273 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_126_865 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6344__A2 _2486_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_3_702 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4355__A1 _0964_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_70_457 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5400_ _1763_ _1775_ _1776_ _1844_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_125_375 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_863 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_340 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_152_172 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6380_ _2244_ _2752_ _2761_ _2241_ _2762_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_11_502 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_768 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5331_ core_0.execute.alu_mul_div.div_cur\[6\] _1761_ _1779_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_23_384 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_239_243 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8050_ _0226_ clknet_leaf_115_i_clk core_0.execute.rf.reg_outputs\[7\]\[5\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_2
XANTENNA__5723__C _2092_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5262_ _1521_ _1522_ _1711_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_4
XFILLER_0_121_581 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_188_2773 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_7001_ _3212_ _3217_ _3218_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__5855__A1 net186 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4213_ _0724_ _0831_ _0832_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_110_1835 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_167_67 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5193_ _1603_ _1623_ _1640_ net223 _1642_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_0_76_98 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4144_ core_0.ew_reg_ie\[0\] _0520_ _0758_ core_0.ew_reg_ie\[1\] _0763_ vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_0_207_151 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_235_471 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6835__B _3083_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5607__A1 _1676_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_223_644 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4075_ _0694_ _0695_ _0696_ _0697_ _0698_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and4_1
XANTENNA__5083__A2 _1491_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7903_ _0094_ clknet_leaf_68_i_clk core_0.decode.i_imm_pass\[12\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_203_2943 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_223_699 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_78_535 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_222_187 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_203_2954 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_148_401 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4830__A2 net40 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_78_568 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7834_ _0027_ clknet_leaf_81_i_clk core_0.fetch.out_buffer_data_instr\[11\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_219_3139 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_19_624 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_101 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_65_229 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7765_ _1068_ _1075_ _3784_ _3840_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_121_1964 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_4977_ _1419_ _1427_ _0120_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__7780__A1 _1136_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6583__A2 _2190_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_136_629 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_176_798 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_191_735 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6716_ core_0.execute.rf.reg_outputs\[5\]\[5\] _3027_ _3016_ _3029_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3928_ net93 _0521_ _0557_ _0562_ _0563_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai22_4
X_7696_ _3794_ _3795_ _3796_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_34_638 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6647_ core_0.execute.rf.reg_outputs\[7\]\[10\] _2962_ _2984_ _2987_ vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_144_651 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7532__A1 _0553_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6335__A2 _1386_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_190_278 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_27_690 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_116_375 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4346__A1 _0883_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7995__CLK clknet_leaf_89_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_150_2316 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6578_ _2930_ _1985_ _2931_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_171_492 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_76_1421 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_8317_ _0493_ clknet_leaf_10_i_clk core_0.dec_jump_cond_code\[2\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_2
X_5529_ _1955_ _1957_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA__6099__A1 _2202_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_30_855 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8248_ _0424_ clknet_leaf_20_i_clk core_0.execute.trap_flag vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_100_732 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5846__A1 net138 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_245_224 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8179_ _0355_ clknet_leaf_127_i_clk core_0.execute.alu_mul_div.mul_res\[5\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_2
XTAP_TAPCELL_ROW_243_3424 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_10_590 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_233_419 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7599__A1 core_0.execute.pc_high_buff_out\[6\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6745__B _3045_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_148_2289 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_214_633 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_161_2445 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6271__A1 core_0.ew_data\[8\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_202_817 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5074__A2 net183 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4282__B1 _0886_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_87_1561 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_96_321 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_213_187 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_167_710 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4821__A2 _1170_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_213_198 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_139_412 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_579 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6023__A1 _1624_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6949__I1 _1754_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_167_754 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_84_527 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_96_387 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_167_765 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7771__A1 core_0.decode.i_instr_l\[8\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_194_584 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_181_201 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_181_212 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_64_240 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5782__B1 _2136_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_126_139 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_37_476 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_52_413 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5096__B _0779_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_181_245 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_182_779 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_24_115 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_80_733 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_865 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_135_673 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4337__A1 core_0.fetch.prev_request_pc\[12\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_52_457 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_190_790 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_172_2574 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_33_671 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_98_1690 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_0_716 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_103_570 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_20_387 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_205_622 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_204_132 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_232_452 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6262__A1 _2281_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4273__B1 _0844_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_88_855 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4812__A2 _1306_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_220_647 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_204_198 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4900_ core_0.execute.alu_mul_div.cbit\[2\] _1366_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__inv_3
XFILLER_0_62_34 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_158_732 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5880_ core_0.dec_sreg_jal_over _2270_ _2273_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_201_850 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6014__A1 _1380_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_62_89 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4831_ _1322_ _1324_ _0077_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_185_562 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_47_1077 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_173_702 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_134_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_28_443 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_173_724 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4576__A1 core_0.ew_data\[2\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7550_ _1209_ _2257_ _3674_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__5718__C _2092_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4762_ _1283_ _1284_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XTAP_TAPCELL_ROW_60_1233 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_117_139 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_145_459 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_172_234 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6501_ _1689_ _2126_ _2127_ _2879_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_0_16_649 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7481_ core_0.execute.sreg_jtr_buff.o_d\[1\] _1398_ _3628_ _3631_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__7514__A1 net215 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4693_ core_0.fetch.out_buffer_data_instr\[4\] net64 _1241_ _1244_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_6432_ _2810_ _2811_ _2133_ _2812_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_114_857 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_141_632 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_153_492 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_107 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_102_95 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4879__A2 _1321_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6363_ _2411_ _2642_ _2744_ _2745_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_101_507 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_855 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8102_ _0278_ clknet_leaf_107_i_clk core_0.execute.rf.reg_outputs\[4\]\[9\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_113_389 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5314_ core_0.execute.alu_mul_div.div_cur\[6\] _1761_ _1762_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__7817__A2 _3806_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6294_ core_0.decode.oc_alu_mode\[2\] _1585_ core_0.decode.oc_alu_mode\[7\] _2678_
+ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_227_202 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5828__A1 _2202_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_8033_ _0210_ clknet_leaf_86_i_clk core_0.ew_reg_ie\[0\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5245_ _1466_ net188 _1694_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_TAPCELL_ROW_71_1362 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4500__A1 _0514_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_227_279 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_215_419 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5176_ _1482_ _1625_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_199_109 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_242_249 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4127_ core_0.execute.prev_pc_high\[7\] _0742_ _0745_ core_0.execute.prev_pc_high\[6\]
+ _0746_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_0_235_290 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5056__A2 net193 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4058_ _0533_ _0541_ _0543_ core_0.execute.rf.reg_outputs\[5\]\[3\] _0682_ vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_0_78_332 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_27_839 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4803__A2 _1307_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_195_326 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_94_803 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_4_10__f_i_clk clknet_3_5_0_i_clk clknet_4_10__leaf_i_clk vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_195_348 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_516 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6005__A1 core_0.execute.pc_high_buff_out\[3\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_66_527 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6005__B2 core_0.execute.alu_flag_reg.o_d\[3\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7817_ _1077_ _3806_ _3876_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__7753__A1 core_0.decode.i_instr_l\[10\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_149_787 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_629 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8023__CLK clknet_leaf_36_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4567__A1 core_0.ew_addr\[0\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7748_ _3825_ _3826_ _0492_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_163_212 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_82_1491 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_191_543 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_117_640 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_435 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7679_ _1082_ _1090_ _1078_ _3779_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_117_673 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_163_278 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4104__I _0723_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_117_695 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_777 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_104_312 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_116_172 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_131_142 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7808__A2 _1134_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4590__I1 core_0.ew_data\[9\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_219_725 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_246_522 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output79_I net79 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5819__A1 net134 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_218_224 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_219_769 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_234_717 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6492__A1 core_0.ew_data\[14\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_21_i_clk_I clknet_4_8__leaf_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_7_597 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6475__B _2851_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_233_227 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_18 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_198_120 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_88_107 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5047__A2 net218 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_199_665 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6795__A2 _3064_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_241_282 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_332 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_186_326 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_201_146 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_97_674 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_84_302 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_97_685 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_84_313 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_398 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_858 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_155_702 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_167_562 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7744__A1 core_0.decode.i_instr_l\[7\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_32_37 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_174_2603 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_84_357 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4558__A1 _1041_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_37_273 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_203_72 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_25_435 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_114_109 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_123_632 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_135_492 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_40_405 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_287 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_122_131 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_123_698 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4730__A1 net48 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_122_197 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_546 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_20_162 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_131_2090 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_209_235 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_185_2732 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6483__A1 _2447_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5286__A2 _1734_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5030_ _1467_ net213 _1478_ _1479_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_4
XANTENNA__4494__B1 _1064_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6235__A1 net86 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5038__A2 _1486_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6235__B2 _2537_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_189_142 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_49_1106 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6981_ _1226_ _1676_ _3199_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_178_827 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6786__A2 _3065_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4797__A1 _1301_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5932_ _2322_ _2323_ net224 _2324_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_88_663 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_200_2913 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7035__I0 _3202_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_105_1767 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_105_1778 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_5863_ net186 _1198_ _2247_ _2256_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_0_180_34 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_75_335 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_118_404 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_196_2861 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_8_613 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_216_3109 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_7602_ net215 _3670_ _3672_ _3719_ _3720_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_29_752 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_118_426 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_145_212 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4814_ _1067_ core_0.fetch.submitable _1313_ _0071_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__4549__A1 _0812_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_7_123 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5794_ _1647_ _2192_ _2193_ _2194_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_0_44_722 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5210__A2 _0768_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8196__CLK clknet_leaf_2_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_113_72 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7533_ core_0.execute.irq_en net18 _1398_ core_0.execute.sreg_irq_flags.o_d\[0\]
+ _3662_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_4745_ _1273_ _0042_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_28_284 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_7_156 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_32_897 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_22_81 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_134_2119 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_160_226 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7464_ net37 _3616_ _3617_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4676_ _1223_ _1225_ _1231_ _1232_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_4
XFILLER_0_126_492 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_31_416 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_113_131 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6415_ core_0.ew_data\[12\] _2486_ _2796_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_189_76 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_31_438 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_4_863 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_113_142 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_98_85 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7395_ _1357_ _1959_ _3546_ _3559_ _3560_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__6710__A2 _3021_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5513__A3 _1172_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_3_384 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6346_ _2113_ _2603_ _2728_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_228_511 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_227_3238 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6277_ _1379_ _2660_ _2661_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_243_503 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8016_ _0193_ clknet_leaf_49_i_clk core_0.ew_data\[15\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_228_588 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5228_ _1625_ _1676_ _1677_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_input30_I i_mem_data[3] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4808__B _1310_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_145_2248 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_4_556 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_5159_ core_0.dec_l_reg_sel\[2\] core_0.dec_l_reg_sel\[1\] _1608_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_4
XANTENNA__5029__A2 net187 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_98_438 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_211_422 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6777__A2 _2934_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4788__A1 _1290_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_84_1520 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output117_I net117 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_67_814 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_137_702 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_67_858 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_149_562 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6529__A2 _1985_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_238_3367 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_109_404 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_426 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_164_521 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_93_154 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_82_839 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_94_699 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_109_448 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_192_863 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4004__A3 _0543_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5201__A2 _1438_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_137_768 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_240_37 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_124_407 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_744 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_221 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_755 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_191_384 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_62_541 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_156_2388 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_34_243 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_470 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7573__C _1950_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_105_632 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_117_492 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4960__B2 _1391_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50_725 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6701__A2 _3000_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6465__A1 _2090_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5268__A2 _1711_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_234_536 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_206_227 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_221_208 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_215_772 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_180_2673 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6768__A2 _3043_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_230_731 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_186_101 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_159_315 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4009__I _0637_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_214_293 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4779__A1 core_0.fetch.prev_request_pc\[7\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_159_337 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4779__B2 net174 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_159_348 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_97_471 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_230_786 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5549__B _1964_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_195 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_128_702 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_174_307 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7717__A1 core_0.decode.i_imm_pass\[3\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_186_189 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_84_143 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_44_1036 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_127_212 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__7906__CLK clknet_leaf_68_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_85_699 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_183_863 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_150_37 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_5_605 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_349 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4251__I0 net63 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_115_418 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_755 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6940__A2 _1715_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4530_ core_0.execute.alu_mul_div.i_mod _1117_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XANTENNA__4951__A1 _1301_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_230_70 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_40_202 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_4_148 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_53_585 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_211_3039 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_80_382 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_224 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_80_393 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4461_ core_0.decode.i_instr_l\[0\] _1039_ _1055_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_0_41_769 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6200_ _2542_ _2585_ _2586_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_7180_ _1926_ _3373_ core_0.execute.alu_mul_div.div_res\[9\] _3375_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_110_123 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4392_ _1001_ _0833_ _0959_ _1002_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_150_292 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6131_ _1831_ _2516_ _2518_ _2412_ _2519_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai211_4
XFILLER_0_110_156 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_0_376 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_237_352 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6456__A1 _2360_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_55_1176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5259__A2 _1702_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6062_ _2445_ _2446_ _2449_ _2450_ _2451_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_0_175_34 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4628__B core_0.execute.alu_flag_reg.o_d\[1\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_0_Left_247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
X_5013_ _1461_ _1382_ _1462_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_0_225_558 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_183_Right_183 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_240_506 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_240_517 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_212_219 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_1_526 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_108_72 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_222_3179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_206_794 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6759__A2 _3042_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_177_101 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_5_Right_5 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_37_956 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6964_ net217 _1650_ _1651_ core_0.execute.alu_mul_div.cbit\[0\] _3184_ vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XANTENNA__5431__A2 _1838_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5915_ _1554_ _1576_ _2307_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_49_858 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_88_493 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_140_2189 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4363__B _0945_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6895_ net95 _3130_ _3124_ _3132_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__7708__A1 _1039_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_146_521 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3993__A2 _0524_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5846_ net138 _2209_ _2240_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_119_746 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_839 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_91_614 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_124_93 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_91 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7184__A2 _3373_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_118_234 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5195__A1 _1558_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_146_576 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5777_ _2074_ _2080_ _2175_ _2177_ _2178_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai31_2
XFILLER_0_17_766 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_161_535 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7516_ net216 _3640_ _3653_ _0433_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_4728_ net47 _1253_ _1265_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_118_1925 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_90_179 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_140_70 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7447_ _3563_ net74 _3553_ _3602_ _3603_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_71_393 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4659_ _1216_ _1217_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_32_769 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_4_682 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_9_615 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5498__A2 _1483_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_9_626 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_31_279 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7378_ _3541_ _3545_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_229_831 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_229_842 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6329_ _1088_ core_0.execute.alu_mul_div.mul_res\[10\] _2712_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_228_341 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_244_801 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_244_823 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6447__B2 net5 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_110_690 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_90_1590 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_150_Right_150 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_169_602 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_243_399 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_169_613 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_99_769 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_196_421 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5958__B1 _2249_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7929__CLK clknet_leaf_24_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_67_611 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_157_808 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_184_605 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_212_797 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_644 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_158_2406 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_94_452 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_368 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3984__A2 _0613_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_67_699 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_109_245 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_137_576 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_192_671 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5186__B2 core_0.execute.rf.reg_outputs\[2\]\[4\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_164_362 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_82_669 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_205_Left_452 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__6922__A2 _3130_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_164_384 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_120_18 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_62_360 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_213 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_90_691 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_462 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_23_769 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6686__A1 _2981_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50_566 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6928__B _3149_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_120_454 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_169_2535 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_169_2546 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_219_352 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6438__A1 _1994_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_182_2702 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_235_834 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_234_311 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_214_Left_461 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_234_355 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_234_366 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4167__C _0785_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7759__B _1101_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_203_720 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_89_235 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_159_101 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_159_112 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_199_292 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_89_279 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_202_263 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5413__A2 _1811_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_225_92 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_34_915 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5279__B _1432_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_34_926 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_3961_ core_0.execute.rf.reg_outputs\[1\]\[11\] _0593_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_230_594 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_85_430 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_159_178 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5700_ _1596_ _2100_ _2101_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_85_452 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_102_1737 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6680_ _2967_ _2999_ _3008_ _0242_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__3975__A2 _0530_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_193_2831 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_46_839 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3892_ _0517_ _0524_ _0527_ _0528_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_4
XPHY_EDGE_ROW_223_Left_470 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_73_636 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_45_338 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5631_ _1761_ _2019_ _2018_ _2032_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_1
XANTENNA__5177__B2 core_0.execute.rf.reg_outputs\[7\]\[5\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_155_362 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_214_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4911__B _1223_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_155_373 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_14_683 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6913__A2 _3135_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_170_310 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_60_308 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5562_ _0964_ _1957_ _1976_ _0156_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__4924__A1 _1195_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_500 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_143_557 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7301_ net76 _3475_ _3476_ _1735_ _3477_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_5_468 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4513_ core_0.decode.i_instr_l\[3\] core_0.decode.i_instr_l\[2\] _1103_ vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_8281_ _0457_ clknet_leaf_29_i_clk core_0.execute.pc_high_buff_out\[2\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5493_ core_0.execute.alu_mul_div.cbit\[0\] _1228_ _1926_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_0_170_387 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7232_ _1430_ _1404_ _2482_ _3391_ _3417_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_111_432 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4444_ core_0.decode.i_instr_l\[1\] _1039_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_123_292 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6838__B _3098_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7163_ _1369_ _1362_ _3358_ _3364_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_4375_ _0892_ _0952_ _0946_ _0988_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_113_1866 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5234__S _1460_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6114_ _2010_ _2152_ _2463_ _2502_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_244_119 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_238_683 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_186_77 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7094_ core_0.execute.alu_mul_div.mul_res\[11\] _3303_ _3189_ _3304_ vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__5101__A1 _1531_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6045_ _2281_ _2434_ _2435_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_clkbuf_leaf_68_i_clk_I clknet_4_15__leaf_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5033__I _1481_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_9_i_clk clknet_4_3__leaf_i_clk clknet_leaf_9_i_clk vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_225_388 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_142_2218 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_21_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_197_218 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_68_1323 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_68_1334 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_96_706 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_178_410 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_240_358 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_206_2985 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_68_419 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_611 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7996_ _0173_ clknet_leaf_90_i_clk net135 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_2
XANTENNA__6601__A1 net29 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5404__A2 _1838_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_178_454 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_95_238 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_166_605 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_178_465 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6947_ _1231_ _1711_ _3168_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4093__B _0520_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_166_627 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_124_1995 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3966__A2 _0524_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_193_457 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_235_3337 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6878_ _2986_ _3108_ _3121_ _0327_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_91_422 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_119_554 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5168__A1 core_0.execute.rf.reg_outputs\[4\]\[7\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_349 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_716 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5168__B2 core_0.execute.rf.reg_outputs\[2\]\[7\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
X_5829_ core_0.execute.rf.reg_outputs\[1\]\[5\] _1615_ _2225_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6904__A2 _3135_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_151_80 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_552 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_134_524 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_146_384 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_161_310 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_134_535 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_162_855 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_32_500 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_161_332 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4540__C _1041_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_153_2347 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_17_596 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_161_354 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_134_579 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output184_I net184 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_32_533 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_79_1463 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4112__I net105 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6668__A1 _2940_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_728 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_102_454 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_246_3466 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_235_119 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_246_3477 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_216_311 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_244_631 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_246_36 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_217_856 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7093__A1 _1561_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7093__B2 _3149_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_164_2476 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_188_207 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_188_229 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_231_347 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7298__C _1736_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_200_701 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_197_763 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7396__A2 _3544_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_212_594 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_72_Left_319 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_157_627 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_95_750 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_156_115 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_67_452 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_200_767 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_200_789 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_625 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_184_457 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_94_271 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_138_863 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_41_1006 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5159__A1 core_0.dec_l_reg_sel\[2\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_37 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_125_524 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_153_833 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8257__CLK clknet_leaf_32_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_54_168 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_180_641 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_35_360 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_11_642 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_125_557 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_511 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_180_663 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_533 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_51_842 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_112_207 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_555 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_106_782 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_140_527 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_152_387 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_50_341 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput208 net208 sr_bus_data_o[8] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XPHY_EDGE_ROW_81_Left_328 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_50_374 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7320__A2 _3492_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_10_238 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_121_774 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5331__A1 core_0.execute.alu_mul_div.div_cur\[6\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_208_801 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_208_812 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4160_ _0778_ _0779_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XTAP_TAPCELL_ROW_52_1135 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3893__A1 core_0.dec_r_reg_sel\[2\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_4_37 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7084__A1 _1909_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_207_344 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4091_ _0568_ core_0.execute.rf.reg_outputs\[3\]\[0\] _0549_ _0712_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_0_65_56 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_128_2051 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_222_303 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6831__A1 core_0.execute.rf.reg_outputs\[2\]\[6\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5634__A2 _1584_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_234_174 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_164_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_188_730 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7850_ _0043_ clknet_leaf_68_i_clk core_0.fetch.out_buffer_data_instr\[27\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_19_742 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_90_Left_337 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_77_216 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6801_ _2983_ _3064_ _3077_ _0294_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_187_273 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4993_ _0782_ _0767_ _1440_ _1441_ _1442_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai31_2
X_7781_ core_0.dec_rf_ie\[4\] _1133_ _3827_ _3843_ _3852_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_147_104 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_58_463 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3944_ _0577_ _0578_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_86_783 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6732_ _2990_ _3022_ _3037_ _0265_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_85_260 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7139__A2 net214 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_86_794 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_84 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_63_1264 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_73_422 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_282 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_14_93 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5737__B core_0.decode.oc_alu_mode\[13\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6663_ _2941_ _2996_ _2997_ _0236_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_162_107 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_6_711 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_190_449 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_73_466 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_128_384 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_33_308 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5614_ _2013_ _2014_ _2015_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XTAP_TAPCELL_ROW_139_2180 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6898__A1 _2951_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_144_855 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6594_ net36 _1148_ _2943_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_26_360 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_254 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_60_127 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_131_505 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5545_ _1004_ _1956_ _1967_ _0148_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__4373__A2 _0966_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_8333_ _0509_ clknet_leaf_91_i_clk core_0.dec_l_reg_sel\[2\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__dffq_2
XTAP_TAPCELL_ROW_230_3267 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_30_81 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_170_173 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_230_3278 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_41_352 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8264_ _0440_ clknet_leaf_37_i_clk core_0.execute.sreg_scratch.o_d\[14\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5476_ _1908_ _1909_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_69_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_197_76 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5472__B _1817_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7215_ _3400_ _3401_ _3402_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_4427_ _0883_ _1028_ _1029_ _0963_ net161 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XANTENNA__5322__A1 core_0.execute.alu_mul_div.div_cur\[1\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_218_609 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8195_ _0371_ clknet_leaf_2_i_clk core_0.execute.alu_mul_div.div_res\[4\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_245_406 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7146_ _3175_ _3350_ _3351_ _3352_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__4676__A3 _1231_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5873__A2 _2264_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4358_ core_0.fetch.prev_request_pc\[13\] _0955_ _0974_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__7075__A1 core_0.execute.alu_mul_div.mul_res\[10\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
X_7077_ _3273_ _3280_ _3287_ _3288_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_4289_ _0836_ _0907_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__5625__A2 _2009_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6028_ _2412_ _2417_ _2418_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_EDGE_ROW_129_Left_376 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_198_527 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_240_122 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_213_347 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_241_667 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_213_358 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_213_369 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_179_752 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_240_177 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_178_251 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_138_104 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7979_ _0156_ clknet_leaf_39_i_clk core_0.execute.mem_stage_pc\[14\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__4107__I net70 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_178_295 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_77_772 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_166_446 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6523__S _2244_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_166_457 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4061__A1 _0533_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_193_276 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_181_416 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_193_287 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_157 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_91_252 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_92_786 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6889__A1 _2996_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_138_Left_385 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__7550__A2 _2257_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_51_127 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_691 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_842 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_122_527 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_134_387 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_161_184 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_32_352 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__7581__C _1950_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6478__B _2856_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5382__B _1817_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_102_251 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7153__I _1747_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_166_2505 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7066__A1 _1224_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_147_Left_394 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_232_601 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_205_826 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_189_538 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_99_352 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_232_667 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_220_807 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4218__S _0824_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_87_536 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_16_701 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_157_402 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_177_2634 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_74_219 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_185_788 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_55_422 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_67_282 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_95_591 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5557__B _1964_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_200_597 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_16_i_clk_I clknet_4_8__leaf_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_82_241 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_222_82 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_83_786 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_126_855 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_137_192 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7541__A2 _1398_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_42_138 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4355__A2 _0966_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5552__A1 _0991_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_141_836 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_23_352 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_141_858 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5330_ core_0.execute.alu_mul_div.div_cur\[5\] _1715_ _1778_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_106_590 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5261_ _1507_ _1512_ _1710_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_TAPCELL_ROW_188_2763 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_227_417 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_188_2774 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_7000_ core_0.execute.alu_mul_div.cbit\[3\] _3216_ _3217_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__nor2_1
Xclkbuf_4_8__f_i_clk clknet_3_4_0_i_clk clknet_4_8__leaf_i_clk vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_4212_ core_0.fetch.out_buffer_data_instr\[23\] _0831_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xclkbuf_leaf_74_i_clk clknet_4_13__leaf_i_clk clknet_leaf_74_i_clk vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_5192_ net186 net202 _1461_ _1641_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_4
XTAP_TAPCELL_ROW_110_1836 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_76_66 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4143_ core_0.ew_reg_ie\[2\] _0760_ _0549_ core_0.ew_reg_ie\[3\] _0534_ _0762_ vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_0_208_664 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5607__A2 _1600_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4074_ _0567_ core_0.execute.rf.reg_outputs\[3\]\[2\] _0548_ _0697_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_222_111 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_222_122 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_207_196 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_222_133 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_89_i_clk clknet_4_6__leaf_i_clk clknet_leaf_89_i_clk vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_7902_ _0093_ clknet_leaf_68_i_clk core_0.decode.i_imm_pass\[11\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_211_818 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_92_65 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4355__C _0963_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_203_2944 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_222_177 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_116_61 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7833_ _0026_ clknet_leaf_59_i_clk core_0.fetch.out_buffer_data_instr\[10\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_116_72 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_148_413 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_148_424 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_148_435 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_12_i_clk clknet_4_9__leaf_i_clk clknet_leaf_12_i_clk vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_148_446 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_176_755 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7764_ _1048_ _1104_ _3761_ _3778_ _3839_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_0_148_457 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4976_ core_0.execute.sreg_priv_control.o_d\[14\] _1393_ _1426_ _1390_ _1427_ vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_TAPCELL_ROW_121_1965 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5467__B _1816_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6715_ _2961_ _3021_ _3028_ _0257_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_3927_ _0558_ _0559_ _0560_ _0561_ _0562_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_4
X_7695_ _1078_ _1095_ _3795_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_163_438 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_175_298 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_191_769 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6646_ _2979_ core_0.ew_data\[10\] _2980_ net22 _2986_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XANTENNA__7532__A2 _3641_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_144_663 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_27_i_clk clknet_4_10__leaf_i_clk clknet_leaf_27_i_clk vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_15_842 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_116_365 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5543__A1 _1008_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_6_585 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_116_387 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_150_2317 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6577_ _2929_ _2930_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_14_352 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_76_1422 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_8316_ _0492_ clknet_leaf_9_i_clk core_0.dec_jump_cond_code\[1\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_2
X_5528_ _1955_ _1956_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA__5914__C _1531_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input60_I i_req_data[2] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_131_379 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5459_ _1886_ _1894_ _1373_ _1895_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_8247_ _0423_ clknet_leaf_20_i_clk net106 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_4
XFILLER_0_218_417 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_112_593 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_246_726 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5846__A2 _2209_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_8178_ _0354_ clknet_leaf_128_i_clk core_0.execute.alu_mul_div.mul_res\[4\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_243_3425 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output147_I net147 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7129_ _3335_ _3336_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_226_461 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7599__A2 _3681_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_161_2446 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6271__A2 _2486_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_214_667 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_202_807 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_241_464 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_87_1551 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_241_475 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4282__A1 core_0.fetch.prev_request_pc\[15\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_213_177 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4282__B2 core_0.fetch.prev_request_pc\[14\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_87_1562 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_243_37 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_96_333 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_139_402 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6949__I2 _1789_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7220__A1 _2440_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_139_468 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_167_777 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_422 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_49_282 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_742 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_126_107 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5782__A1 _1121_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5782__B2 _2139_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_181_224 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_92_561 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_9_390 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_855 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_37_488 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_181_257 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_18_680 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_92_594 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_107_343 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7523__A2 _3646_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_107_365 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_181_279 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_21_770 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_122_302 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_123_836 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_172_2575 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_122_335 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_123_858 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_98_1691 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_33_683 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7287__A1 _3384_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6001__B _2346_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_155_Left_402 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_237_748 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_207_3000 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_236_247 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6428__S _1625_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_205_612 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_125_2010 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_204_122 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_189_346 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6262__A2 _2646_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_160 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_204_166 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_204_177 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_99_182 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_153_48 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6671__B _2984_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_153_59 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7211__A1 _1742_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_47_208 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6014__A2 core_0.execute.sreg_irq_pc.o_d\[3\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_201_862 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_164_Left_411 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_157_232 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4830_ _1280_ net40 _1170_ _1323_ _1324_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_0_75_539 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_47_1078 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_200_383 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_107 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_145_416 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4576__A2 net157 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_8_839 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4761_ _1051_ _1283_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_185_596 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_172_213 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_338 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_145_438 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_157_298 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_60_1234 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_127_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_28_477 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_349 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6500_ _1059_ _2872_ _2594_ _2815_ _2878_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_138_490 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_126_641 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7480_ net201 _1398_ _3630_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4692_ _1243_ _0019_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7514__A2 _3640_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_136_2150 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4328__A2 _0942_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_43_458 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6431_ _2113_ _2669_ _2811_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_153_471 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_126_696 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_11_72 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_102_85 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_3_544 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_3_555 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6362_ _1059_ _2052_ _2743_ _2744_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_113_346 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_87_10 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_178_34 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_11_322 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7278__A1 _1400_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5313_ _1760_ _1761_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
X_8101_ _0277_ clknet_leaf_107_i_clk core_0.execute.rf.reg_outputs\[4\]\[8\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_2
XANTENNA__7278__B2 _1430_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_344 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_173_Left_420 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
X_6293_ _2036_ _2676_ _2677_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_87_76 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5244_ net189 net205 _1460_ _1693_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_4
X_8032_ _0209_ clknet_leaf_53_i_clk net121 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_227_225 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6846__B _3098_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5175_ _1531_ _1624_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XTAP_TAPCELL_ROW_71_1363 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4500__A2 _1078_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_208_461 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4126_ core_0.execute.pc_high_out\[6\] _0732_ _0745_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_194_77 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_194_88 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7450__A1 _3581_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6253__A2 _1620_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4057_ core_0.execute.rf.reg_outputs\[1\]\[3\] _0681_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_36_80 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_223_475 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6005__A2 _2249_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7816_ _1098_ _3874_ _1141_ _3875_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__4016__A1 _0533_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_66_539 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_422 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7753__A2 _0514_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_149_799 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_108_107 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_136_416 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_176_585 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4567__A2 core_0.ew_mem_width vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5764__A1 _1754_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7747_ core_0.decode.i_instr_l\[8\] _0514_ _1070_ _3826_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_4959_ _1414_ _0626_ _1415_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_46_241 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_108_129 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_163_224 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_46_252 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_82_1492 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_74_583 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_652 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_46_285 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_62_734 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7678_ _1042_ _1092_ _1078_ _3778_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_151_419 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_34_447 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6629_ core_0.execute.rf.reg_outputs\[7\]\[6\] _2962_ _1978_ _2973_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_105_858 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_131_110 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_171_290 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_131_132 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7269__A1 _1742_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_197_Right_197 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_120_839 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_30_664 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_30_675 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_219_737 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5819__A2 _2209_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_238_37 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6756__B _3045_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_246_556 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_218_247 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6492__A2 _2486_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_7_598 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_242_751 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_214_442 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7441__A1 _3563_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_300 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_202_626 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_201_103 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_241_294 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_97_664 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4007__A1 net102 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_96_174 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_96_185 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_38_731 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7744__A2 _0514_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_139_254 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_194_371 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_174_2604 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5755__A1 _1515_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_72_509 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4558__A2 _1066_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_84_369 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_154_235 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_25_447 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_4_319 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_142_419 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5507__A1 _1223_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_53_767 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_255 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_80_575 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_150_430 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_213_3070 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_40_428 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_80_597 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xmax_cap218 _1484_ net218 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XPHY_EDGE_ROW_164_Right_164 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__4730__A2 _1253_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_141 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_110_349 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_131_2080 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_20_174 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_148_37 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_237_534 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_185_2733 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_209_247 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_209_258 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4965__I _1283_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6483__A2 _2860_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5140__C1 core_0.execute.rf.reg_outputs\[6\]\[8\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6158__S _2123_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7680__A1 _1113_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4494__A1 _1061_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_224_217 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4494__B2 _1086_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6235__A2 _2531_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7432__A1 _3581_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_189_132 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6980_ _3192_ _3196_ _3197_ _3198_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_232_261 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7985__CLK clknet_leaf_29_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_232_272 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7497__B _3516_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5931_ _1689_ _1652_ _1559_ _2323_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__5994__A1 _2281_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_76_804 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_244_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_200_2914 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_48_506 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_244_91 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_539 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_105_1768 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_5862_ core_0.execute.pc_high_buff_out\[0\] _2249_ _2250_ core_0.execute.sreg_irq_flags.o_d\[0\]
+ core_0.execute.sreg_scratch.o_d\[0\] _2254_ _2255_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi222_2
XFILLER_0_87_196 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_196_2862 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_7601_ _3670_ _3718_ _3719_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4813_ _0866_ core_0.fetch.submitable _1313_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_185_371 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_764 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_200_191 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_185_393 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5793_ core_0.execute.rf.reg_outputs\[3\]\[1\] _1606_ _1615_ core_0.execute.rf.reg_outputs\[1\]\[1\]
+ _2193_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_145_224 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4205__I core_0.fetch.out_buffer_valid vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_8_658 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5210__A3 _0776_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7532_ _0553_ _3641_ _3661_ _0441_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_4744_ core_0.fetch.out_buffer_data_instr\[26\] net56 _1236_ _1273_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_44_734 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_56_594 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_145_268 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_43_222 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_32_898 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_7463_ core_0.execute.mem_stage_pc\[14\] _3616_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_4675_ _1227_ _1230_ _1231_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_6414_ _2346_ net197 _2784_ _2794_ _2795_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__6171__A1 _1613_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_98_75 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_141_463 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7394_ _1357_ core_0.execute.mem_stage_pc\[2\] _3559_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_98_97 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_102_839 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_113_165 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_114_699 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6345_ _2576_ _2726_ _2727_ _0188_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XPHY_EDGE_ROW_131_Right_131 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_141_496 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_12_664 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_101_349 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6276_ net87 _2531_ _2659_ _2537_ _2660_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_TAPCELL_ROW_227_3239 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_11_185 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_51_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_216_707 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8015_ _0192_ clknet_leaf_53_i_clk core_0.ew_data\[14\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_2
X_5227_ _0690_ net219 _1670_ _1675_ _1676_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XANTENNA__7671__A1 _1078_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6295__C _2638_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4485__A1 core_0.decode.i_instr_l\[6\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_209_792 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_138_81 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5158_ core_0.execute.rf.reg_outputs\[5\]\[6\] _1604_ _1605_ core_0.execute.rf.reg_outputs\[7\]\[6\]
+ _1606_ core_0.execute.rf.reg_outputs\[3\]\[6\] _1607_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_0_243_559 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_4_557 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_145_2249 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input23_I i_mem_data[11] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7423__A1 _3563_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4109_ net19 net18 core_0.execute.irq_en _0729_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__4237__A1 _0824_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5089_ core_0.execute.rf.reg_outputs\[6\]\[14\] _1435_ _1486_ core_0.execute.rf.reg_outputs\[5\]\[14\]
+ _1538_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_169_839 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5985__A1 _1603_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_84_1521 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7200__B _1414_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_78_174 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_79_697 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_149_552 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_78_185 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_238_3368 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_94_656 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_807 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_94_667 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5737__A1 _1715_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_137_736 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_191_352 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_34_211 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_35_767 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_151_216 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_156_2389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4960__A2 _1394_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_255 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_564 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_62_586 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_737 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_62_597 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6162__A1 _2022_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_132_452 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output91_I net91 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_95_1650 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_160_783 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_105_699 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_132_496 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_219_512 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_246_342 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5268__A3 _1713_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6465__A2 _2843_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_100_371 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7662__A1 _1132_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_118_18 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4476__A1 core_0.decode.i_instr_l\[3\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_206_239 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_215_751 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7414__A1 _3543_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_230_710 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4228__A1 _0726_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_215_795 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_180_2674 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_214_283 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4779__A2 _1285_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_804 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5976__A1 _1121_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_187_658 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_163 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_111 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__7717__A2 _1064_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_167_360 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_128_725 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_44_1037 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5728__A1 _2123_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_233_Right_233 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_85_689 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_183_842 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_72_317 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__7764__C _3778_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_594 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_26_745 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5565__B _1978_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_53_564 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4460_ _1034_ _1050_ _1054_ _0004_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__6153__A1 _1378_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_151_772 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_247 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_68_34 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4391_ _0951_ _1000_ _1001_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__5900__A1 _1458_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_159_58 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6130_ _1601_ _2309_ _2517_ _1831_ _2518_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_0_111_669 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_238_843 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_238_865 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_194_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_55_1177 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6456__A2 _2825_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6061_ core_0.execute.sreg_scratch.o_d\[4\] _2254_ _2264_ core_0.execute.sreg_irq_pc.o_d\[4\]
+ _2450_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__7653__A1 _3758_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8013__CLK clknet_leaf_53_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4467__A1 _1034_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5012_ _1460_ _1461_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_8
XANTENNA__7004__C _3177_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7405__A1 _1357_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_205_261 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_1_527 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_178_636 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_221_754 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_191_34 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6963_ _1439_ _1448_ _1449_ _1226_ _3183_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XANTENNA__8163__CLK clknet_leaf_89_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5967__A1 _2356_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_37_957 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_76_601 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_177_124 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_191_56 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_177_135 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5914_ _1554_ _1568_ _2305_ _1531_ _2306_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai211_2
XANTENNA__4363__C _0823_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_48_336 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6894_ _2940_ _3129_ _3131_ _0333_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__7708__A2 _1084_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_64_807 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5719__A1 _1124_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_8_411 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_76_667 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_75_155 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5845_ _2236_ _2238_ _2239_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__3993__A3 _0527_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_76_689 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_200_Right_200 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_119_758 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_712 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_8_466 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5195__A2 _1553_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6392__A1 core_0.decode.oc_alu_mode\[11\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_90_125 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_91_648 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_173_352 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_56_380 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5776_ _2072_ _2176_ _2177_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_clkbuf_leaf_64_i_clk_I clknet_4_15__leaf_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_173_374 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_99_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_EDGE_ROW_101_Left_348 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
X_7515_ core_0.execute.sreg_scratch.o_d\[7\] _3646_ _3651_ _3653_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_16_244 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_90_158 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4727_ _0840_ _1237_ _1264_ _0033_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_173_396 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_118_1926 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_71_361 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6150__I _2245_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_44_586 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7446_ _3547_ _3601_ _3602_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_114_452 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4658_ _0722_ _1216_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_114_485 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_142_794 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_9_616 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_141_282 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7377_ _3540_ _3544_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
X_4589_ _1159_ net153 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_12_461 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6328_ _2697_ _2705_ _2710_ _2711_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and3_2
XANTENNA__4819__B _1316_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6447__A2 _2579_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7644__A1 core_0.execute.pc_high_buff_out\[6\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6259_ _1059_ _2040_ _2641_ _2643_ _2644_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XTAP_TAPCELL_ROW_90_1591 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_110_Left_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_216_559 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_203_209 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_99_748 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_98_236 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_224_592 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_98_247 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_169_625 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_168_102 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5958__B2 core_0.execute.pc_high_buff_out\[2\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_212_776 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_67_623 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_196_466 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_158_2407 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4630__A1 core_0.execute.alu_flag_reg.o_d\[1\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_11_Right_11 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_177_691 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_165_842 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_54_317 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_637 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_164_341 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5186__A2 _1434_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_81_136 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_35_553 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_137_599 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_105_430 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_90_681 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_133_772 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_22_247 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6995__I core_0.execute.alu_mul_div.mul_res\[4\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6686__A2 _2999_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_169_2536 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_20_Right_20 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__7635__A1 net204 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_37 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4449__A1 _1038_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_246_172 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_209_72 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_207_559 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_234_345 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6944__B _1230_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_89_203 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_145_38 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_215_570 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7759__C core_0.decode.i_instr_l\[3\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_203_732 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_47 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_89_258 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_199_282 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_187_422 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5949__A1 core_0.dec_sreg_irt vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_230_540 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_203_754 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_202_231 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_225_60 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_58_601 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_148_809 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6610__A2 _2941_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_159_146 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_187_466 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_202_275 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3960_ _0592_ net197 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XTAP_TAPCELL_ROW_34_916 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4621__A1 core_0.execute.alu_flag_reg.o_d\[2\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_175_628 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_807 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_58_667 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_102_1738 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_3891_ _0526_ _0527_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_8
XTAP_TAPCELL_ROW_193_2832 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_57_177 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_156_853 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5630_ _1715_ _1934_ _2022_ _2031_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA__5177__A2 _1604_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_73_648 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_183_672 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_38_391 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_14_684 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5295__B _0731_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_183_694 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_241_92 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5561_ core_0.execute.mem_stage_pc\[14\] _1955_ _1964_ _1976_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_5_436 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_170_333 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_207_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_26_586 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7300_ net76 _3475_ _3476_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_14_737 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_26_597 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_692 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4512_ _1101_ _1046_ _1102_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_8280_ _0456_ clknet_leaf_27_i_clk core_0.execute.pc_high_buff_out\[1\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5492_ _1923_ _1924_ _1229_ _1925_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_170_399 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7231_ net82 _3398_ _3399_ _3415_ _3416_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__6677__A2 _3006_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_123_271 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_41_578 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_123_282 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4443_ core_0.decode.i_instr_l\[0\] _1038_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_110_96 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4374_ net73 _0987_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_0_1_675 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7162_ core_0.execute.alu_mul_div.div_res\[3\] _3363_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_186_34 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_111_477 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_113_1867 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_226_802 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7626__A1 _0735_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6113_ _2500_ _2501_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_4
X_7093_ _1561_ _1566_ _3209_ _3302_ _3149_ _3303_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai32_1
XFILLER_0_226_824 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_95_98 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_119_61 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6044_ _2419_ _2430_ _2433_ _2434_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_4
XANTENNA__5101__A2 _1549_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_119_72 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_142_2219 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_241_838 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_178_400 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_68_1324 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_206_2986 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_96_718 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_178_422 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_7995_ _0172_ clknet_leaf_89_i_clk net134 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_4
X_6946_ _1713_ _1926_ _3167_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_178_477 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_124_1996 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7685__B _1084_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_119_522 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_235_3327 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_193_447 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3966__A3 _0527_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6877_ core_0.execute.rf.reg_outputs\[1\]\[10\] _3114_ _3112_ _3121_ vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_147_842 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_165_138 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_317 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_235_3338 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_63_103 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_76_497 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_174_650 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5168__A2 _1436_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_48_199 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6365__A1 _2734_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5828_ _2202_ _2223_ _2224_ _0173_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_146_374 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_180_119 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_227 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5759_ _2149_ _2154_ _2159_ _2160_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_134_547 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_153_2348 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_44_372 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8059__CLK clknet_leaf_99_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_115_772 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_71_191 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_79_1464 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_60_865 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4128__B1 net112 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6668__A2 _2999_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_102_411 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_output177_I net177 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7429_ _3563_ net86 _3553_ _3587_ _3588_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_32_589 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_92_1620 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4679__A1 _1221_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5876__B1 _2268_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_102_499 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_246_3467 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_246_3478 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_216_334 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7093__A2 _1566_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_216_356 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6764__B _3045_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_216_378 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6840__A2 _3092_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_164_2477 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4851__A1 _0914_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_87_718 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_99_578 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_169_422 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_86_228 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_86_239 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_67_431 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_95_740 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_28_807 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5894__I core_0.decode.oc_alu_mode\[7\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_95_784 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_27_328 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_165_650 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_41_1007 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5159__A2 core_0.dec_l_reg_sel\[1\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_131_18 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_137_352 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_136 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_165_683 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_152_311 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_11_643 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_82_489 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_164_193 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_152_377 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xoutput209 net209 sr_bus_data_o[9] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA__6659__A2 _2935_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_10_206 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_58 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5331__A2 _1761_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7608__A1 core_0.execute.pc_high_buff_out\[7\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_208_824 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_52_1136 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_235_632 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3893__A2 core_0.dec_r_reg_sel\[1\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_12_i_clk_I clknet_4_9__leaf_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7084__A2 _1576_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_156_37 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4090_ _0565_ _0535_ _0536_ core_0.execute.rf.reg_outputs\[6\]\[0\] _0711_ vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_0_235_654 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6674__B _3004_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_128_2052 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_65_68 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_223_838 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_207_389 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6831__A2 _3092_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4842__A1 _1280_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_222_337 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4693__I1 net64 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_19_743 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_203_562 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_157_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6800_ core_0.execute.rf.reg_outputs\[3\]\[9\] _3070_ _3072_ _3077_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_81_45 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6595__A1 net28 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_188_786 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7780_ _1136_ _3851_ _0499_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_4992_ _0770_ _0767_ core_0.execute.rf.reg_outputs\[7\]\[0\] _1441_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_187_296 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_58_453 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6731_ core_0.execute.rf.reg_outputs\[5\]\[12\] _3027_ _3031_ _3037_ vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3943_ core_0.dec_r_reg_sel\[2\] core_0.dec_r_reg_sel\[1\] _0518_ _0577_ vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_0_129_842 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_147_138 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_317 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_46_648 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_63_1265 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_105_96 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_144_801 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_73_434 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__8201__CLK clknet_leaf_2_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6662_ core_0.execute.rf.reg_outputs\[7\]\[15\] _2935_ _2984_ _2997_ vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_116_503 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_171_620 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5613_ _1479_ _1665_ _2014_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__6898__A2 _3129_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_139_2181 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6593_ _2936_ _2940_ _2942_ _0221_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_143_344 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7725__S _1946_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_26_372 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8332_ _0508_ clknet_leaf_91_i_clk core_0.dec_l_reg_sel\[1\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__dffq_4
X_5544_ core_0.execute.mem_stage_pc\[6\] _1957_ _1964_ _1967_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_103_208 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_865 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_230_3268 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_8263_ _0439_ clknet_leaf_37_i_clk core_0.execute.sreg_scratch.o_d\[13\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5475_ core_0.execute.alu_mul_div.cbit\[0\] _1908_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
X_7214_ net79 net72 net80 _3401_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_197_66 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7919__CLK clknet_4_3__leaf_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4426_ net72 _0882_ _1029_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_8194_ _0370_ clknet_leaf_129_i_clk core_0.execute.alu_mul_div.div_res\[3\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__4369__B _0945_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1_483 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7145_ _3343_ _3339_ _3349_ _3351_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4357_ _0934_ _0942_ _0945_ _0830_ _0973_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XANTENNA__7075__A2 _3285_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4288_ _0835_ _0906_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_7076_ core_0.execute.alu_mul_div.mul_res\[9\] _3279_ _3287_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_225_142 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_198_506 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6027_ _1601_ _2414_ _2416_ _1831_ _2417_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__6822__A2 _3087_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_241_624 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_240_101 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_241_646 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4833__A1 _1280_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_240_134 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_69_718 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_178_230 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_179_764 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5389__A2 _1814_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7978_ _0155_ clknet_leaf_56_i_clk core_0.execute.mem_stage_pc\[13\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_166_403 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7783__B1 _3827_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_221_392 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_178_285 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6929_ _1915_ _1221_ _3151_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_83_209 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_138_138 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4061__A2 _0524_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6338__A1 net73 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_76_294 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_119_352 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6338__B2 _2537_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_107_536 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6889__A2 _3108_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_174_491 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_146_193 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_45_670 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_558 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_150_804 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5561__A2 _1955_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_161_174 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_242_Left_489 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_103_731 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6478__C _2332_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_102_241 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_166_2506 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_3_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_229_492 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5077__A1 _1467_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6274__B1 _2577_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4793__I _1283_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_217_698 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_205_838 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_231_123 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7102__C _1372_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_375 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_59_228 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_16_702 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_240_690 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_212_392 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_200_532 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6941__C _1367_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_185_756 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_28_615 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_67_250 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_177_2635 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_55_401 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_157_458 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_184_244 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_184_255 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6329__A1 _1088_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_83_754 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_165_480 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_629 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_222_94 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5001__A1 _1439_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_82_286 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_128 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_8_i_clk clknet_4_3__leaf_i_clk clknet_leaf_8_i_clk vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_125_377 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5552__A2 _1956_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_51_640 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_24_865 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_23_342 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_51_651 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6669__B _2984_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_140_314 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_152_174 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_2_247 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6501__A1 _1689_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5260_ core_0.decode.oc_alu_mode\[12\] _1520_ _1708_ _1709_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_11_559 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_188_2764 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_239_278 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4211_ _0723_ net59 _0829_ _0830_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_4
XFILLER_0_167_47 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5191_ _1596_ _1624_ _1639_ _1640_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_0_76_45 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_110_1837 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_167_69 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4142_ core_0.ew_reg_ie\[6\] _0760_ _0549_ core_0.ew_reg_ie\[7\] _0539_ _0761_ vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XANTENNA__5068__A1 _1513_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4073_ _0567_ core_0.execute.rf.reg_outputs\[4\]\[2\] net228 _0696_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__6804__A2 _3070_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_222_101 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7901_ _0092_ clknet_leaf_74_i_clk core_0.decode.i_imm_pass\[10\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_203_2945 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_7832_ _0025_ clknet_leaf_60_i_clk core_0.fetch.out_buffer_data_instr\[9\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_92_99 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_59_751 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7763_ _1057_ _1140_ _3796_ _3838_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_0_58_261 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_784 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_4975_ _1400_ _0563_ _1426_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_6714_ core_0.execute.rf.reg_outputs\[5\]\[4\] _3027_ _3016_ _3028_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_121_1966 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_73_220 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3926_ _0534_ _0542_ _0544_ core_0.execute.rf.reg_outputs\[5\]\[14\] _0561_ vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_4
X_7694_ _1055_ _1049_ _3794_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_190_214 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_73_242 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_128_171 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_178_Right_178 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_191_759 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_190_236 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_144_631 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_190_247 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6645_ _2936_ _2983_ _2985_ _0230_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_61_404 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_46_489 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_6_575 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6576_ core_0.ew_mem_access _2929_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XANTENNA__5543__A2 _1956_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_150_2307 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_143_174 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_150_2318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_42_651 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_6_597 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_116_399 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_143_185 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_802 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8315_ _0491_ clknet_leaf_9_i_clk core_0.dec_jump_cond_code\[0\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_76_1423 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_5527_ _0810_ _1955_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_42_684 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_131_369 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8246_ _0422_ clknet_leaf_18_i_clk core_0.execute.sreg_jtr_buff.o_d\[2\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5458_ _1892_ _1893_ _1894_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA_input53_I i_req_data[23] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_100_734 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4409_ _0835_ _0947_ _0970_ _1016_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_8177_ _0353_ clknet_leaf_129_i_clk core_0.execute.alu_mul_div.mul_res\[3\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_10_570 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5389_ core_0.execute.alu_mul_div.div_cur\[2\] _1814_ _1816_ _1834_ _1835_ vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XTAP_TAPCELL_ROW_243_3426 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_7128_ _2797_ _3328_ _3335_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__5059__A1 _1466_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4319__S _0725_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7059_ _3257_ _3271_ _3189_ _3272_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__4806__A1 _0944_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_161_2447 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4282__A2 _0827_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_87_1552 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6008__B1 _2257_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_243_16 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_96_312 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_241_487 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6534__S _2906_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6559__A1 _2209_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_559 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_96_356 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7220__A2 _3391_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6949__I3 _1752_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_210_863 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_518 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_84_529 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_96_389 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5231__A1 _1601_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3957__I net91 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_167_767 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7771__A3 _3842_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_194_575 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_182_737 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_64_242 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_135_620 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_145_Right_145 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_64_264 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_629 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_52_415 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4990__B1 _1436_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4990__C2 _1438_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_21_760 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5534__A2 _1956_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_640 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_122_314 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_134_174 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_135_697 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_172_2576 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_150_645 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_98_1692 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_150_667 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_33_695 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5298__A1 core_0.decode.o_submit vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_236_226 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_207_3001 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_236_259 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_205_602 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_37 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_245_782 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_204_101 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_125_2011 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_217_50 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_244_292 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_88_802 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_232_454 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4273__A2 _0843_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5470__A1 _1374_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_29_860 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_201_830 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_158_734 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_185_520 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4025__A2 _0594_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5222__A1 core_0.execute.rf.reg_outputs\[1\]\[2\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_157_244 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_8_807 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_218_3130 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_47_1079 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_28_423 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_592 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_306 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_55_220 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4760_ _1282_ _0048_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_200_395 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_60_1235 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_71_702 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_83_562 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_138_480 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_112_Right_112 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
X_4691_ core_0.fetch.out_buffer_data_instr\[3\] net63 _1241_ _1243_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_55_275 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_136_2140 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6430_ _2293_ _2809_ _2810_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_71_757 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_126_675 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6722__A1 _2977_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_125_163 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5525__A2 _1953_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_113_314 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_141_623 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6361_ _1686_ _2171_ _2739_ _1752_ _2742_ _2743_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai221_2
XFILLER_0_180_291 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_EDGE_ROW_49_Right_49 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_3_578 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8100_ _0276_ clknet_leaf_113_i_clk core_0.execute.rf.reg_outputs\[4\]\[7\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5312_ _1515_ _1516_ _1760_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_51_492 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_194 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_140_177 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6292_ _2164_ _2634_ _2676_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_8031_ _0208_ clknet_leaf_57_i_clk net120 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_121_380 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5243_ _1477_ _1685_ _1691_ _1692_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_0_227_259 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_208_440 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_194_34 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5174_ _1531_ _1622_ _1623_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_71_1364 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_4125_ core_0.execute.prev_pc_high\[4\] _0744_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_235_270 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_147_2280 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_223_454 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4056_ core_0.execute.rf.reg_outputs\[7\]\[3\] _0530_ _0680_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__and2_1
XPHY_EDGE_ROW_58_Right_58 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__6862__B _3112_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4264__A2 core_0.decode.i_flush vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5461__A1 core_0.execute.alu_mul_div.div_cur\[12\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_195_306 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_211_649 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xclkbuf_leaf_109_i_clk clknet_4_5__leaf_i_clk clknet_leaf_109_i_clk vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_7815_ _1139_ _1094_ _1119_ _3874_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__4016__A2 _0541_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_148_244 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_52_80 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7746_ core_0.dec_jump_cond_code\[1\] _1062_ _3825_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_46_231 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_164_737 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4958_ _1381_ _1414_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XTAP_TAPCELL_ROW_82_1493 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_163_236 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_573 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3909_ _0539_ _0542_ _0544_ core_0.execute.rf.reg_outputs\[1\]\[15\] _0545_ vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_0_46_275 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_415 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_19_489 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_62_724 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7677_ _1139_ _1094_ _3777_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4889_ _1357_ _0805_ net20 core_0.ew_submit _1358_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or4_1
XFILLER_0_191_578 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_212 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6628_ _2930_ core_0.ew_data\[6\] _2971_ _2972_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_4
XFILLER_0_116_152 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_144_461 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_15_640 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_67_Right_67 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_104_314 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_116_174 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6564__I1 core_0.ew_reg_ie\[2\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_6_383 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_116_185 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6559_ _2209_ _2893_ _2920_ _0209_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_120_807 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_132_667 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_104_369 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_30_654 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_246_502 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5941__B _2279_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_8229_ _0405_ clknet_leaf_13_i_clk core_0.execute.sreg_irq_pc.o_d\[1\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_218_237 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_168_90 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_227_760 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_100_597 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_199_601 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_7_599 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_59_i_clk_I clknet_4_14__leaf_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_227_793 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_76_Right_76 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_226_292 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_198_111 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_88_109 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7441__A2 net73 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_214_Right_214 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_214_465 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5452__A1 core_0.execute.alu_mul_div.div_cur\[11\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_97_632 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_186_317 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_96_120 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_198_177 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_186_339 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_26_830 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_57_518 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_167_531 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_85_838 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_97_698 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4007__A2 _0578_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5204__A1 _1558_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_139_244 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_127_406 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_220 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_174_2605 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_139_277 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6952__A1 core_0.decode.o_submit vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4558__A3 _1048_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_73_i_clk clknet_4_13__leaf_i_clk clknet_leaf_73_i_clk vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_154_225 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_37_253 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_562 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_38_787 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_154_247 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_108_653 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_85_Right_85 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_92_381 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_108_664 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_142_409 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_25_437 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_108_675 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_135_461 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5507__A2 _1939_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_107_174 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_135_483 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_587 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_213_3071 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_88_i_clk clknet_4_12__leaf_i_clk clknet_leaf_88_i_clk vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_123_678 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_492 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_110_317 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_122_177 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4318__I0 net69 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6468__B1 net214 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_131_2081 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_237_524 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_21_698 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_185_2734 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_11_i_clk clknet_4_9__leaf_i_clk clknet_leaf_11_i_clk vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__5140__B1 _1486_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5140__C2 _1435_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7680__A2 _1116_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_94_Right_94 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_218_771 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4494__A2 _1062_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_205_454 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_232_240 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_26_i_clk clknet_4_10__leaf_i_clk clknet_leaf_26_i_clk vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_178_807 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5443__A1 _1374_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_178_829 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4981__I _1209_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6491__I0 _0563_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5930_ _1819_ _1676_ _2322_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_220_435 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87_131 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_200_2915 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_220_457 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_158_531 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5861_ _2253_ _2254_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XTAP_TAPCELL_ROW_105_1769 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7196__A1 _1051_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_237_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7600_ _3682_ _3716_ _3717_ _3718_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_196_2863 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_14_Left_261 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
X_4812_ _0940_ _1306_ _1312_ _0070_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_8_626 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5792_ core_0.execute.rf.reg_outputs\[5\]\[1\] _1604_ _2192_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_113_30 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_146_737 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_158_597 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_7_114 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7531_ core_0.execute.sreg_scratch.o_d\[15\] _3639_ _3651_ _3661_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_145_236 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_4743_ _1272_ _0041_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_28_264 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_329 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_173_556 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_43_212 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_44_746 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_32_899 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_113_96 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_160_206 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7499__A2 _3641_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7462_ _3581_ _3615_ _0417_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_4674_ _1229_ _1230_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XANTENNA__6546__I1 _2690_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6413_ _2244_ _2793_ core_0.dec_mem_access _2794_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_43_278 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_189_67 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_114_656 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_342 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_865 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_102_807 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_114_667 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7393_ _1980_ _3558_ _0405_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__7733__S _1946_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4182__A1 _0799_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_101_306 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6344_ core_0.ew_data\[10\] _2486_ _2727_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6857__B _3098_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_113_188 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_12_676 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_23_Left_270 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
X_6275_ _2447_ _2657_ _2658_ _2659_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_12_698 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_228_546 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8014_ _0191_ clknet_leaf_53_i_clk core_0.ew_data\[13\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_2
X_5226_ _1671_ _1672_ _1673_ _1674_ _1675_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and4_2
XANTENNA__4377__B _0970_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_44_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA_clkbuf_leaf_60_i_clk_I clknet_4_14__leaf_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5157_ _0770_ _0773_ _1606_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_4
XANTENNA__5052__I _1500_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_4_558 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_98_407 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7423__A2 net85 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4108_ net37 core_0.execute.sreg_irq_flags.i_d\[2\] _0728_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_223_251 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6592__B _1978_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5088_ _0789_ core_0.execute.rf.reg_outputs\[4\]\[14\] _0779_ _1537_ vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA_input16_I i_core_int_sreg[9] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5434__A1 _1375_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4039_ _0516_ _0540_ _0518_ core_0.execute.rf.reg_outputs\[1\]\[5\] _0665_ vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_1
XTAP_TAPCELL_ROW_84_1522 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_195_136 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3996__A1 _0619_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_687 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_67_838 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_94_613 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_195_158 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7187__A1 _1748_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_93_112 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_149_564 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_109_406 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_238_3369 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_19_220 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_109_417 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6934__A1 _1223_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_109_428 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_109_439 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_562 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_192_865 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7729_ net193 core_0.decode.i_imm_pass\[9\] _1946_ _3816_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_34_201 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_124_409 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_152_718 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_297 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_156_2379 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_34_234 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_670 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_90_863 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_623 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_22_407 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_50_716 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_104_111 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_144_280 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_278 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_22_418 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_132_442 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_492 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_95_1651 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_160_795 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_output84_I net84 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6767__B _3057_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_30_451 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_104_199 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_120_659 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3920__A1 _0534_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7111__A1 _2778_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_219_546 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7662__A2 _1048_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_100_383 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_246_376 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4476__A2 core_0.decode.i_instr_l\[2\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_234_538 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_192_Left_439 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_89_418 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_215_763 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_214_240 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5425__A1 _1812_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_180_2675 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_69_142 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_202_457 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7178__A1 _1231_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_84_101 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_326 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_57_348 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_44_1038 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_85_679 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6925__A1 net94 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_128_737 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_72_307 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_38_584 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_183_865 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_5_607 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7617__I _3729_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_25_212 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_25_223 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_5_618 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_392 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_117 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7725__I0 net191 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_4_128 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_716 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_133_2110 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_80_384 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7350__A1 _1458_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7350__B2 _1549_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4164__A1 _0767_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4390_ core_0.fetch.prev_request_pc\[6\] _0950_ core_0.fetch.prev_request_pc\[7\]
+ _1000_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_238_811 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6677__B _3004_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_111_648 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_150_283 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3911__A1 core_0.dec_r_reg_sel\[1\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7102__A1 _1225_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_55_1167 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7952__CLK clknet_leaf_4_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6060_ core_0.execute.pc_high_buff_out\[4\] _2249_ _2257_ core_0.execute.pc_high_out\[4\]
+ _2448_ _2449_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XTAP_TAPCELL_ROW_55_1178 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input8_I i_core_int_sreg[1] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_187_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_225_527 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5011_ _1459_ _1460_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_84_45 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_108_30 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_240_519 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_84_89 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_1_528 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5416__A1 _1233_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_221_722 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_72 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6962_ _3173_ _3182_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_220_221 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5600__I _1676_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_37_958 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_5913_ _1554_ _1501_ _2305_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__3978__A1 _0534_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_838 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7169__A1 _3358_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6893_ net88 _3130_ _3124_ _3131_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_88_495 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_186_681 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5844_ _2227_ _2230_ _2237_ _2238_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_124_73 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_29_540 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5719__A2 _1585_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6916__A1 _2986_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_158_383 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_562 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_17_702 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_90_104 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_118_247 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5775_ _2073_ _2067_ _2176_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_146_578 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7514_ net215 _3640_ _3652_ _0432_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_161_515 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4726_ net46 _1253_ _1264_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_72_863 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_118_1927 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_161_559 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7445_ core_0.execute.mem_stage_pc\[11\] _3601_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_114_442 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7341__A1 core_0.execute.alu_flag_reg.o_d\[1\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4657_ _1172_ _1215_ _0754_ _0013_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_142_773 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_150 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4155__A1 _0773_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_141_261 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_9_617 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_102_637 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7376_ _3542_ _3543_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
X_4588_ core_0.ew_data\[0\] core_0.ew_data\[8\] net157 _1159_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_101_114 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4886__I _1283_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6327_ _2090_ _2382_ _2709_ _2626_ _2710_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_0_229_844 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7644__A2 _3731_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_216_505 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6258_ _1602_ _2642_ _2643_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_110_692 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5655__A1 _1508_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_228_387 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_216_527 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5209_ _1655_ _1656_ _1657_ _0769_ _1658_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai31_2
XTAP_TAPCELL_ROW_90_1592 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_209_590 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6189_ _2202_ _2574_ _2575_ _0184_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_99_716 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_212_711 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5407__A1 core_0.execute.alu_mul_div.div_cur\[6\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output122_I net122 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4554__C _1136_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_169_648 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5958__A2 _1385_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6080__A1 _1603_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3969__A1 _0517_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_211_276 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4630__A2 core_0.execute.alu_flag_reg.o_d\[0\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_158_2408 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_66_123 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6542__S _2906_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_137_512 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_94_454 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6907__A1 _2972_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_149_372 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_165_832 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_183_139 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_4_8__f_i_clk_I clknet_3_4_0_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_81_104 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_109_247 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_109_258 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_192_662 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7580__A1 core_0.execute.pc_high_out\[3\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4394__A1 _0883_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_62_340 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_191_183 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_118_792 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_90_660 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_180_857 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_117_291 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_50_524 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_62_384 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6135__A2 _2521_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7332__A1 _2646_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_210_3030 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_105_486 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_120_412 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_50_579 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_132_283 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_238_107 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_120_434 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_169_2537 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_30_270 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_207_516 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4449__A2 _1043_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_235_858 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_54_26 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_54_37 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_187_412 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_221_3170 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_225_50 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_202_243 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_225_72 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_203_788 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_34_917 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_202_287 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4621__A2 core_0.execute.alu_flag_reg.o_d\[0\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_202_298 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3890_ _0525_ _0526_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_58_679 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_102_1739 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_193_2833 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_57_189 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_156_865 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7571__A1 net221 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_14_685 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_5560_ _0972_ _1957_ _1975_ _0155_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_5_426 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_182_172 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_115_228 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_143_537 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_41_502 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_143_559 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_373 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_4511_ core_0.decode.i_instr_l\[5\] _1035_ _1101_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_0_79_34 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5491_ _0690_ net219 _1670_ _1675_ _1908_ _1924_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_0_102_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4700__S _1246_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7230_ _3413_ _3414_ _3415_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_13_248 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4137__A1 core_0.decode.i_flush vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4442_ _1036_ _1037_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_1_632 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7161_ _3360_ _3362_ _3357_ _0369_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_4373_ _0982_ _0966_ _0986_ _0963_ net163 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_4
X_6112_ _2298_ _2499_ _2293_ _2500_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_111_489 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_113_1868 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7626__A2 _3729_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7092_ core_0.execute.alu_mul_div.mul_res\[11\] _3300_ _3301_ _3302_ vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_95_66 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8130__CLK clknet_leaf_111_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6043_ _2296_ _2432_ _2433_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_0_95_88 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_225_346 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4860__A2 _1306_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_68_1325 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_240_349 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_206_2987 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_7994_ _0171_ clknet_leaf_89_i_clk net133 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_4
XFILLER_0_89_760 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_95_218 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_135_72 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6945_ _1915_ _1702_ _3165_ _3166_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_48_101 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_88_281 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6876_ _2983_ _3107_ _3120_ _0326_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_124_1997 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_119_534 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_235_3328 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_91_402 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5827_ net135 _2209_ _2224_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_146_342 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4390__B core_0.fetch.prev_request_pc\[7\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7562__A1 _3682_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_63_126 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_119_578 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_174_662 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_63_137 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4376__A1 _0892_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_63_159 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5758_ _2017_ _1620_ _2158_ _2159_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_60_80 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_239 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_72_671 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_134_559 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_153_2349 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_4709_ _1236_ _1253_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA__7314__A1 _1977_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_44_384 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_32_524 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_161_367 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5689_ _2089_ _2090_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_121_209 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_60_855 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_79_1465 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_7428_ _3547_ _3586_ _3587_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_20_708 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5933__C _1624_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_92_1621 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5876__A1 _2245_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5876__B2 net72 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7359_ _3525_ _3526_ _3527_ _3528_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor3_2
XTAP_TAPCELL_ROW_246_3468 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_246_3479 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_229_696 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7093__A3 _3209_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_244_655 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_244_677 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_99_524 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_164_2478 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_99_557 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_169_401 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4851__A2 _1306_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_231_349 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5240__I _1625_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6053__A1 _2346_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6780__B _3057_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_157_607 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_wire219_I _1483_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_169_478 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_197_798 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_157_629 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_149_180 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_138_865 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_137_342 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7553__A1 core_0.execute.pc_high_buff_out\[0\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_41_1008 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_55_649 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_94_295 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4367__A1 _0977_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_54_148 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_82_457 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_36_863 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_159 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_70_608 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_125_537 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_164_172 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_192_492 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_11_644 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_125_559 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_50_310 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7305__A1 _1431_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_211_85 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_773 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_112_209 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4119__A1 core_0.execute.pc_high_out\[0\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5867__A1 _1196_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_120_231 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5619__A1 _1761_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_52_1137 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_235_622 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3893__A3 _0518_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_65_47 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5095__A2 _1438_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_128_2053 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_234_165 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_179_209 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4842__A2 net43 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_236_82 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_159_Right_159 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_19_744 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_172_37 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4991_ core_0.execute.rf.reg_outputs\[5\]\[0\] _1440_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_86_730 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7792__A1 _0542_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_175_404 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_86_741 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6730_ _2988_ _3022_ _3036_ _0264_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_187_286 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3942_ net92 _0576_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__inv_2
XFILLER_0_46_616 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_73_402 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_86_785 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_58_487 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6661_ _2979_ core_0.ew_data\[15\] _2980_ net27 _2996_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XTAP_TAPCELL_ROW_63_1266 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_45_126 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_156_662 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7544__A1 _3663_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_116_515 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4358__A1 core_0.fetch.prev_request_pc\[13\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5612_ _1929_ _1683_ _2013_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_0_143_312 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_5_212 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6592_ core_0.execute.rf.reg_outputs\[7\]\[0\] _2941_ _1978_ _2942_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_139_2182 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_60_107 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_8331_ _0507_ clknet_leaf_90_i_clk core_0.dec_l_reg_sel\[0\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__dffq_4
X_5543_ _1008_ _1956_ _1966_ _0147_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_30_61 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_42_855 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_171_698 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_230_3269 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_41_343 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_83 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8262_ _0438_ clknet_leaf_39_i_clk core_0.execute.sreg_scratch.o_d\[12\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_112_721 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_124_592 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5474_ _1906_ _1907_ _0137_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_7213_ net80 net79 net72 _3400_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and3_1
X_4425_ core_0.fetch.prev_request_pc\[0\] _0851_ _0946_ _1028_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_1_440 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8193_ _0369_ clknet_leaf_2_i_clk core_0.execute.alu_mul_div.div_res\[2\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5322__A3 _1557_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4369__C _0854_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7741__S _1063_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_4_14__f_i_clk_I clknet_3_7_0_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_112_798 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7144_ _3343_ _3339_ _3349_ _3350_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_0_111_286 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4356_ net76 _0972_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XANTENNA__6865__B _3112_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_74_1395 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_7075_ core_0.execute.alu_mul_div.mul_res\[10\] _3285_ _3286_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_4287_ _0903_ _0836_ _0838_ _0904_ _0905_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__6283__A1 _2113_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6026_ _1601_ _1624_ _2415_ _2416_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_213_316 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_213_338 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_241_669 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6035__A1 _1765_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_126_Right_126 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_178_220 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7232__B1 _2482_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_6_Left_253 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_96_527 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_96_538 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_178_242 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7977_ _0154_ clknet_leaf_39_i_clk core_0.execute.mem_stage_pc\[12\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_193_212 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6928_ _1227_ _1841_ _3149_ _3150_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_49_465 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_49_476 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_76_262 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_36_104 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4061__A3 _0526_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_147_640 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6338__A2 _2531_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_9_562 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6859_ core_0.execute.rf.reg_outputs\[1\]\[2\] _3108_ _3098_ _3111_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_107_504 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_64_457 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_92_766 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_162_610 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_36_159 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_146_172 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_863 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_340 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_51_107 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_161_142 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_134_389 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_32_343 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_60_663 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_161_197 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_527 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_130_540 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_387 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_130_573 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4521__A1 _1109_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_166_2507 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6775__B _3057_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_129_i_clk_I clknet_4_0__leaf_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_244_452 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5077__A2 net181 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6026__A1 _1601_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_169_220 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_185_702 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_197_562 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_16_703 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_68_730 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_68_741 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_157_426 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_169_286 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_67_240 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_68_763 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5785__B1 _1615_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_129_128 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_177_2636 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_185_768 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_138_640 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_200_588 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7526__A1 _0592_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6329__A2 core_0.execute.alu_mul_div.mul_res\[10\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_83_766 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_165_470 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_43_619 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_265 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_153_632 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_165_492 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_70_416 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_125_334 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5001__A2 _1448_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_125_356 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_855 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_180_473 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4250__S _0724_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_121_562 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4210_ _0723_ _0828_ _0829_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_188_2765 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_228_Right_228 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_227_419 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4512__A1 _1101_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5190_ _1625_ _1631_ _1638_ _1639_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA__6685__B _3004_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_110_1827 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_110_1838 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_76_57 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4984__I core_0.execute.alu_mul_div.i_mul vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4141_ _0542_ _0544_ _0760_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_4072_ core_0.execute.rf.reg_outputs\[7\]\[2\] _0529_ _0695_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_208_699 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_223_636 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_92_34 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7900_ _0091_ clknet_leaf_74_i_clk core_0.decode.i_imm_pass\[9\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_223_669 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_78_505 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_116_30 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6017__A1 _2356_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_78_527 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_203_2946 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_7831_ _0024_ clknet_leaf_58_i_clk core_0.fetch.out_buffer_data_instr\[8\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_203_360 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7765__A1 _1068_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_25_72 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6704__I _3020_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_763 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_175_212 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7762_ _1097_ _3836_ _3837_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_4974_ _1419_ _1425_ _0119_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_58_251 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_58_273 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6713_ _3020_ _3027_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
X_3925_ _0539_ core_0.execute.rf.reg_outputs\[3\]\[14\] _0549_ _0560_ vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_2
XTAP_TAPCELL_ROW_121_1967 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_7693_ _1049_ _1139_ _1092_ _1037_ _3793_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_163_418 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_457 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6644_ core_0.execute.rf.reg_outputs\[7\]\[9\] _2962_ _2984_ _2985_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_116_312 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_521 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_73_276 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_143_142 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_310 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_144_676 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6575_ _2928_ _0217_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_171_462 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7535__I _1283_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_150_2308 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_14_332 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5526_ _1740_ _1954_ _1284_ _0142_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_8314_ _0490_ clknet_leaf_76_i_clk net184 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_4
XFILLER_0_42_663 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_76_1424 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_14_387 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_8245_ _0421_ clknet_leaf_20_i_clk core_0.execute.sreg_jtr_buff.o_d\[1\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5457_ _1797_ _1799_ _1893_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_246_706 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_112_573 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_100_724 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4408_ _0959_ _1014_ _1015_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__4503__A1 _1084_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_8176_ _0352_ clknet_leaf_128_i_clk core_0.execute.alu_mul_div.mul_res\[2\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5388_ _1375_ _1832_ _1833_ _1822_ _1834_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA_input46_I i_req_data[17] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_245_238 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7127_ _2797_ _3181_ _3334_ _0363_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_243_3427 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_4339_ core_0.fetch.prev_request_pc\[14\] _0956_ _0957_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6256__A1 _2287_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5059__A2 _0608_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7058_ _3259_ _3269_ _3270_ _3271_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_199_816 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_66_90 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_241_422 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4806__A2 _1306_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_199_849 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6009_ _2395_ _2396_ _2397_ _2398_ _2399_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_0_214_658 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_161_2448 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_87_1553 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6008__B2 core_0.execute.pc_high_out\[3\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_97_858 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_179_562 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6559__A2 _2893_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7756__A1 core_0.dec_jump_cond_code\[4\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output202_I net202 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_167_757 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_402 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_166_256 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_167_779 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_108_802 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6550__S _2906_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_181_226 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_182_749 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_135_632 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_181_237 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_18_660 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_405 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_24_107 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_107_334 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_55_i_clk_I clknet_4_14__leaf_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_118 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_52_427 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6192__B1 _2577_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_21_761 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3973__I _0604_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6731__A2 _3027_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_150_613 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_162_473 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_172_2577 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_33_652 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_663 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_98_1693 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_122_348 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_21_836 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_103_551 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_21_858 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_103_562 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5298__A2 _0801_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_236_216 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_207_3002 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6247__A1 _2010_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_69_Left_316 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_205_636 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6798__A2 _3070_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_125_2012 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_205_669 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_99_151 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_217_95 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_29_861 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_99_184 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7747__A1 core_0.decode.i_instr_l\[8\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_62_37 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_157_212 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_197_392 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5222__A2 _1615_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_233_72 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_218_3131 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_157_278 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_457 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_83_552 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_60_1236 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_4690_ _1242_ _0018_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XPHY_EDGE_ROW_78_Left_325 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_43_416 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_107 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_153_440 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_224 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_125_142 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_136_2141 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6722__A2 _3021_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_71_769 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6399__C _2332_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_153_484 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_181_793 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6360_ _1568_ _2740_ _2741_ _2742_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_102_98 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5311_ core_0.execute.alu_mul_div.div_cur\[7\] _1758_ _1759_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__or2_1
X_6291_ _1121_ _2674_ _2675_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_8030_ _0207_ clknet_leaf_57_i_clk net119 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_228_717 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6486__A1 _1380_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_87_67 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5242_ _1686_ _1687_ _1688_ _1689_ _1472_ _1690_ _1691_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai222_1
XTAP_TAPCELL_ROW_229_3260 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_5173_ _1553_ _1613_ _1621_ _1622_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XPHY_EDGE_ROW_87_Left_334 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_71_1365 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_242_208 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_208_452 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4124_ _0743_ net112 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_235_260 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_208_485 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6789__A2 _3070_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_223_422 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_147_2281 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
Xinput1 i_core_int_sreg[0] net1 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_4055_ _0679_ net204 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_127_84 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_36_82 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_79_836 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_78_313 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5461__A2 _1838_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_858 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_149_702 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_204_680 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_210_138 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_78_368 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7814_ _3793_ _3798_ _3873_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_94_839 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_176_543 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6410__A1 _1379_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4016__A3 _0543_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5213__A2 _1615_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_413 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_143_72 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4957_ _1301_ _1413_ _0114_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_93_349 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_96_Left_343 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
X_7745_ _3823_ _3824_ _0491_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_163_204 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_19_446 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_47_766 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_703 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_82_1494 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_3908_ _0543_ _0544_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_117_632 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_129_492 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4972__A1 _1400_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_191_557 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_265 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_799 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_7676_ _3663_ _3776_ _0470_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_163_248 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4888_ net37 _1357_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_116_142 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_117_665 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6627_ _2929_ _2969_ _2970_ _2971_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_0_105_816 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_62_769 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_116_164 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4724__A1 net45 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6558_ net121 _1985_ _2920_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_116_197 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_696 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5509_ _1375_ _1820_ _1941_ _1942_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_6489_ _2866_ _2867_ _2868_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_131_189 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_100_521 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8228_ _0404_ clknet_leaf_13_i_clk core_0.execute.sreg_irq_pc.o_d\[0\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_218_216 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4838__B _1170_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7214__B net80 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_8159_ _0335_ clknet_leaf_88_i_clk net96 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_4
XANTENNA__6229__A1 core_0.ew_data\[7\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_199_613 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_214_422 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_198_101 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_214_444 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_199_646 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_7_i_clk clknet_4_2__leaf_i_clk clknet_leaf_7_i_clk vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_241_263 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_202_617 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5452__A2 _1814_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_198_167 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_26_820 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_139_212 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5388__C _1822_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_96_154 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_195_863 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5204__A2 _1652_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6401__A1 _2279_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_194_351 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_167_576 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_127_418 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_174_2606 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_167_598 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4963__B2 _1391_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_80_500 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_107_142 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_53_769 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_213_3072 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_122_123 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_61_780 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_150_487 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6468__A1 _2286_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_143 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6468__B2 _1455_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_103_392 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_131_2082 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_209_216 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_185_2735 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_237_558 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_217_260 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_205_422 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6640__A1 core_0.execute.rf.reg_outputs\[7\]\[8\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_232_274 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_73_69 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_232_285 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_158_510 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_200_2916 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_5860_ _1382_ net186 _1201_ _2252_ _2253_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_0_76_839 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7196__A2 _1392_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_201_672 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4811_ core_0.decode.i_instr_l\[4\] _1307_ _1312_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_180_37 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_200_160 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_87_198 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_196_2864 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_185_362 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_349 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_118_418 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5791_ _2191_ _0169_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_185_373 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_132_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_145_204 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_185_384 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_28_232 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_118_429 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_173_524 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4742_ core_0.fetch.out_buffer_data_instr\[25\] net55 _1246_ _1272_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_7530_ _0563_ _3641_ _3660_ _0440_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__4954__A1 _1301_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_56_574 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_51 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_7_148 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_28_298 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_16_438 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7461_ core_0.execute.sreg_irq_pc.o_d\[13\] _3542_ _3614_ _3615_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_44_758 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4673_ _1228_ _1229_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_43_246 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_126_484 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6412_ _2786_ _2792_ _2793_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_98_33 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_855 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_71_588 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7392_ core_0.execute.sreg_irq_pc.o_d\[1\] _3543_ _3557_ _3558_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_3_332 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_71_599 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_114_679 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6343_ _2346_ net195 _2717_ _2725_ _2726_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_98_88 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_51_290 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6459__A1 _2576_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6274_ core_0.execute.sreg_priv_control.o_d\[9\] _1386_ _2577_ core_0.execute.sreg_irq_pc.o_d\[9\]
+ _2658_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_TAPCELL_ROW_116_1899 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_110_863 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8013_ _0190_ clknet_leaf_53_i_clk core_0.ew_data\[12\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_2
X_5225_ _0782_ _0768_ _0776_ core_0.execute.rf.reg_outputs\[2\]\[2\] _1674_ vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_0_215_208 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_209_772 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5156_ _0770_ core_0.dec_l_reg_sel\[1\] _1605_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_4
XFILLER_0_243_539 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_138_83 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_37_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6873__B _3112_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_138_94 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_236_591 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4107_ net70 _0727_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XTAP_TAPCELL_ROW_4_559 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_79_600 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5087_ core_0.execute.rf.reg_outputs\[1\]\[14\] _1484_ _1536_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6631__A1 net27 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4038_ core_0.execute.rf.reg_outputs\[6\]\[5\] _0661_ _0662_ core_0.execute.rf.reg_outputs\[5\]\[5\]
+ core_0.execute.rf.reg_outputs\[4\]\[5\] _0663_ _0664_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi222_2
XTAP_TAPCELL_ROW_84_1523 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_196_649 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3996__A2 _0624_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_78_187 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5198__A1 _0770_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5709__S _2102_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6934__A2 _1369_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5989_ _2002_ _2364_ _2368_ _2003_ _2379_ _2380_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_0_192_855 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7728_ _3815_ _0483_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4945__A1 _1301_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_62_500 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_276 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_736 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7209__B _3395_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_35_769 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7659_ core_0.dec_mem_width _1053_ _1064_ _3764_ _3765_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_34_257 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_7_693 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_144_270 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_132_421 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_120_605 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5370__A1 core_0.execute.alu_mul_div.div_cur\[1\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_95_1652 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_104_167 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3920__A2 _0535_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7111__A2 _3313_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_246_322 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output77_I net77 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_219_558 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput190 net190 sr_bus_addr[6] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_234_517 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6870__A1 _2972_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6622__A1 _2930_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_180_2676 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_187_627 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_202_436 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_186_126 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_230_778 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3987__A2 _0530_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_839 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7178__A2 _3373_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_85_625 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_97_485 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_187 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_97_496 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_168_863 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5189__A1 _1482_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_44_1039 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_182_310 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_194_181 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_26_703 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4936__A1 net201 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_194_192 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_65_360 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_758 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_842 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_4_107 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_170_527 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_182_387 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7725__I1 core_0.decode.i_imm_pass\[7\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_230_62 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_577 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_133_2111 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_163_590 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_419 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_111_605 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4164__A2 _0769_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1_836 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_110_104 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_123_487 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_110_126 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_858 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_leaf_108_i_clk clknet_4_5__leaf_i_clk clknet_leaf_108_i_clk vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__3911__A2 _0518_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_55_1168 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_226_3230 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_5010_ core_0.dec_r_bus_imm _1459_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_3
XANTENNA__6693__B _3004_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_240_509 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_206_753 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_144_2240 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6613__A1 net31 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_1_529 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_178_605 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7301__C _1735_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_233_594 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6961_ _3176_ _3181_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XTAP_TAPCELL_ROW_37_959 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_5912_ _1550_ _2301_ _2303_ _1559_ _2304_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai22_4
XFILLER_0_220_255 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_305 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3978__A2 _0535_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6892_ _3128_ _3130_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_124_41 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_75_135 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5843_ _2203_ _2231_ _2237_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_174_811 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_146_513 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_33_72 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_119_738 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6916__A2 _3130_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_29_585 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_8_457 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5774_ _2168_ _2169_ _2174_ _2175_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_146_568 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_522 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_382 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7513_ core_0.execute.sreg_scratch.o_d\[6\] _3646_ _3651_ _3652_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4725_ _0849_ _1237_ _1263_ _0032_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_17_758 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_114_410 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_71_352 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_118_1928 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_7444_ _3581_ _3600_ _0414_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_4656_ core_0.dec_jump_cond_code\[4\] _1194_ _1214_ _1204_ _1215_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_71_385 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7341__A2 _3510_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_102_605 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput70 i_req_data_valid net70 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__4155__A2 _0769_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5352__A1 core_0.execute.alu_mul_div.div_cur\[12\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
X_4587_ _1158_ net152 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_101_104 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7375_ _3541_ _3542_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_40_750 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_9_618 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_40_761 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_452 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_102_649 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5491__C _1908_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6326_ _2294_ _2545_ _2708_ _2090_ _2709_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai211_2
XANTENNA__3902__A2 _0528_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4388__B _0970_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_228_333 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6257_ _2412_ _1765_ _2642_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_228_377 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_216_517 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5208_ _0782_ _0767_ core_0.execute.rf.reg_outputs\[3\]\[3\] _1657_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__and3_1
XANTENNA__5655__A2 _1509_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6852__A1 core_0.ew_reg_ie\[1\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_72_i_clk clknet_4_13__leaf_i_clk clknet_leaf_72_i_clk vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_6188_ core_0.ew_data\[6\] _2486_ _2575_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_90_1593 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_243_358 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5139_ core_0.execute.rf.reg_outputs\[7\]\[8\] net235 _1443_ core_0.execute.rf.reg_outputs\[3\]\[8\]
+ _1588_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_0_212_701 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5407__A2 _1761_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_165_81 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_168_104 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_87_i_clk clknet_4_12__leaf_i_clk clknet_leaf_87_i_clk vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA_output115_I net115 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3969__A2 _0524_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_196_457 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4091__A1 _0568_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_66_102 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_168_159 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_636 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_158_2409 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6907__A2 _3129_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_176_170 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_54_319 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_10_i_clk clknet_4_3__leaf_i_clk clknet_leaf_10_i_clk vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_47_360 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_47_371 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7580__A2 _3672_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_63_842 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_152_505 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_152_527 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_164_387 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_35_566 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7332__A2 _2684_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_132_240 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_25_i_clk clknet_4_10__leaf_i_clk clknet_leaf_25_i_clk vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_22_238 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_132_251 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_210_3031 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5343__A1 core_0.execute.alu_mul_div.div_cur\[11\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_31_761 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_120_424 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_772 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_120_457 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_169_2538 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_219_333 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_30_282 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7096__A1 core_0.execute.alu_mul_div.mul_res\[11\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_235_804 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_235_826 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6843__A1 _2988_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_219_388 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_234_358 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_209_96 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7402__B _3545_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_234_369 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_42_Left_289 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_215_550 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_89_216 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_199_251 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_221_3160 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_98_761 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6071__A2 _2423_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_187_457 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4082__A1 _0533_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_85_400 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_98_794 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_225_95 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_34_918 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_97_282 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_230_597 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_58_658 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_156_811 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_174_107 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_128_513 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_37 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_193_2823 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_193_2834 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_85_488 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_127 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7571__A2 _3675_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_241_72 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_14_675 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_115_207 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_170_302 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_14_686 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_5_416 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_51_Left_298 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__5582__A1 _1051_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_171_836 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_241_94 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_352 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4510_ _1098_ _1099_ _1100_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_171_858 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7791__C _1133_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5490_ net217 _1650_ _1651_ _1226_ _1923_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XANTENNA__7323__A2 _3495_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_170_368 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_124_774 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_79_68 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4441_ core_0.decode.i_instr_l\[5\] _1035_ _1036_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_41_558 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3891__I _0526_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1_611 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_111_402 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6382__I0 core_0.ew_data\[11\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_9_Right_9 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_110_65 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_123_295 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_7160_ _1369_ _3358_ _3361_ _3362_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_4372_ _0965_ _0983_ _0985_ _0986_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_0_21_282 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6111_ _2498_ _2431_ _2102_ _2499_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_238_653 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_113_1869 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_226_804 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7091_ core_0.execute.alu_mul_div.mul_res\[10\] _3285_ _3290_ _3301_ vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_1_699 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_238_664 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_238_675 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_226_815 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_186_69 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5098__B1 _1486_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_238_686 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XPHY_EDGE_ROW_107_Right_107 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__5098__C2 _1435_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6834__A1 _2977_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6042_ _2431_ _2297_ _2102_ _2432_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__5637__A2 _1592_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_119_41 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_94 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_240_317 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4655__C _0753_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_233_380 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_68_1326 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_206_2988 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_7993_ _0170_ clknet_leaf_49_i_clk net132 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_178_413 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7739__S _1063_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_95_208 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_89_772 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6944_ _1915_ _1803_ _1230_ _3165_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_178_457 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4073__A1 _0567_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_647 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6875_ core_0.execute.rf.reg_outputs\[1\]\[9\] _3114_ _3112_ _3120_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_124_1998 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_146_321 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_235_3329 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_9_744 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_48_168 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_158_181 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_17_500 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_91_414 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5826_ _2219_ _2222_ _2223_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_45_842 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5573__A1 _1980_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_161_302 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5757_ _2155_ _2157_ _2158_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_17_555 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_134_527 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_146_387 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_161_313 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_566 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_115_730 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_127_590 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_161_346 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4708_ core_0.fetch.out_buffer_data_instr\[11\] _1252_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_5688_ _1479_ _2088_ _2089_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__6598__B _1978_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_79_1455 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4897__I core_0.execute.alu_mul_div.cbit\[1\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_79_1466 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4128__A2 _0742_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7427_ core_0.execute.mem_stage_pc\[8\] _3586_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_142_571 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4639_ net185 net178 _1197_ _1198_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_2
XTAP_TAPCELL_ROW_92_1611 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_13_772 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_8_93 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_92_1622 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_229_620 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7358_ _2854_ _2888_ _3527_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_102_457 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_229_653 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6309_ core_0.ew_data\[9\] _2486_ _2693_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7289_ net74 _3454_ net75 _3466_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__5089__B1 _1486_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_246_3469 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_217_826 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6825__A1 _2956_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_228_174 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_228_185 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_216_325 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_216_336 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4846__B _1170_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_216_347 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_232_807 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_164_2479 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_212_531 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_240_862 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_196_221 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_197_788 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_157_619 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_212_597 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_200_737 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_67_433 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_67_444 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_156_107 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_55_617 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_94_263 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_67_488 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_138_855 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_41_1009 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_137_354 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7942__CLK clknet_leaf_43_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_125_i_clk_I clknet_4_1__leaf_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_164_140 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4367__A2 _0966_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_125_516 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_35_352 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_125_549 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_153_858 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_209_Right_209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_23_503 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_11_645 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_51_812 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_62_160 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_62_171 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_140_519 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_23_547 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_2_419 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4119__A2 net105 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_62_193 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5316__A1 _1461_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_180_699 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_105_273 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_239_417 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_377 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_295 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7116__C _1367_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_121_766 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_120_243 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_219_152 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5619__A2 _2019_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_52_1138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_234_100 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_65_26 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_207_336 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_128_2043 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_128_2054 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_234_177 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_222_317 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_188_711 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_141_2210 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7241__A1 _3384_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_19_745 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_77_208 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4990_ core_0.execute.rf.reg_outputs\[6\]\[0\] _1435_ _1436_ core_0.execute.rf.reg_outputs\[4\]\[0\]
+ core_0.execute.rf.reg_outputs\[2\]\[0\] _1438_ _1439_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_0_188_788 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_187_254 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_98_591 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7792__A2 _1134_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_187_265 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_230_383 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_69 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3941_ _0571_ _0572_ _0573_ _0574_ _0575_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_0_105_43 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_606 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_18_308 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6660_ _2941_ _2994_ _2995_ _0235_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_39_680 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_58_499 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_63_1267 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_45_138 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_155_151 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_171_600 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_27_842 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5611_ _2010_ _2011_ _2012_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_128_376 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_5_202 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_116_527 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_128_387 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4602__I0 core_0.ew_data\[7\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_212_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6591_ _2935_ _2941_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XTAP_TAPCELL_ROW_139_2183 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_26_352 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_171_644 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8330_ _0506_ clknet_leaf_91_i_clk core_0.dec_r_reg_sel\[2\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__dffq_4
X_5542_ core_0.execute.mem_stage_pc\[5\] _1957_ _1964_ _1966_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_41_311 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_257 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_480 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_112_700 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5307__A1 core_0.execute.alu_mul_div.div_cur\[9\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
X_8261_ _0437_ clknet_leaf_37_i_clk core_0.execute.sreg_scratch.o_d\[11\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5473_ core_0.execute.alu_mul_div.div_cur\[15\] _1812_ _1841_ _1907_ vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_170_187 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_112_733 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4424_ _1024_ _0970_ _1026_ _1027_ _0877_ net168 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi221_4
X_7212_ _1172_ _1739_ _1734_ _3399_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_0_10_720 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8192_ _0368_ clknet_leaf_129_i_clk core_0.execute.alu_mul_div.div_res\[1\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4355_ _0964_ _0966_ _0969_ _0971_ _0963_ net166 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi221_4
X_7143_ core_0.execute.alu_mul_div.mul_res\[15\] _3348_ _3349_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_111_298 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_74_1396 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6807__A1 _2990_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7074_ _1372_ _1224_ _1928_ _3284_ _3285_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai31_4
XFILLER_0_39_93 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4286_ core_0.fetch.prev_request_pc\[6\] _0904_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_214_807 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7042__B _3189_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7480__A1 net201 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6025_ _2315_ _2321_ _1603_ _2415_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_198_508 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_198_519 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_240_114 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_709 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6881__B _3112_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_241_3399 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_96_506 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7232__A1 _1430_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6035__A2 _1665_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7232__B2 _3391_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_240_169 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7976_ _0153_ clknet_leaf_55_i_clk core_0.execute.mem_stage_pc\[11\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_221_361 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7783__A2 _1133_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6927_ core_0.decode.o_submit _1088_ _3149_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_4
XFILLER_0_76_230 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_77_764 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_193_224 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_606 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_166_438 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_178_298 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xclkbuf_4_13__f_i_clk clknet_3_6_0_i_clk clknet_4_13__leaf_i_clk vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_37_628 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_488 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6858_ _2946_ _3107_ _3110_ _0318_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_193_268 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5809_ _2204_ _2207_ _2208_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_6789_ core_0.execute.rf.reg_outputs\[3\]\[4\] _3070_ _3057_ _3071_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_17_352 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5717__S _1554_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_135_858 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_51_119 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_160 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_17_385 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7299__A1 _1742_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_44_193 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_output182_I net182 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6121__B _1458_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_60_675 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_102_210 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_107_Left_354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__4420__I net79 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_4_290 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_102_232 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_32_399 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_103_788 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4521__A2 _1062_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_166_2508 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_217_623 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6274__A2 _1386_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7471__A1 _3547_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_244_464 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_217_678 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_205_818 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_51_i_clk_I clknet_4_12__leaf_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_204_317 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_216_177 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6026__A2 _1624_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_213_862 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_208 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_116_Left_363 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_16_704 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7774__A2 _3842_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_129_107 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5785__A1 core_0.execute.rf.reg_outputs\[3\]\[0\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_184_213 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_68_775 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_177_2637 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5200__B _1446_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_138_630 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_67_274 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_68_797 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_82_200 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_126_803 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_138_663 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7526__A2 _3641_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_127 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8120__CLK clknet_leaf_103_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_683 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_3_706 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_480 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_35_193 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_125_Left_372 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_2_227 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4330__I core_0.fetch.prev_request_pc\[3\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_192_Right_192 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_121_585 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_227_409 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_188_2766 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4512__A2 _1046_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_208_601 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_110_1828 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_4140_ core_0.ew_reg_ie\[4\] _0520_ _0758_ core_0.ew_reg_ie\[5\] _0759_ vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_0_207_133 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_208_667 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5068__A3 _1515_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6265__A2 _0798_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7462__A1 _3581_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4071_ _0532_ _0523_ _0526_ core_0.execute.rf.reg_outputs\[6\]\[2\] _0694_ vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_1
XANTENNA__4276__A1 core_0.fetch.prev_request_pc\[11\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_134_Left_381 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_162_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__7214__A1 net79 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_204_862 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4706__S _1246_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7830_ _0023_ clknet_leaf_58_i_clk core_0.fetch.out_buffer_data_instr\[7\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_222_169 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_203_2947 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_78_539 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_116_53 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_231_681 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_148_405 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7761_ _1038_ _3760_ _1116_ _3835_ _3836_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai211_2
X_4973_ core_0.execute.sreg_priv_control.o_d\[13\] _1393_ _1424_ _1390_ _1425_ vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_TAPCELL_ROW_199_2895 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4823__I0 _0936_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_628 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6712_ _2956_ _3021_ _3026_ _0256_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_73_200 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3924_ _0539_ core_0.execute.rf.reg_outputs\[4\]\[14\] _0520_ _0559_ vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_129_652 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_86_594 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_121_1968 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_7692_ _3790_ _3791_ _3792_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__7517__A2 _3646_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_117_814 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_191_739 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6643_ _1963_ _2984_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_41_72 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_73_266 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_117_858 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_171_430 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6720__I _1963_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_143_Left_390 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__4200__A1 _0725_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6574_ core_0.dec_rf_ie\[7\] core_0.ew_reg_ie\[7\] _2201_ _2928_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_143_154 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_150_2309 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_132_839 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_8313_ _0489_ clknet_leaf_77_i_clk net183 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_2
X_5525_ core_0.execute.mem_stage_pc\[0\] _1953_ _1954_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4751__A2 _1238_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_30_804 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_14_355 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_42_675 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_76_1425 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_131_338 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_112_541 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_8244_ _0420_ clknet_leaf_20_i_clk core_0.execute.sreg_jtr_buff.o_d\[0\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5456_ _1796_ _1800_ _1891_ _1892_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_67_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_4407_ _0909_ _1009_ _1014_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__4503__A2 _1092_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_8175_ _0351_ clknet_leaf_124_i_clk core_0.execute.alu_mul_div.mul_res\[1\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5700__A1 _1596_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1_282 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5387_ _1374_ _1826_ _1833_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_7126_ _3189_ _3333_ _3334_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_243_3428 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_4338_ core_0.fetch.prev_request_pc\[13\] _0955_ _0956_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_10_594 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_5_72 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_input39_I i_req_data[10] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7453__A1 _3563_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5059__A3 _0613_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_226_453 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4269_ core_0.fetch.prev_request_pc\[12\] _0823_ _0830_ core_0.fetch.prev_request_pc\[13\]
+ _0887_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
Xclkbuf_3_5_0_i_clk clknet_0_i_clk clknet_3_5_0_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_7057_ _3259_ _3269_ _3175_ _3270_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__4267__A1 _0723_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_66_80 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_157_93 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_214_637 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6008_ core_0.execute.sreg_scratch.o_d\[3\] _2254_ _2257_ core_0.execute.pc_high_out\[3\]
+ _2398_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_213_136 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_161_2449 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6008__A2 _2254_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7205__A1 _1381_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_241_467 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_87_1554 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_96_314 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_241_489 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4019__A1 net101 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7756__A2 _3766_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_139_416 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5767__A1 _2161_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8143__CLK clknet_leaf_119_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7959_ _0137_ clknet_leaf_17_i_clk core_0.execute.alu_mul_div.div_cur\[15\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_210_865 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5020__B _1467_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_37_414 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_65_723 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_135_600 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_182_728 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_360 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_80_704 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_382 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_80_715 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4990__A2 _1435_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7873__D core_0.fetch.submitable vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_64_266 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_181_249 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_190_750 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_92_597 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8293__CLK clknet_leaf_12_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6192__A1 core_0.execute.pc_high_out\[7\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6192__B2 core_0.execute.sreg_irq_pc.o_d\[7\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_21_762 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_135_677 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_123_828 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_135_699 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_172_2578 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_98_1683 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5790__I1 _2188_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_98_1694 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4150__I core_0.dec_l_reg_sel\[0\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6786__B _3057_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_130_360 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_236_228 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_236_239 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_245_740 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7444__A1 _3581_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6247__A2 _2013_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_217_486 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_125_2013 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_88_804 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_217_85 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_153_18 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_201_810 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_29_862 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7747__A2 _0514_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_212_191 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_201_854 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_157_235 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_185_566 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_218_3132 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_68_594 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_185_588 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_222 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_55_233 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_166_791 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_60_1237 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_70_203 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_125_132 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6183__A1 core_0.execute.alu_mul_div.div_cur\[6\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_136_2142 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_181_772 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_70_247 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_140_102 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_125_187 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_153_496 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5930__A1 _1819_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_113_338 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_3_547 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5310_ _1513_ _1514_ _1758_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_4
XFILLER_0_23_174 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_11_314 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6290_ _2048_ _2629_ _2039_ _2674_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_178_37 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_23_196 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6696__B _3016_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5241_ core_0.decode.oc_alu_mode\[6\] _1690_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_3
XFILLER_0_227_206 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_121_382 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4497__A1 _1088_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_229_3261 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_5172_ _1553_ _1620_ _1621_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_71_1366 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7435__A1 _3563_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4123_ core_0.execute.pc_high_out\[4\] _0732_ _0743_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_194_69 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_147_2271 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_147_2282 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
Xinput2 i_core_int_sreg[10] net2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4054_ _0672_ _0677_ _0678_ _0679_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_235_294 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8166__CLK clknet_leaf_88_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_61 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_72 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_78_336 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_176_500 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_94_807 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_7813_ _1034_ _3863_ _3872_ _0511_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__5749__A1 _2010_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_176_522 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_203_191 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7744_ core_0.decode.i_instr_l\[7\] _0514_ _1070_ _3824_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_4956_ core_0.execute.sreg_priv_control.o_d\[8\] _1394_ _1412_ _1391_ _1413_ vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_74_520 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_136_408 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_163_216 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_46_244 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3907_ _0518_ _0543_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_8
XTAP_TAPCELL_ROW_82_1495 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_7675_ core_0.dec_sreg_load _3766_ _3775_ _3776_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__4972__A2 _0580_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_7_842 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4887_ _1356_ _0101_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_144_430 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_62_737 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6626_ net33 _1149_ _2970_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6174__A1 _1600_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_74_597 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_61_236 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_6_363 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_247 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_699 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_172_794 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6557_ _2919_ _0208_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4724__A2 _1253_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5921__A1 _1625_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_171_282 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_601 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_132_647 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_42_461 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_612 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5508_ _1223_ _1922_ _1940_ _1941_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_4
X_6488_ _2834_ _2865_ _2243_ _2867_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_219_718 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5134__C1 core_0.execute.rf.reg_outputs\[6\]\[9\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_30_667 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6477__A2 _2855_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7674__A1 _1133_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_8227_ _0403_ clknet_leaf_24_i_clk core_0.execute.irq_en vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_219_729 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_112_382 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5439_ _1876_ _1877_ _0132_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__4488__A1 _1037_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_246_526 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_218_228 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8158_ _0334_ clknet_leaf_88_i_clk net95 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_4
XANTENNA__6229__A2 _2486_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7426__A1 _3581_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7109_ _3189_ _3317_ _3318_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_199_603 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8089_ _0265_ clknet_leaf_99_i_clk core_0.execute.rf.reg_outputs\[5\]\[12\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5988__A1 _1480_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_198_124 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_303 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_199_669 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_97_623 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_241_286 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_69_336 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4660__A1 _1217_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_198_179 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_186_319 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_201_139 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_26_821 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_84_306 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_194_330 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_167_544 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_96_177 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_210_673 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_194_363 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_139_279 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_239_Left_486 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_46_1070 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_37_244 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4963__A2 _1394_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_154_238 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_203_65 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_277 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_135_441 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_163_772 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_52_247 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_567 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_122_102 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_409 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_123_636 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_150_422 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5912__B2 _1559_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_107_198 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_213_3073 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5905__S _1625_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8039__CLK clknet_leaf_81_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_60_291 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_20_133 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6468__A2 _1713_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7665__A1 _1066_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_131_2083 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4479__A1 _1069_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_177 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_185_2736 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_209_239 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5140__A2 net218 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7417__A1 _3563_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_224_209 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_218_795 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6963__C _1226_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_6_590 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_232_220 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_189_124 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6640__A2 _2962_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_87_100 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_205_489 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4651__A1 _1209_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_220_437 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_244_72 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_220_448 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_200_2917 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_76_807 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_88_667 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_158_522 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4810_ _1040_ core_0.fetch.submitable _1311_ _0069_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_158_555 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_200 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_75_339 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7794__C _1279_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_196_2865 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4403__A1 _0959_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5790_ core_0.ew_addr_high\[0\] _2188_ _2190_ _2191_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_8_617 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_756 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4741_ _1271_ _0040_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_90_309 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_173_536 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3894__I _0529_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_7_127 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_138 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_125_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_44_726 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_417 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_737 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_56_597 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_71_523 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7460_ _0580_ _3546_ _3541_ _3613_ _3614_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_22_85 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_4_801 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4672_ core_0.execute.alu_mul_div.cbit\[1\] _1228_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__inv_2
X_6411_ _1380_ _2790_ _2791_ _2792_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_113_113 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_126_496 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_153_282 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_7391_ _0709_ _3544_ _3545_ _3556_ _3557_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_189_69 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_113_135 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6342_ _2244_ _2724_ core_0.dec_mem_access _2725_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_113_157 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_101_308 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_12_645 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_11_133 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_12_667 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6273_ core_0.execute.sreg_scratch.o_d\[9\] _2579_ _2534_ net16 _2657_ vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_TAPCELL_ROW_149_2300 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_8012_ _0189_ clknet_leaf_49_i_clk core_0.ew_data\[11\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_2
X_5224_ _0771_ core_0.execute.rf.reg_outputs\[4\]\[2\] _0779_ _1673_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__5131__A2 _1438_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_243_507 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_209_762 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7408__A1 core_0.execute.sreg_irq_pc.o_d\[4\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5155_ _0782_ _0767_ _1604_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_4106_ _0725_ _0726_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
X_5086_ _1533_ _1534_ _1535_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_223_231 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_clkbuf_leaf_98_i_clk_I clknet_4_7__leaf_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_211_404 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4037_ _0532_ _0519_ _0663_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_0_79_623 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4642__A1 net187 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_2_73 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_84_1524 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_177_842 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_66_317 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_78_177 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_149_544 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_4_1__f_i_clk clknet_3_0_0_i_clk clknet_4_1__leaf_i_clk vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_137_706 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5198__A2 _0767_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_380 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6395__A1 _1107_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5988_ _1480_ _2372_ _2378_ _1684_ _2379_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_109_419 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_81_309 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7727_ net192 core_0.decode.i_imm_pass\[8\] _1946_ _3815_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4939_ _1400_ net212 _1401_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_35_715 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_191_344 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_62_523 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_748 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_34_225 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7658_ _1043_ _3760_ _3763_ _3764_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_35_759 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_145_772 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_34_247 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_865 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_117_474 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_144_260 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_707 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6609_ _2930_ core_0.ew_data\[3\] _2955_ _2956_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_4
XTAP_TAPCELL_ROW_31_890 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_6_171 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6698__A2 _2998_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7589_ _3673_ _3707_ _3708_ _1950_ _0451_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_15_461 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5952__C _2242_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5370__A2 _1603_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_95_1653 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_132_488 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_442 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7647__A1 net216 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_113_680 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_101_842 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3920__A3 _0536_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput180 net180 sr_bus_addr[11] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
Xoutput191 net191 sr_bus_addr[7] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_206_209 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6556__S _2189_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6870__A2 _3107_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_227_581 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4881__A1 _0827_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_214_220 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_199_422 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_230_702 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_215_787 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6622__A2 core_0.ew_data\[5\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_100 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_180_2677 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_159_319 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_807 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_69_155 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5189__A2 _1637_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_167_352 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_104_1760 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_38_531 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_194_160 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_167_396 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4936__A2 _1398_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6304__B _2279_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4603__I _1166_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_25_203 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_597 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_441 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_65_394 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6138__A1 _1117_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_92_191 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_247 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_123_400 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6689__A2 _3006_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_123_422 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_133_2112 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_68_37 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7638__A1 _0748_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_486 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6310__A1 _2576_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5113__A2 _1438_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_55_1169 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_226_3220 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7789__C _1133_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_218_592 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_108_32 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3889__I _0518_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_144_2241 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_233_562 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_205_253 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_1_519 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_108_65 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_205_264 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_206_798 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6960_ core_0.execute.alu_mul_div.mul_res\[1\] _3180_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_221_746 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5911_ _1542_ _2302_ _1482_ _2303_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_159_831 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_177_127 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_242_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__3978__A3 _0536_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6891_ _3128_ _3129_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_159_842 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_186_650 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_76_637 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6377__A1 _1380_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5842_ _0638_ _1444_ _1614_ _2236_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_8_403 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_201_492 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_29_542 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_29_553 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_237_3360 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_124_97 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5773_ _2171_ _2173_ _2174_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_7512_ _0722_ _3651_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
X_4724_ net45 _1253_ _1263_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6129__A1 _1601_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_127_772 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_16_236 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_247 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_72_865 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_173_399 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7443_ core_0.execute.sreg_irq_pc.o_d\[10\] _3542_ _3599_ _3600_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_44_578 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_118_1929 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_155_2370 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_4655_ net106 _1207_ _1213_ _0753_ _1214_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai211_4
XFILLER_0_31_206 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput60 i_req_data[2] net60 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_4_664 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_114_466 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput71 i_rst net71 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_4_675 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5352__A2 _1701_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7374_ _1953_ _3540_ _0731_ _3541_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_4
X_4586_ core_0.ew_data\[7\] net157 _1158_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_4_686 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_141_263 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7629__A1 _3732_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_9_619 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6325_ _2123_ _2706_ _2707_ _2294_ _2708_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_0_101_138 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_110_650 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_497 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6256_ _2287_ _2164_ _2640_ _2641_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__5104__A2 _1552_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_149_72 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6884__B _3124_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_81 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5207_ core_0.execute.rf.reg_outputs\[7\]\[3\] _1605_ _1656_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__5655__A3 _2053_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6852__A2 _2934_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_244_849 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_209_570 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6187_ _2346_ net206 _2573_ _2574_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__4863__A1 core_0.decode.i_imm_pass\[7\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_90_1594 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_5138_ _0789_ core_0.execute.rf.reg_outputs\[4\]\[8\] _0779_ _1587_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA_input21_I i_mem_data[0] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_165_60 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6604__A2 _2941_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5069_ _1466_ net189 _1518_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_169_617 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_211_212 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_196_425 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3969__A3 _0527_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_67_615 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4091__A2 core_0.execute.rf.reg_outputs\[3\]\[0\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6368__A1 core_0.execute.alu_mul_div.div_res\[11\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_183_108 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_164_311 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_181_92 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_164_333 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_192_653 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_192_664 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_118_761 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_124_208 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_191_163 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_331 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_662 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_23_718 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_132_230 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_210_3032 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_50_559 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5343__A2 _1752_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_160_594 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_169_2539 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7096__A2 _3300_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_246_142 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6794__B _3072_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_235_838 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_234_304 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6843__A2 _3087_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_121_i_clk_I clknet_4_3__leaf_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4854__A1 core_0.decode.i_imm_pass\[3\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6056__B1 _2265_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_215_562 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_203_702 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5203__B _1651_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_89_239 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8227__CLK clknet_leaf_24_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_221_3161 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_230_532 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_199_296 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_225_63 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_97_250 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_159_138 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4082__A2 _0524_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_230_576 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_202_267 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_34_919 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_85_412 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_434 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_156_801 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_193_2824 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_155_322 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_167_182 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_167_193 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_361 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_383 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_394 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_26_534 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_14_676 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_182_152 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_109_772 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_155_377 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5582__A2 _1953_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_183_686 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_81_640 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_170_314 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_54_865 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_46_i_clk_I clknet_4_9__leaf_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_170_336 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_161 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4440_ core_0.decode.i_instr_l\[6\] core_0.decode.i_instr_l\[4\] _1035_ vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_0_151_594 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_111_436 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4371_ _0946_ _0954_ _0984_ _0985_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_0_111_469 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6110_ _2104_ _2098_ _1625_ _2498_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_186_37 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_7090_ _1222_ _3204_ _3299_ _3300_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_237_142 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_192_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6834__A2 _3086_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6041_ _2107_ _2105_ _1482_ _2431_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__4845__A1 _0726_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_28_73 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_240_307 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_68_1327 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_7992_ _0169_ clknet_leaf_49_i_clk core_0.ew_addr_high\[0\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__7795__B1 _1092_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_206_2989 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6943_ _3163_ _3164_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_49_615 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5270__A1 _1543_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_626 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_178_469 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6874_ _2981_ _3107_ _3119_ _0325_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_9_712 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_124_1999 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_5825_ _2220_ _2221_ _2222_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_174_631 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_8_222 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_64_629 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_119_558 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_151_40 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_8_244 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_29_383 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_692 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_60 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_63_139 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_174_675 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5756_ _2156_ _2019_ _2157_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5573__A2 _0748_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6770__A1 _2990_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_106_219 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_151_84 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6879__B _3112_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_97_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_134_539 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_173_174 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4707_ _1251_ _0026_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_72_662 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_504 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5687_ _1124_ _1700_ _2088_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_79_1456 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_130_701 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7426_ _3581_ _3585_ _0411_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_4_461 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_194 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_102_403 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4638_ net189 net188 net191 net190 _1197_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or4_4
XANTENNA_input69_I i_req_data[9] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_130_734 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_92_1612 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_7357_ _2711_ _2747_ _3526_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_4569_ _1148_ _1149_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__inv_2
XFILLER_0_229_632 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6308_ _0626_ _2691_ _2242_ _2692_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_40_592 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_294 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7288_ _3460_ _3461_ _3465_ _0393_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_246_3459 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_228_142 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__7503__B _3516_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6239_ _2616_ _2622_ _2624_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__6825__A2 _3086_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4836__A1 core_0.decode.i_instr_l\[13\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5884__I0 core_0.ew_data\[0\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6589__A1 _2930_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_559 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_169_403 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_224_381 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_212_521 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_197_767 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_79_261 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_212_576 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_94_231 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_leaf_107_i_clk clknet_4_4__leaf_i_clk clknet_leaf_107_i_clk vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_67_456 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_95_765 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_629 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5013__A1 _1461_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_101_1730 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_165_642 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_153_804 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_180_601 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_47_180 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_137_377 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6761__A1 _2981_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_152_303 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_153_837 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_865 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6789__B _3057_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_164_174 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_165_697 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_173_Right_173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_152_325 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_11_646 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_164_196 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_515 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_695 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_180_667 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_50_312 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_106_775 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_23_559 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5316__A2 net213 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_133_572 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7710__B1 _3758_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_189_Left_436 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_120_255 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_208_816 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7413__B _3516_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_52_1139 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_207_348 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_128_2044 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_65_49 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_141_2200 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_188_734 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_188_745 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6044__A3 _2433_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_19_735 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_198_Left_445 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_19_746 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_58_401 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_188_778 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_230_373 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_175_406 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3940_ _0534_ _0535_ _0536_ core_0.execute.rf.reg_outputs\[6\]\[13\] _0574_ vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_0_187_277 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_105_55 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_86_798 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_426 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_63_1268 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_156_664 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5610_ _1695_ _1637_ _2011_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_6_715 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6590_ _2930_ core_0.ew_data\[0\] _2939_ _2940_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_4
XANTENNA__5555__A2 _1955_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_171_612 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_leaf_71_i_clk clknet_4_13__leaf_i_clk clknet_leaf_71_i_clk vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__4602__I1 core_0.ew_data\[15\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_26_342 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_737 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_EDGE_ROW_140_Right_140 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_42_802 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_662 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_139_2184 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_170_111 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_26_364 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5541_ _1013_ _1956_ _1965_ _0146_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_205_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_121_65 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_131_509 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_171_678 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_81_492 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_152_2340 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_8260_ _0436_ clknet_leaf_36_i_clk core_0.execute.sreg_scratch.o_d\[10\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__6504__A1 _2294_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5307__A2 _1754_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5472_ core_0.execute.alu_mul_div.div_cur\[14\] _1814_ _1817_ _1905_ _1906_ vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_170_177 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6211__C _2412_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_356 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7211_ _1742_ _3397_ _3398_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_0_124_594 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4423_ _0842_ _0947_ _0970_ _1027_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_111_222 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_8191_ _0367_ clknet_leaf_3_i_clk core_0.execute.alu_mul_div.div_res\[0\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_112_756 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_86_i_clk clknet_4_12__leaf_i_clk clknet_leaf_86_i_clk vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_22_581 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_10_732 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7142_ _3249_ _3347_ _1372_ _3348_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4354_ _0847_ _0947_ _0970_ _0971_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_1_475 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_39_50 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6268__B1 _2652_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_72 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_83 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_10_787 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_74_1397 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6807__A2 _3065_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7323__B _1955_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7073_ _1367_ _1937_ _3283_ _1372_ _3284_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_0_226_635 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4285_ core_0.fetch.prev_request_pc\[5\] _0903_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__inv_1
XANTENNA__4818__A1 _0935_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6024_ _2308_ _2413_ _1596_ _2414_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__7480__A2 _1398_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_207_860 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4294__A2 _0860_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_241_649 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5618__I0 net100 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_240_137 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_7975_ _0152_ clknet_leaf_55_i_clk core_0.execute.mem_stage_pc\[10\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_12_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_96_529 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_179_756 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_leaf_24_i_clk clknet_4_8__leaf_i_clk clknet_leaf_24_i_clk vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_178_244 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7549__I _3672_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_412 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6926_ _2996_ _3130_ _3148_ _0348_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_166_406 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_194_737 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6991__A1 _3149_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_76_242 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6857_ core_0.execute.rf.reg_outputs\[1\]\[1\] _3108_ _3098_ _3110_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_119_344 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_147_653 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_202_Left_449 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_91_212 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5808_ _2205_ _2206_ _2207_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_146_152 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xclkbuf_leaf_39_i_clk clknet_4_11__leaf_i_clk clknet_leaf_39_i_clk vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_45_640 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6743__A1 _2940_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6788_ _3063_ _3070_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_134_314 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_18_865 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_3_1_0_i_clk clknet_0_i_clk clknet_3_1_0_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_146_174 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_162_634 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5739_ _1439_ _1448_ _2140_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__6402__B _2782_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_150_807 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_162_667 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_695 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7299__A2 _3467_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_142_380 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_102_222 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4506__B1 _1095_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7409_ _3543_ _3570_ _3571_ _0408_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA_output175_I net175 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8072__CLK clknet_leaf_103_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_130_597 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_166_2509 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_211_Left_458 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_187_91 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_216_101 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5532__I net80 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4809__A1 _0870_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_217_646 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__7471__A2 net78 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_244_454 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_99_323 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4148__I core_0.dec_l_reg_sel\[1\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6564__S _1985_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_242_Right_242 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_240_660 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_16_705 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_212_373 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_212_384 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_200_524 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_185_726 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_67_220 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_184_203 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6982__A1 _1908_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5785__A2 _1606_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_157_428 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_220_Left_467 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_83_702 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_177_2638 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_184_247 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_82_212 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_95_595 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_138_675 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_139 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6734__A1 _2992_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5537__A2 _1172_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_651 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_70_407 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4596__I0 core_0.ew_data\[4\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_802 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_137_196 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_153_656 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7408__B _3516_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_125_358 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_152_144 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_51_621 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_51_632 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_63_492 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_140_317 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_23_345 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_152_177 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_106_594 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_239_204 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_133_380 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_121_542 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_188_2767 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_121_597 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_76_37 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_110_1829 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_76_59 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4070_ core_0.execute.rf.reg_outputs\[2\]\[2\] _0691_ _0662_ core_0.execute.rf.reg_outputs\[5\]\[2\]
+ _0692_ core_0.execute.rf.reg_outputs\[1\]\[2\] _0693_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XANTENNA__4276__A2 _0854_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5473__A1 core_0.execute.alu_mul_div.div_cur\[15\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_235_487 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_204_830 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_222_137 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__7214__A2 net72 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_116_32 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_92_69 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_203_2948 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5225__A1 _0782_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_155_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_231_693 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7760_ _1083_ _1080_ _1105_ _3834_ _3835_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_2
X_4972_ _1400_ _0580_ _1424_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_188_597 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_59_765 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_199_2896 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_25_96 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_148_439 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4823__I1 core_0.decode.i_instr_l\[9\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6711_ core_0.execute.rf.reg_outputs\[5\]\[3\] _3022_ _3016_ _3026_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3923_ _0539_ _0542_ _0544_ core_0.execute.rf.reg_outputs\[1\]\[14\] _0558_ vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_4
X_7691_ _1084_ _1080_ _1102_ _1065_ _1105_ _3791_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XTAP_TAPCELL_ROW_121_1969 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_73_212 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6642_ _2979_ core_0.ew_data\[9\] _2980_ net36 _2983_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_0_18_139 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_234 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_132_53 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_144_601 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_156_461 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_116_314 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_128_185 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_183_291 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6573_ _2927_ _0216_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6222__B _1114_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_132_807 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_144_667 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_172 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_312 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8312_ _0488_ clknet_leaf_76_i_clk net182 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_4
XFILLER_0_6_589 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5524_ _0797_ _0808_ _1952_ _1953_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_4
XFILLER_0_171_486 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_41_142 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_76_1426 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_8243_ _0419_ clknet_leaf_43_i_clk core_0.execute.sreg_irq_pc.o_d\[15\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_41_164 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5455_ core_0.execute.alu_mul_div.div_cur\[12\] _1803_ _1891_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__7150__A1 _1980_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4406_ net82 _1013_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_3
X_8174_ _0350_ clknet_leaf_129_i_clk core_0.execute.alu_mul_div.mul_res\[0\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5161__B1 _1437_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5386_ core_0.execute.alu_mul_div.div_cur\[3\] _1831_ _1773_ _1832_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_100_737 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_112_597 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_10_551 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_562 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7125_ _1994_ _3209_ _3330_ _3332_ _3333_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_4337_ core_0.fetch.prev_request_pc\[12\] _0954_ _0955_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_TAPCELL_ROW_243_3429 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7932__CLK clknet_leaf_24_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7453__A2 net75 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7056_ _3267_ _3268_ _3269_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_157_72 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4268_ _0723_ net61 _0885_ _0886_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_4
XFILLER_0_66_70 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6007_ net10 _2260_ _2264_ core_0.execute.sreg_irq_pc.o_d\[3\] _2397_ vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_198_317 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4199_ _0724_ net49 _0818_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_161_2439 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_97_816 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_96_304 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7205__A2 net202 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_241_479 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_87_1555 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4019__A2 _0578_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5216__A1 net97 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_222_671 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_96_337 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_194_523 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6964__A1 net217 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_82_91 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7958_ _0136_ clknet_leaf_17_i_clk core_0.execute.alu_mul_div.div_cur\[14\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_167_748 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_77_562 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_264 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6909_ net101 _3135_ _3139_ _3140_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_166_247 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7889_ _0080_ clknet_leaf_77_i_clk core_0.decode.i_instr_l\[14\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_49_286 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_77_595 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_92_521 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_804 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_65_746 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5519__A2 _0807_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_107_314 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_64_256 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_119_174 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_107_347 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6192__A2 _2257_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_45_470 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_64_289 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_21_763 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_107_369 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5527__I _0810_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4431__I _0733_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_632 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_134_155 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_45_492 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_122_317 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_134_177 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_172_2579 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_33_654 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_32_131 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_32_142 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_451 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_98_1684 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3950__A1 _0568_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_687 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7141__A1 _1225_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6358__I _1455_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_244_251 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5455__A1 core_0.execute.alu_mul_div.div_cur\[12\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_245_796 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_125_2014 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_204_126 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_99_142 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_232_457 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_99_164 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_213_671 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_198_862 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_29_863 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5758__A2 _1620_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6955__A1 _3175_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_158_737 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_185_534 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_107_1791 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_157_258 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_218_3133 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_55_212 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_95_381 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_543 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_172_217 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_60_1227 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_60_1238 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_43_407 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_102_34 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6183__A2 _2279_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_126_667 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_136_2143 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_126_689 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_153_475 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5930__A2 _1676_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_180_283 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_142 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_3_559 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_87_14 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5240_ _1625_ _1689_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_228_719 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_87_69 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7683__A2 _3778_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5694__A1 _1123_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4497__A2 _1062_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_229_3262 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_227_229 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_EDGE_ROW_18_Right_18 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
X_5171_ _1619_ _1620_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
X_4122_ core_0.execute.pc_high_out\[7\] _0732_ _0742_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_194_37 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_71_1367 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7435__A2 net87 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_208_454 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_235_251 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5446__A1 core_0.execute.alu_mul_div.div_cur\[10\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_235_273 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_147_2272 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_4053_ net98 _0578_ _0678_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xinput3 i_core_int_sreg[11] net3 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5997__A2 _0798_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7812_ core_0.dec_alu_flags_ie _1052_ _3872_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_188_372 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5749__A2 _2013_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6946__A1 _1713_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_47_702 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_562 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7743_ core_0.dec_jump_cond_code\[0\] _1062_ _3823_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4955_ _1400_ _0637_ _1412_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XPHY_EDGE_ROW_27_Right_27 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_93_329 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_148_247 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4421__A2 core_0.fetch.prev_request_pc\[0\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_176_578 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_129_450 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3906_ _0541_ _0542_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_8
X_7674_ _1133_ _1048_ _1104_ _3775_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_0_62_705 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_82_1496 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_117_623 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_163_228 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4886_ _1283_ _1356_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_46_256 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_191_559 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_62_716 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6625_ net26 _1148_ _2969_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_74_587 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_116_122 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_156_291 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_331 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_656 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_689 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_94_i_clk_I clknet_4_7__leaf_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6556_ net120 _2859_ _2189_ _2919_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_104_317 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_116_177 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5921__A2 _1592_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_42_451 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5507_ _1223_ _1939_ _1940_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__3932__A1 _0565_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6487_ _2834_ _2865_ _2866_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_14_186 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5134__B1 _1486_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_8226_ _0402_ clknet_leaf_8_i_clk core_0.execute.alu_flag_reg.o_d\[4\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_2
X_5438_ core_0.execute.alu_mul_div.div_cur\[10\] _1812_ _1841_ _1877_ vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__7674__A2 _1048_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_36_Right_36 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__5134__C2 _1435_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input51_I i_req_data[21] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_218_218 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8157_ _0333_ clknet_leaf_84_i_clk net88 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_4
X_5369_ _1816_ _1817_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
X_7108_ _3149_ _3315_ _3316_ _1501_ _3209_ _3317_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai32_1
X_8088_ _0264_ clknet_leaf_104_i_clk core_0.execute.rf.reg_outputs\[5\]\[11\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5437__A1 core_0.execute.alu_mul_div.div_cur\[9\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_242_722 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_199_615 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_242_733 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_226_284 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7039_ _3243_ _3252_ _3253_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA_output138_I net138 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5810__I _2201_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_242_755 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_198_136 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3999__A1 core_0.execute.rf.reg_outputs\[7\]\[8\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_202_619 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_93_90 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4660__A2 _1214_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_241_298 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_195_821 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8260__CLK clknet_leaf_36_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_195_832 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_45_Right_45 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_26_822 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_195_865 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_96_189 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_139_247 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7828__CLK clknet_leaf_53_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_37_212 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_77_381 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_167_578 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_46_1060 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_203_22 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_194_375 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7737__I0 net182 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_203_55 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_418 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_645 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_163_740 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_524 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_108_667 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4176__B2 _0771_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_123_626 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_213_3063 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_190_592 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_579 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_213_3074 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_150_434 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3923__A1 _0539_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_101 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7114__A1 _1227_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_54_Right_54 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_110_309 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_122_169 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5125__B1 _1443_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7665__A2 _1069_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_131_2084 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_185_2737 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7417__A2 net84 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_218_763 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_217_262 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_6_580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_109_1820 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_233_766 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_205_457 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__7140__C _1225_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_63_Right_63 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__6037__B _1061_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4651__A2 net192 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_200_2907 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_200_2918 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6928__A1 _1227_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_185_320 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_196_2866 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4403__A2 _0950_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_96_690 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_158_578 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_113_22 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4740_ core_0.fetch.out_buffer_data_instr\[24\] net54 _1246_ _1271_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_7_106 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_200_195 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_29_768 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_863 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_145_228 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_185_397 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_138_280 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_clkbuf_leaf_116_i_clk_I clknet_4_4__leaf_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4671_ _1226_ _1227_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_113_88 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_43_226 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_83_395 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7353__A1 _1217_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_154_762 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_118_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_126_464 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6410_ _1379_ core_0.execute.sreg_irq_pc.o_d\[12\] _2791_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_189_26 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_141_401 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_153_261 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7390_ _1357_ net79 _3553_ _3555_ _3556_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__5903__A2 _2133_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_72_Right_72 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
X_6341_ _2663_ _2723_ _2724_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_12_613 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__3914__A1 _0539_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7105__A1 _2778_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_98_79 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_141_467 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_367 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_112 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_141_489 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5116__B1 _1486_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6272_ _2576_ _2655_ _2656_ _0186_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__5116__C2 _1435_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_149_2301 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_8011_ _0188_ clknet_leaf_53_i_clk core_0.ew_data\[10\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_2
XANTENNA__5667__A1 _1803_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5223_ _0771_ _0768_ _0776_ core_0.execute.rf.reg_outputs\[6\]\[2\] _1672_ vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_0_110_865 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_209_730 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5831__S _2219_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5154_ _1596_ _1603_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XANTENNA__7408__A2 _3542_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5419__A1 _1747_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_47_72 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_4105_ _0724_ _0725_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_5085_ core_0.execute.rf.reg_outputs\[7\]\[14\] net233 _1443_ core_0.execute.rf.reg_outputs\[3\]\[14\]
+ _1534_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XPHY_EDGE_ROW_81_Right_81 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__6092__A1 core_0.execute.alu_mul_div.div_cur\[4\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_223_243 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4036_ _0515_ core_0.dec_r_reg_sel\[1\] _0525_ _0662_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_4
XANTENNA__4642__A2 net192 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_196_629 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_84_1525 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6919__A1 net91 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_149_556 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7592__A1 core_0.execute.pc_high_buff_out\[5\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_192_802 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5987_ _2300_ _2374_ _2377_ _1624_ _1480_ _2378_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_0_93_126 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_212 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_109_409 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_234 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_176_375 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7726_ _3814_ _0482_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4938_ _1381_ _1400_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA__7719__I0 net188 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_176_397 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_164_559 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_7_640 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4869_ _0837_ _1348_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_7657_ _3761_ _3762_ _3763_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_62_535 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_90_Right_90 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_7_673 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_855 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_105_615 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4158__A1 _0768_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6608_ _2929_ _2953_ _2954_ _2955_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_2
XTAP_TAPCELL_ROW_31_880 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_7588_ core_0.execute.pc_high_out\[4\] _3672_ _3708_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_172_592 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_659 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6539_ _2910_ _0199_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7506__B _3516_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_70_590 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_95_1654 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_113_692 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5658__A1 _1754_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_8209_ _0385_ clknet_leaf_31_i_clk net81 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_4
Xoutput170 net170 o_req_addr[3] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
Xoutput181 net181 sr_bus_addr[12] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
Xoutput192 net192 sr_bus_addr[8] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA__4881__A2 _1321_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_215_755 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6083__A1 _1137_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_3_550 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_180_2667 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_187_607 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_180_2678 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_214_276 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_187_629 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4156__I core_0.dec_l_reg_sel\[0\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4633__A2 core_0.execute.alu_flag_reg.o_d\[3\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_134 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6572__S _2201_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_161_Left_408 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_230_758 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_39_980 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_97_465 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_167 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_318 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_168_865 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_38_521 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_183_813 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_104_1761 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_167_364 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4397__A1 _0959_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_195_684 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_127_206 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_194_172 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_183_835 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_863 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_705 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4936__A3 _1390_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_26_716 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_362 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_26_749 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_81_833 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6138__A2 _2524_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7335__A1 net194 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_230_53 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_259 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_80_354 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_133_2113 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5897__A1 _1456_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_80_387 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_170_Left_417 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_150_242 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_151_776 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_111_629 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_123_489 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7638__A2 _3729_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_115_1890 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_226_3221 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_225_508 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4321__A1 _0935_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_206_700 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_218_571 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_206_733 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4872__A2 _1341_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_42_i_clk_I clknet_4_9__leaf_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_233_541 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_206_755 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_144_2242 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_88_410 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7810__A2 _1053_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4066__I net212 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_205_298 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_187_Right_187 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
X_5910_ _1531_ _1491_ _2302_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_221_758 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6890_ core_0.ew_reg_ie\[0\] _2934_ _3128_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_76_605 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_177_139 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5841_ _2232_ _2234_ _2235_ _0175_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__7574__A1 core_0.execute.pc_high_out\[3\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7377__I _3540_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_174_802 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_235_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_185_150 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_75_137 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_174_813 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4388__A1 _0843_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_185_161 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_33_74 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_8_415 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_66_1299 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_75_159 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5772_ _2172_ _2056_ _2173_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_TAPCELL_ROW_237_3361 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_185_183 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_185_194 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_660 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_107 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_173_334 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_671 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7511_ _3649_ _3650_ _0431_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_16_204 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_8_459 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4723_ _1261_ _1237_ _1262_ _0031_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_44_524 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_127_751 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6129__A2 _1624_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7326__A1 _2565_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_72_855 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_83_192 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7442_ _0615_ _3546_ _3545_ _3598_ _3599_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai211_1
XTAP_TAPCELL_ROW_155_2371 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_4654_ net106 _1212_ _1213_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_71_365 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_154_592 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_632 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_140_86 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput50 i_req_data[20] net50 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput61 i_req_data[30] net61 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_7373_ _1209_ _2577_ _3540_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_4
X_4585_ _1157_ net151 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_3_142 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_114_478 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_12_432 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_114_489 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_142_798 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6324_ _2123_ _2096_ _2707_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_12_454 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_141_286 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_465 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6255_ _1061_ _2037_ _2637_ _1109_ _2639_ _2640_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_0_0_860 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6301__A2 core_0.execute.alu_mul_div.mul_res\[9\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
X_5206_ _0771_ _0773_ core_0.execute.rf.reg_outputs\[5\]\[3\] _1655_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_0_110_695 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6186_ _2544_ _2572_ core_0.dec_mem_access _2573_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_42_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_90_1595 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4863__A2 _1341_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5137_ core_0.execute.rf.reg_outputs\[2\]\[8\] _1438_ _1586_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_165_50 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6065__A1 _1378_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_165_72 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5068_ _1513_ _1514_ _1515_ _1516_ _1517_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and4_1
XANTENNA_input14_I i_core_int_sreg[7] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5812__A1 _2202_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_169_629 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4019_ net101 _0578_ _0647_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_212_769 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_154_Right_154 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__4091__A3 _0549_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_94_402 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_36_950 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_66_104 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_67_627 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_177_640 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7565__A1 _3673_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6368__A2 _2332_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_0_Right_0 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__6191__I _2264_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_94_457 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_48_863 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_80 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_191_120 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_43_1030 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_47_373 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_164_345 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_191_142 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7709_ _1085_ _1098_ _3763_ _3805_ _3806_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and4_1
XANTENNA__7317__A1 _3409_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_62_321 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_74_181 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_164_378 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_35_557 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_652 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_118_784 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_412 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_492 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_22_207 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_50_516 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_376 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_132_220 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_50_527 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_62_387 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_22_229 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_200_34 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6140__B core_0.dec_mem_access vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_160_562 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_210_3033 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_105_478 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_output82_I net82 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_30_251 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_219_302 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_101_640 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_207_508 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_101_695 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_207_519 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_246_176 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4854__A2 _1307_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_234_349 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_243_850 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_199_220 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_54_18 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_89_207 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6056__B2 core_0.execute.alu_flag_reg.o_d\[4\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_230_511 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_203_736 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_202_213 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_221_3162 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4815__S _1305_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_98_763 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_230_544 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_187_437 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_159_128 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_121_Right_121 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__4082__A3 _0527_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_202_279 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3939__B _0520_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_211_780 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6359__A2 _1620_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7556__A1 core_0.execute.pc_high_out\[0\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_193_2825 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_183_632 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_195_492 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_183_643 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_129 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7308__A1 net77 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_53_310 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_183_676 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_14_677 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_115_209 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_155_389 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_183_698 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4790__A1 _1290_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_123_220 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_80_173 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_110_34 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_232_3291 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_151_562 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_110_45 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_124_798 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4370_ core_0.fetch.prev_request_pc\[11\] _0953_ _0984_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__5098__A2 _1484_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6040_ _1665_ _2420_ _1999_ _2424_ _2429_ _2430_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai221_4
XANTENNA__6295__B2 _1754_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input6_I i_core_int_sreg[14] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_185_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_206_563 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6598__A2 _2941_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7991_ _0168_ clknet_leaf_20_i_clk net159 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_2
XTAP_TAPCELL_ROW_206_2979 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_68_1328 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7795__B2 _1037_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_178_426 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6942_ _3158_ _3159_ _3161_ _3162_ _1223_ _3163_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XANTENNA__5270__A2 _1548_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_159_640 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_48_104 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_193_418 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7547__A1 _3637_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6873_ core_0.execute.rf.reg_outputs\[1\]\[8\] _3114_ _3112_ _3119_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_9_702 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_49_649 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_88_295 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_119_526 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_157_2400 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_5824_ _2195_ _2203_ _2207_ _2215_ _2221_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor4_2
XFILLER_0_151_30 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5022__A2 _1469_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_9_768 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5755_ _1515_ _1516_ _2156_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_173_142 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_44_321 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_84_490 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6770__A2 _3043_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_115_710 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4706_ core_0.fetch.out_buffer_data_instr\[10\] net39 _1246_ _1251_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_44_354 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_803 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4781__B2 net175 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5686_ _1711_ _1549_ _1992_ _2086_ _2087_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai22_2
XFILLER_0_32_516 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_387 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_32_527 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_440 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_115_765 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_79_1457 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_4637_ net186 _1196_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__inv_2
X_7425_ core_0.execute.sreg_irq_pc.o_d\[7\] _3543_ _3584_ _3585_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__4399__C _0877_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_102_415 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4533__A1 _1056_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_4_495 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_229_600 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4568_ _1147_ _1148_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
X_7356_ _2646_ _2684_ _3524_ _3525_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor3_1
XTAP_TAPCELL_ROW_92_1613 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6895__B _3124_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_130_768 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6307_ _2663_ _2665_ _2690_ _2360_ _2691_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_7287_ _3384_ _3464_ _3465_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_229_655 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4499_ _1038_ _1039_ _1069_ _1090_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_4
XANTENNA__6286__A1 _2294_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5089__A2 _1435_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_223_Right_223 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
X_6238_ _2616_ _2622_ _2623_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4836__A2 _1307_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6169_ _1761_ _1613_ _1686_ _2556_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_176_93 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6038__B2 _1831_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_197_702 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7786__A1 _1136_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output120_I net120 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_224_393 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_169_426 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_67_413 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_79_273 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_212_588 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_39_126 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7538__A1 _3663_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4434__I _0742_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_94_243 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_149_172 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_177_481 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_101_1720 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_177_492 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6210__A1 net223 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_48_671 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_107 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5013__A2 _1382_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_164_142 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_192_462 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_165_687 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_855 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6761__A2 _3042_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_192_484 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_663 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_11_647 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7010__I0 _2001_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_211_66 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_836 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_51_858 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_133_562 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_16_590 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5265__I core_0.decode.oc_alu_mode\[12\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7710__A1 _2242_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7710__B2 _3806_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4524__A1 _1065_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_160_381 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_239_419 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_105_297 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6277__A1 _1379_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_208_828 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_112_1860 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_101_492 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_235_636 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_235_647 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_128_2045 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6029__A1 _1480_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_216_861 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_243_680 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_141_2201 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7777__A1 _1136_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_243_691 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_231_842 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_187_212 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_19_736 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_5_i_clk clknet_4_2__leaf_i_clk clknet_leaf_5_i_clk vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_203_566 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5252__A2 _1527_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_81_49 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_86_744 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_175_418 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_457 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_156_610 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_85_276 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5004__A2 core_0.decode.oc_alu_mode\[11\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_63_1269 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_234_3320 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_155_142 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_170 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_26_332 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6752__A2 _3049_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_183_473 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_170_101 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_139_2185 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_5540_ core_0.execute.mem_stage_pc\[4\] _1957_ _1964_ _1965_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_143_348 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_170_123 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_41_302 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_5_248 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_30_53 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_527 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_26_398 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_112_702 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5471_ _1375_ _1903_ _1904_ _1822_ _1905_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XTAP_TAPCELL_ROW_152_2341 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5175__I _1531_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_100_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_30_86 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_124_584 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4422_ _0959_ _1025_ _1026_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__4515__A1 _1101_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7210_ _0810_ _1734_ _3397_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__5108__C _1460_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_8190_ _0366_ clknet_leaf_18_i_clk core_0.execute.next_ready_delayed vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_151_392 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_443 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_7141_ _1225_ _3297_ _3346_ _3347_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_4353_ _0965_ _0970_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_111_278 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_238_452 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_487 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_226_603 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6268__B2 _2356_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_62 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7072_ _1224_ _1914_ _3283_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA_clkbuf_4_7__f_i_clk_I clknet_3_3_0_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4284_ core_0.fetch.prev_request_pc\[7\] _0833_ _0901_ core_0.fetch.prev_request_pc\[6\]
+ _0902_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_TAPCELL_ROW_74_1398 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_10_799 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4818__A2 core_0.fetch.submitable vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6023_ _1624_ _2313_ _2413_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5124__B _0778_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5491__A2 net219 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_241_628 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7768__A1 core_0.decode.i_instr_l\[8\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_222_831 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_163_2470 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_55_83 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_178_212 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7974_ _0151_ clknet_leaf_56_i_clk core_0.execute.mem_stage_pc\[9\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_178_234 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_221_352 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6440__A1 _2812_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_179_768 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_76_210 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6925_ net94 _3128_ _3139_ _3148_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__6991__A2 _1819_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_178_289 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_193_226 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_147_621 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_76_254 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_92_714 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6856_ _2940_ _3107_ _3109_ _0317_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_147_632 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_159_492 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_36_107 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_92_725 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5807_ core_0.execute.rf.reg_outputs\[1\]\[2\] _1615_ _2206_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_119_367 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_92_758 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_162_602 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3999_ core_0.execute.rf.reg_outputs\[7\]\[8\] _0530_ _0628_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_18_855 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6787_ _2956_ _3064_ _3069_ _0288_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__6743__A2 _3042_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_174_473 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_147_698 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_652 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_161_112 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_174_495 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_45_674 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5738_ _1698_ _1722_ _2138_ _2139_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_0_161_123 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_17_376 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_836 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_32_313 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_493 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_858 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_32_335 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_115_562 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5669_ _1752_ _1568_ _2070_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_60_655 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8217__CLK clknet_leaf_36_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4506__A1 _1043_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7408_ core_0.execute.sreg_irq_pc.o_d\[4\] _3542_ _3516_ _3571_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_13_582 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output168_I net168 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7339_ _2183_ _3502_ _3511_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6259__A1 _1059_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_229_463 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_229_485 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_229_496 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4809__A2 core_0.fetch.submitable vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4429__I _0736_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_244_466 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7759__A1 _1045_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_89_i_clk_I clknet_4_6__leaf_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_213_842 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_99_368 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_169_212 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6431__A1 _2113_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_240_683 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_16_706 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_240_694 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_157_418 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_206_99 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_200_536 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_197_598 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6982__A2 _1931_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6580__S _2201_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_177_2639 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4993__A1 _0782_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_82_202 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_184_259 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_298 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6195__B1 _2534_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_83_758 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6734__A2 _3022_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_165_484 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_125_326 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4596__I1 core_0.ew_data\[12\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_222_98 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_63_460 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_125_348 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_708 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_23_324 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5209__B _0769_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_51_644 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_51_655 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6498__A1 _2287_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_133_392 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_121_554 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7424__B _3545_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_39_Left_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_188_2768 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_208_603 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_76_49 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_235_422 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6670__A1 _2946_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5473__A2 _1812_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_188_521 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_240_3390 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_203_2949 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_203_352 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4028__A3 _0543_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5225__A2 _0768_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_48_Left_295 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
X_4971_ _1419_ _1423_ _0118_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_230_171 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_59_755 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_129_610 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_148_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_199_2897 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6710_ _2951_ _3021_ _3025_ _0255_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_19_608 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3922_ _0554_ _0528_ _0555_ _0556_ _0557_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai211_4
XFILLER_0_129_632 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_58_265 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7690_ _1084_ _1092_ _1119_ _1140_ _3790_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_18_107 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_58_276 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_121_1959 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_184_760 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6641_ _2936_ _2981_ _2982_ _0229_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__6725__A2 _3027_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_117_838 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_rebuffer4_I net223 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_171_410 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_144_635 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4802__I _1305_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6572_ core_0.dec_rf_ie\[6\] core_0.ew_reg_ie\[6\] _2201_ _2927_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_41_96 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_15_836 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8311_ _0487_ clknet_leaf_68_i_clk net181 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_4
XFILLER_0_54_493 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5523_ core_0.decode.i_flush _1951_ _1952_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_15_858 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_76_1427 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_42_677 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5454_ _1889_ _1890_ _0134_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_8242_ _0418_ clknet_leaf_43_i_clk core_0.execute.sreg_irq_pc.o_d\[14\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_42_688 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_379 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_30_839 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7150__A2 _0807_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_140_863 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4405_ _1008_ _0966_ _1011_ _1012_ _0877_ net172 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XANTENNA__5161__A1 core_0.execute.rf.reg_outputs\[4\]\[6\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5161__B2 core_0.execute.rf.reg_outputs\[2\]\[6\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
X_8173_ _0349_ clknet_leaf_0_i_clk core_0.execute.alu_mul_div.cbit\[0\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_4
X_5385_ _1765_ _1831_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_239_761 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_239_772 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4336_ core_0.fetch.prev_request_pc\[11\] _0953_ _0954_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
X_7124_ _3175_ _3331_ _3332_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xclkbuf_leaf_106_i_clk clknet_4_5__leaf_i_clk clknet_leaf_106_i_clk vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_10_574 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_226_433 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7055_ _2648_ _3265_ _3268_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4267_ _0723_ _0845_ _0885_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6006_ core_0.execute.sreg_long_ptr_en _1385_ _2250_ core_0.execute.sreg_irq_flags.o_d\[3\]
+ _2396_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__6661__B2 net27 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_214_639 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4198_ core_0.fetch.out_buffer_data_instr\[1\] _0817_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__inv_1
XANTENNA_clkbuf_leaf_90_i_clk_I clknet_4_6__leaf_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_241_458 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_87_1556 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6413__A1 _2244_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5216__A2 _1492_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_173_72 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7957_ _0135_ clknet_leaf_5_i_clk core_0.execute.alu_mul_div.div_cur\[13\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__6964__A2 _1650_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6908_ _0722_ _3139_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA__4975__A1 _1400_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7888_ _0079_ clknet_leaf_83_i_clk core_0.decode.i_instr_l\[13\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_194_579 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_119_142 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_181_207 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6839_ _2983_ _3086_ _3099_ _0310_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_147_462 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6413__B core_0.dec_mem_access vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6716__A2 _3027_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_134_101 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_175_793 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_181_229 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_92_577 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_92_588 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_162 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_780 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_21_764 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_33_644 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_162_476 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_98_1685 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_33_699 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7244__B net84 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_130_362 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_229_282 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_217_422 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6101__B1 _2264_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_70_i_clk clknet_4_15__leaf_i_clk clknet_leaf_70_i_clk vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__5455__A2 _1803_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6652__B2 net24 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_125_2015 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_198_830 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_88_839 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5207__A2 _1605_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_29_864 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_213_683 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_87_338 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_197_384 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_185_524 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_leaf_85_i_clk clknet_4_12__leaf_i_clk clknet_leaf_85_i_clk vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__4966__A1 _1400_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_107_1792 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4823__S _1305_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_4_13__f_i_clk_I clknet_3_6_0_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_83_500 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_218_3123 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_173_708 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_218_3134 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_28_427 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6707__A2 _3022_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_60_1228 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_55_279 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_126_657 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_70_216 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_136_2144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_24_633 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4194__A2 _0812_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_140_104 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_141_627 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_66 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_140_115 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_12_839 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_24_699 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_140_159 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_122_863 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7154__B _3357_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_23_i_clk clknet_4_8__leaf_i_clk clknet_leaf_23_i_clk vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__5694__A2 _1620_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5170_ net101 _1618_ _1446_ _1619_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_229_3263 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6993__B _3189_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_236_731 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4121_ core_0.execute.prev_pc_high\[2\] _0735_ _0736_ core_0.execute.prev_pc_high\[1\]
+ _0740_ _0741_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai221_4
XFILLER_0_208_444 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_clkbuf_leaf_112_i_clk_I clknet_4_4__leaf_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_71_1368 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_38_i_clk clknet_4_11__leaf_i_clk clknet_leaf_38_i_clk vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_208_477 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5446__A2 _1814_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4052_ _0673_ _0674_ _0675_ _0676_ _0677_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and4_1
XTAP_TAPCELL_ROW_147_2273 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
Xinput4 i_core_int_sreg[12] net4 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_235_296 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_223_458 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_63 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_56_Left_303 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_78_305 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_96 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7199__A2 _2334_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7811_ _1034_ _3870_ _3871_ _0510_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__6946__A2 _1926_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_188_384 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_176_524 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4957__A1 _1301_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8062__CLK clknet_leaf_109_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7742_ _3822_ _0490_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4954_ _1301_ _1411_ _0113_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_19_438 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3905_ _0540_ _0541_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_46_235 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7673_ _1034_ _3773_ _3774_ _0469_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4885_ _1279_ _1285_ _0883_ _0100_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_1
XTAP_TAPCELL_ROW_82_1497 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_191_549 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6624_ _2936_ _2967_ _2968_ _0226_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_46_279 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_37_i_clk_I clknet_4_11__leaf_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_482 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_65_Left_312 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__5382__A1 core_0.execute.alu_mul_div.div_cur\[1\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_171_251 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6555_ _2918_ _0207_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_15_644 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_249 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_6_387 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5506_ _1367_ _1928_ _1938_ _1939_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA__7659__B1 _1064_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3932__A2 _0541_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6486_ _1380_ _2863_ _2864_ _2865_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_42_485 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5134__A1 core_0.execute.rf.reg_outputs\[1\]\[9\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
X_8225_ _0401_ clknet_leaf_12_i_clk core_0.execute.alu_flag_reg.o_d\[3\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5437_ core_0.execute.alu_mul_div.div_cur\[9\] _1814_ _1817_ _1875_ _1876_ vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_246_506 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_112_384 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_218_208 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_593 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_100_535 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_112_395 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6882__A1 _2990_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5368_ _1232_ _1815_ core_0.execute.alu_mul_div.comp _0801_ _1816_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__oai211_4
X_8156_ _0332_ clknet_leaf_79_i_clk core_0.execute.rf.reg_outputs\[1\]\[15\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_2
XANTENNA_input44_I i_req_data[15] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_77_81 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_100_568 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7107_ _3305_ _3307_ _3314_ _3316_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and3_1
X_4319_ net39 core_0.fetch.out_buffer_data_instr\[10\] _0725_ _0937_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_8087_ _0263_ clknet_leaf_100_i_clk core_0.execute.rf.reg_outputs\[5\]\[10\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5299_ _1746_ _1747_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__6634__A1 _2930_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5437__A2 _1814_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_227_797 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_7038_ _3251_ _3252_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XPHY_EDGE_ROW_74_Left_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_184_82 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_241_244 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3999__A2 _0530_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_241_255 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_201_119 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_26_823 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_139_204 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_output200_I net200 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_167_535 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_195_855 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4948__A1 _1301_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_77_360 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_194_343 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_46_1061 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_93_842 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_108_602 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_37_246 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_65_555 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5538__I _0722_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_182_527 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7737__I1 core_0.decode.i_imm_pass\[13\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_37_257 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_65_566 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_37_279 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_83_Left_330 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_107_134 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_108_657 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_163_752 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_46_791 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_135_465 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5373__A1 _1374_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_122_104 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_135_487 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_213_3064 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3923__A2 _0542_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_122_137 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__7114__A2 _1501_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_104_863 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_496 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_150_479 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_131_693 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_209_219 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_131_2085 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_185_2727 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_185_2738 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_168_Right_168 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__6625__A1 net26 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_205_414 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_6_581 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_109_1821 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5222__B net219 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_232_244 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_232_255 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_87_102 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_87_113 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_88_647 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_200_2908 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_87_135 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_88_669 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6928__A2 _1841_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_158_524 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7050__A1 _1224_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4939__A1 _1400_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5876__C core_0.dec_sreg_irt vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_200_141 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_158_557 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_196_2867 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_8_619 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_113_34 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_341 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_7_129 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_56_566 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_268 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_16_419 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4670_ core_0.execute.alu_mul_div.cbit\[0\] _1226_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__inv_4
XANTENNA__7922__CLK clknet_leaf_8_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_43_238 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_141_413 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_452 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6340_ _1379_ core_0.execute.sreg_irq_pc.o_d\[10\] _2722_ _2723_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_3_346 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_783 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7105__A2 _3313_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_51_282 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6271_ core_0.ew_data\[8\] _2486_ _2656_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_12_658 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8010_ _0187_ clknet_leaf_55_i_clk core_0.ew_data\[9\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_2
X_5222_ core_0.execute.rf.reg_outputs\[1\]\[2\] _1615_ net219 _1671_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__5667__A2 _1501_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_149_2302 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_110_855 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_11_179 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_209_742 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5153_ _1560_ _1597_ _1601_ _1602_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_243_509 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_135_Right_135 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_208_241 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_236_561 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4104_ _0723_ _0724_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_5084_ core_0.execute.rf.reg_outputs\[2\]\[14\] _1438_ _1533_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5132__B _0779_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4035_ _0515_ _0540_ _0518_ _0661_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_4
XANTENNA__6092__A2 _1432_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_223_255 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_211_417 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4642__A3 _1199_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_189_671 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_2_75 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_84_1515 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_84_1526 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6919__A2 _3135_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7041__A1 _3149_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_63_72 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_78_157 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_94_617 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5986_ _2300_ _2376_ _2377_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_137_708 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7592__A2 _3682_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_75_842 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_93_138 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7059__B _3189_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7725_ net191 core_0.decode.i_imm_pass\[7\] _1946_ _3814_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_164_527 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_4937_ _1397_ _1399_ _1284_ _0108_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_176_387 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_246 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_191_335 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7656_ _1074_ _1080_ _1037_ _3762_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4868_ _1347_ _0091_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6607_ net30 _1149_ _2954_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4158__A2 _0776_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_249 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_31_881 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_105_627 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7587_ net204 _3675_ _3706_ _3707_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_144_284 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_160_733 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4799_ _1146_ _1237_ _1304_ _0065_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_43_772 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_132_446 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6538_ net126 _2526_ _2906_ _2910_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_15_485 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_70_580 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_95_1655 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5107__A1 _1466_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6469_ _1137_ _2179_ _2846_ _1109_ _2847_ _2848_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_0_179_93 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8208_ _0384_ clknet_leaf_32_i_clk net80 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_4
XANTENNA__5658__A2 _1585_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_100_321 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xoutput160 net160 o_req_active vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_246_336 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput171 net171 o_req_addr[4] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_11_680 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput182 net182 sr_bus_addr[13] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
Xoutput193 net193 sr_bus_addr[9] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
X_8139_ _0315_ clknet_leaf_97_i_clk core_0.execute.rf.reg_outputs\[2\]\[14\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_100_387 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XPHY_EDGE_ROW_102_Right_102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__6607__A1 net30 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_215_723 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_242_520 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_242_542 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7280__A1 _3409_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_215_767 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6083__A2 _1683_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_214_244 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_3_551 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_180_2668 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_97_422 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_230_737 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_242_597 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_186_107 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_186_118 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_39_981 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_69_146 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7032__A1 _1226_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_85_617 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_168_855 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5696__C _2092_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_210_450 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_78_691 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_104_1762 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5594__A1 _1702_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_182_302 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_194_184 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_65_352 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_182_335 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_588 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_728 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_80_311 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7335__A2 _3495_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_108_465 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_182_379 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_80_333 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5346__A1 core_0.execute.alu_mul_div.div_cur\[10\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_123_402 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_136_785 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_133_2103 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_237_Right_237 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_133_2114 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_40_208 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_33_282 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_422 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7099__A1 _1230_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_110_107 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_150_287 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_103_181 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_238_859 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_115_1891 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_226_3222 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4321__A2 _0936_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_84_49 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_45 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7271__A1 net87 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_205_233 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4347__I net77 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_144_2243 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4085__A1 _0567_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_205_266 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_221_726 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_205_277 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5821__A2 _1615_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4624__A3 core_0.execute.alu_flag_reg.o_d\[0\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_220_225 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7023__A1 _1372_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5840_ net137 _2209_ _2235_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_57_842 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4388__A2 _0947_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_186_685 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_173_302 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_237_3351 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_185_173 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5771_ _2170_ _1568_ _2172_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_130_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_146_527 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_158_387 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_237_3362 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_228_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_17_706 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7510_ core_0.execute.sreg_scratch.o_d\[5\] _3641_ _1217_ _3650_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_44_514 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4722_ net44 _1253_ _1262_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_173_346 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_84_683 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7326__A2 _2606_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_83_171 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_322 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_161_519 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7441_ _3563_ net73 _3553_ _3597_ _3598_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai211_2
XANTENNA__5337__A1 core_0.execute.alu_mul_div.div_cur\[9\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6385__I0 _2122_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4653_ core_0.execute.sreg_jtr_buff.o_d\[0\] _1208_ _1211_ _1172_ _0731_ _1212_ vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_0_4_622 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_155_2372 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_204_Right_204 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
Xinput40 i_req_data[11] net40 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_25_772 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_3_121 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput51 i_req_data[21] net51 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_140_98 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7372_ _3538_ _3539_ _1395_ _0403_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
Xinput62 i_req_data[31] net62 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_4584_ core_0.ew_data\[6\] net157 _1157_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_142_777 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6323_ _2121_ _2706_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA_clkbuf_0_i_clk_I i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_797 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6254_ _1592_ _1455_ _2638_ _2639_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_12_499 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_110_663 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_228_347 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5205_ _1644_ _1653_ _1654_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_149_96 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_216_509 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_209_550 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6185_ _2360_ _2571_ _2572_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_209_572 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_90_1596 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_5136_ _1579_ _1584_ _1585_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_0_209_594 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_224_531 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_35_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7262__A1 _2652_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5067_ _0652_ _0657_ _0659_ _1459_ _1516_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai31_4
XFILLER_0_212_715 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_212_737 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_4018_ _0642_ _0643_ _0644_ _0645_ _0646_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_4
XTAP_TAPCELL_ROW_0_510 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4615__A3 core_0.execute.alu_flag_reg.o_d\[2\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_168_107 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_196_449 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_36_940 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_149_343 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_94_436 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_181_72 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_137_516 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_176_162 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5576__A1 _1051_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5969_ _2356_ _2360_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_47_352 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_43_1031 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_165_858 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_192_655 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_47_363 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_118_741 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7708_ _1039_ _1084_ _1103_ _3805_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_117_240 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7517__B _3651_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_62_333 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_74_193 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5328__A1 core_0.execute.alu_mul_div.div_cur\[4\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
X_7639_ net227 _3733_ _3749_ _3750_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_62_344 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_191_187 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_145_593 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_133_766 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4000__A1 _0565_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_90 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_210_3034 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_43_591 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_282 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_120_416 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_120_438 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6828__A1 _2961_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_8_610 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_246_122 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output75_I net75 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_101_663 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5500__A1 _1908_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_3_2_0_i_clk_I clknet_0_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_54_1160 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_246_166 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_234_317 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_209_66 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_209_88 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_209_99 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7253__A1 _1742_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6056__A2 _1385_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_243_862 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_199_232 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_242_350 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_242_361 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_221_3163 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_187_416 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_98_753 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_202_247 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_11_Left_258 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__7556__A2 _3673_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_842 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_57_138 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5567__A1 _1419_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_128_527 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_155_302 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_210_291 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_193_2826 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_66_683 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7308__A2 net76 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_26_536 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_14_678 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_124_711 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6516__B1 _2534_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_136_582 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_170_327 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_151_530 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_117_1920 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_123_243 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_232_3292 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_22_731 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_20_Left_267 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_110_79 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6819__A1 _2940_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_104_490 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_238_645 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_237_133 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_226_807 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_238_667 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6295__A2 _1455_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_218_380 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7244__A1 net83 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6047__A2 _2436_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_178_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4058__A1 _0533_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7990_ _0167_ clknet_leaf_19_i_clk core_0.execute.prev_sys vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_233_383 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_68_1329 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6941_ _1231_ _1758_ _1761_ _1926_ _1367_ _3162_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_0_221_556 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_221_567 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_617 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_76_403 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5410__B _1817_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_44_85 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6872_ _2977_ _3107_ _3118_ _0324_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_159_663 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_202_781 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_33_910 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5558__A1 _0977_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5823_ _2212_ _2215_ _2220_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_TAPCELL_ROW_157_2401 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_147_836 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_29_341 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_650 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_147_858 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_45_812 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_17_503 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5754_ _2017_ _1619_ _2155_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_17_536 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_162_839 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4705_ _1250_ _0025_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4781__A2 _1285_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_115_722 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_127_582 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_72_664 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5685_ _1990_ _1991_ _1996_ _2085_ _2086_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_44_366 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_114_232 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7424_ _0648_ _3544_ _3545_ _3583_ _3584_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_4636_ core_0.dec_sreg_irt _1195_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_4
XFILLER_0_71_185 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_79_1458 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_4_463 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5730__A1 _1689_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7355_ _2821_ _2777_ _3524_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__4533__A2 _1068_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4567_ core_0.ew_addr\[0\] core_0.ew_mem_width _1147_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_8_85 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_92_1614 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6306_ _2687_ _2688_ _2689_ _2690_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_4
XFILLER_0_229_634 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_229_645 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7286_ net74 _3462_ _3463_ _1735_ _3464_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_40_594 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4498_ _1063_ _0514_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XTAP_TAPCELL_ROW_168_2530 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6237_ _1379_ core_0.execute.sreg_irq_pc.o_d\[8\] _2621_ _2622_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__5371__I _1554_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_228_177 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_216_317 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_216_339 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6168_ _1137_ _2156_ _1456_ _2555_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_85_81 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_243_158 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5119_ _1567_ _1568_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
X_6099_ _2202_ _2485_ _2487_ _0182_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_212_534 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_240_854 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_output113_I net113 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5320__B core_0.execute.alu_mul_div.div_cur\[1\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_197_769 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_192_93 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_94_211 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_138_803 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_436 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6135__C _0799_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_184_419 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_39_138 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_149_162 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_801 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_101_1721 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6210__A2 _2414_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_137_346 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_620 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_125_508 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_153_817 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_192_474 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_106_711 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_153_839 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_165_699 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_62_130 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_11_648 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_118_593 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_180_647 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_517 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4450__I core_0.decode.i_instr_l\[2\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7010__I1 _1665_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_62_163 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_23_528 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_133_541 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_85_i_clk_I clknet_4_12__leaf_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_23_539 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_325 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_211_89 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_133_574 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7710__A2 _1134_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_239_409 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4524__A2 _1039_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_160_371 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_219_122 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7474__A1 _3581_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_112_1861 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_235_626 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_65_18 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_128_2046 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7226__A1 _3384_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6029__A2 _2411_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_215_361 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_141_2202 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_236_86 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_187_202 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5788__A1 _1051_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_19_737 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5230__B _1624_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_86_734 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7529__A2 _3646_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4460__A1 _1034_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_129_836 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_105_68 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_156_622 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_406 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_123_1990 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_129_858 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_183_441 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_234_3321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_128_357 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_183_452 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_480 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_128_368 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7157__B _3357_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_54_642 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_144_839 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_5_216 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_139_2175 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_42_804 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_54_664 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_121_34 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_139_2186 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_109_593 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_152_2331 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_5470_ _1374_ _1899_ _1904_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_121_89 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_152_2342 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7701__A2 _3766_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_347 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4421_ core_0.fetch.prev_request_pc\[1\] core_0.fetch.prev_request_pc\[0\] _1025_
+ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__5712__A1 _1600_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1_422 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_112_758 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_112_769 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7140_ _1364_ _3322_ _3345_ _1225_ _3346_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_0_111_246 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4352_ _0957_ _0968_ _0969_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_22_594 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_10_734 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7465__A1 _3563_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4283_ _0838_ _0901_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_7071_ _3282_ _0359_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_74_1399 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_245_3450 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6022_ _1682_ _1683_ _2412_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_0_226_659 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7217__A1 _1736_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7620__B _1216_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4736__S _1246_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7768__A2 core_0.decode.i_instr_l\[7\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_163_2471 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_7973_ _0150_ clknet_leaf_38_i_clk core_0.execute.mem_stage_pc\[8\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_233_191 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4535__I core_0.decode.oc_alu_mode\[11\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6924_ _2994_ _3130_ _3147_ _0347_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__4451__A1 core_0.decode.i_instr_l\[3\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_76_244 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6855_ core_0.execute.rf.reg_outputs\[1\]\[0\] _3108_ _3098_ _3109_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_18_801 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_147_644 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_91_203 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5806_ _1666_ _1669_ _2205_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_147_655 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4203__A1 _0723_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_45_620 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6786_ core_0.execute.rf.reg_outputs\[3\]\[3\] _3065_ _3057_ _3069_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3998_ core_0.execute.rf.reg_outputs\[1\]\[8\] _0627_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__inv_1
XANTENNA_clkbuf_leaf_107_i_clk_I clknet_4_4__leaf_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4754__A2 _1241_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5737_ _1715_ _2137_ core_0.decode.oc_alu_mode\[13\] _2138_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__5366__I _1809_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_60_601 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_44_163 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_115_552 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5668_ _2067_ _2068_ _2069_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_5_772 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_32_347 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_667 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_102_202 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_142_371 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7407_ net204 _3544_ _3569_ _3570_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__5703__A1 _1123_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4619_ _1175_ core_0.execute.alu_flag_reg.o_d\[1\] _1178_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_130_522 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4506__A2 _1094_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5599_ _1676_ _1641_ _2000_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_130_544 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7338_ _1172_ _3509_ _3510_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_0_229_431 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_130_577 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7456__A1 _3581_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7269_ _1742_ _3439_ _3449_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_51_1130 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_213_832 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_231_139 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_197_522 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_206_34 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4445__I core_0.decode.i_instr_l\[3\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_169_246 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_200_504 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_197_566 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_16_707 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_68_734 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_206_89 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_745 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_95_531 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_200_548 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_28_609 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_184_227 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4993__A2 _0767_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_67_266 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_55_417 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_138_644 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_138_655 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6195__A1 core_0.execute.pc_high_buff_out\[7\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_138_677 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6195__B2 net14 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_193_772 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_36_631 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_82_236 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_153_603 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_126_839 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_222_77 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_24_795 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_24_804 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_82_269 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5942__A1 core_0.execute.alu_mul_div.div_cur\[1\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_51_601 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4180__I _0798_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_35_174 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_23_336 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_152_168 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_106_574 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_121_500 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_51_667 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6498__A2 _1719_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7695__A1 _1078_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7705__B _1284_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50_155 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_50_188 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7447__A1 _3563_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_188_2769 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8311__CLK clknet_leaf_68_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_102_780 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_207_125 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_235_467 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_223_618 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6670__A2 _2999_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_235_489 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_223_629 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4681__A1 _0813_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_216_692 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_78_509 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6958__B1 _3178_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_240_3391 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4028__A4 core_0.execute.rf.reg_outputs\[5\]\[6\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5225__A3 _0776_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_203_364 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_58_200 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4970_ core_0.execute.sreg_priv_control.o_d\[12\] _1393_ _1422_ _1390_ _1423_ vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_86_531 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_EDGE_ROW_103_Left_350 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_175_216 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_58_244 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3921_ core_0.execute.rf.reg_outputs\[7\]\[14\] _0530_ _0556_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_199_2898 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6640_ core_0.execute.rf.reg_outputs\[7\]\[8\] _2962_ _1978_ _2982_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__6503__C _2113_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_144_625 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_73_258 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_210_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5933__A1 _1603_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6571_ _2926_ _0215_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_171_422 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_601 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_116_349 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_144_669 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8310_ _0486_ clknet_leaf_75_i_clk net180 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_4
XFILLER_0_26_174 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5522_ core_0.execute.hold_valid core_0.decode.o_submit _0754_ _1951_ vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__7615__B _1953_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_42_667 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_30_807 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_8241_ _0417_ clknet_4_9__leaf_i_clk core_0.execute.sreg_irq_pc.o_d\[13\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_76_1428 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_112_522 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5453_ core_0.execute.alu_mul_div.div_cur\[12\] _1812_ _1841_ _1890_ vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_2_731 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_112_533 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4404_ _0836_ _0947_ _0970_ _1012_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_8172_ _0348_ clknet_leaf_87_i_clk net94 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_4
XANTENNA__5161__A2 _1436_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5384_ core_0.execute.alu_mul_div.div_cur\[3\] _1811_ _1830_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__7438__A1 _3581_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7123_ _3320_ _3316_ _3329_ _3331_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4335_ _0892_ _0952_ _0953_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_10_553 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_10_597 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_7054_ _3266_ _3267_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_4266_ core_0.fetch.prev_request_pc\[15\] _0827_ _0884_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__4121__B1 _0736_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6005_ core_0.execute.pc_high_buff_out\[3\] _2249_ _2265_ core_0.execute.alu_flag_reg.o_d\[3\]
+ _2395_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__6661__A2 core_0.ew_data\[15\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_33_i_clk_I clknet_4_10__leaf_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_66_94 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4197_ _0725_ net38 _0815_ _0816_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_4
XFILLER_0_241_426 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_207_692 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_87_1557 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_96_317 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_222_673 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7610__A1 net216 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_173_62 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_96_339 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7956_ _0134_ clknet_leaf_19_i_clk core_0.execute.alu_mul_div.div_cur\[12\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_2
XANTENNA__4424__A1 _1024_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_139_408 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6907_ _2972_ _3129_ _3138_ _0339_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_7887_ _0078_ clknet_leaf_78_i_clk core_0.decode.i_instr_l\[12\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_2
XANTENNA__4975__A2 _0563_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_37_406 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_65_715 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_166_249 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_37_428 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6838_ core_0.execute.rf.reg_outputs\[2\]\[9\] _3092_ _3098_ _3099_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_9_352 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_175_772 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_64_236 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_108_839 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4727__A2 _1237_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5924__A1 _1559_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_64_269 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_664 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_80_729 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6769_ core_0.execute.rf.reg_outputs\[4\]\[12\] _3049_ _3057_ _3059_ vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_107_349 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_21_765 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_72_291 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_103_500 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output180_I net180 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7525__B _3651_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_667 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_143_680 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_149_Right_149 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_98_1686 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_32_155 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_60_475 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3950__A3 _0549_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_131_842 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_20_317 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_328 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_4_i_clk clknet_4_2__leaf_i_clk clknet_leaf_4_i_clk vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_13_391 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7429__A1 _3563_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6101__A1 net12 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_245_754 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6652__A2 core_0.ew_data\[12\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_205_618 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_125_2016 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_232_448 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_88_807 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_217_99 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_29_865 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_197_352 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_213_695 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_158_728 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_240_481 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_240_492 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4966__A2 _0604_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_107_1793 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_200_356 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_28_406 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6604__B _1978_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_218_3124 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_200_367 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_203 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4903__I _1225_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_56_737 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_68_597 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6168__A1 _1137_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_225 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_166_761 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_60_1229 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_83_556 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_153_411 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5915__A1 _1554_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_71_718 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_125_113 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_153_422 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_165_282 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_125_146 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_136_2145 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_102_69 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_23_122 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_125_179 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_153_488 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_807 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__7435__B _3553_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_667 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XPHY_EDGE_ROW_116_Right_116 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__7668__A1 core_0.dec_sreg_jal_over vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_106_382 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87_16 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_106_393 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_11_328 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6340__A1 _1379_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_121_352 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_229_3264 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_208_423 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4120_ core_0.execute.prev_pc_high\[0\] _0739_ _0740_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_236_754 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_235_231 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_71_1369 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_242_3420 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_235_264 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4051_ core_0.execute.rf.reg_outputs\[7\]\[4\] _0529_ _0676_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_236_798 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_223_415 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_208_489 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_147_2274 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4654__A1 net106 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput5 i_core_int_sreg[13] net5 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_36_53 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_127_66 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_160_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_189_842 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_160_2430 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_78_317 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7810_ core_0.dec_alu_carry_en _1053_ _3871_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_203_150 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_188_341 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_149_706 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__8207__CLK clknet_leaf_12_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_176_514 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_231_492 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_203_183 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_59_542 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7741_ net184 core_0.decode.i_imm_pass\[15\] _1063_ _3822_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4953_ core_0.execute.sreg_priv_control.o_d\[7\] _1394_ _1410_ _1391_ _1411_ vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__6514__B _1432_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_176_547 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_417 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_129_430 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_74_512 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_86_372 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3904_ core_0.dec_r_reg_sel\[1\] _0540_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__inv_4
XFILLER_0_129_441 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6159__A1 _2293_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7672_ _1431_ _1053_ _3774_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_163_208 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4884_ _1279_ _0727_ _1355_ _0099_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_0_52_96 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_191_539 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_247 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_82_1498 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_129_485 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_46_258 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6623_ core_0.execute.rf.reg_outputs\[7\]\[5\] _2962_ _1978_ _2968_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_117_636 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_156_271 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_46_269 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5906__A1 _2102_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_144_422 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_117_658 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_117_669 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_228 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_116_146 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_171_241 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6554_ net119 _2825_ _2906_ _2918_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__7108__B1 _1501_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5382__A2 _1814_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_116_168 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_54_291 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5505_ _1367_ _1937_ _1938_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_30_604 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_171_2570 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3932__A3 _0543_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_113_842 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6485_ _1380_ core_0.execute.sreg_irq_pc.o_d\[14\] _2864_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_30_615 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_14_177 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_112_341 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8224_ _0400_ clknet_leaf_16_i_clk core_0.execute.alu_flag_reg.o_d\[2\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_2
X_5436_ _1873_ _1874_ _1838_ _1875_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__5134__A2 net218 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_65_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6882__A2 _3108_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_8155_ _0331_ clknet_leaf_79_i_clk core_0.execute.rf.reg_outputs\[1\]\[14\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_77_60 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5367_ _1749_ _1808_ _1815_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7106_ _3305_ _3307_ _3314_ _3315_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_4318_ net69 core_0.fetch.out_buffer_data_instr\[9\] _0725_ _0936_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_77_93 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8086_ _0262_ clknet_leaf_105_i_clk core_0.execute.rf.reg_outputs\[5\]\[9\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5298_ core_0.decode.o_submit _0801_ _1746_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA_input37_I i_mem_exception vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_226_242 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6634__A2 core_0.ew_data\[7\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7037_ core_0.execute.alu_mul_div.mul_res\[7\] _3250_ _3251_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_4249_ net64 core_0.fetch.out_buffer_data_instr\[4\] _0724_ _0868_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_214_426 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4645__A1 _1195_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_241_212 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_184_72 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_241_267 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_179_341 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_179_352 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_195_812 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_179_374 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_26_824 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_96_158 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_84_309 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_218_Right_218 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
X_7939_ _0117_ clknet_leaf_41_i_clk core_0.execute.sreg_priv_control.o_d\[11\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5070__A1 _1461_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_46_1062 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_37_236 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_135_422 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_147_282 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_162_241 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_150_403 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_33_431 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_740 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_559 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_208_Left_455 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_213_3065 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_190_594 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_61_762 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_150_436 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_61_784 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3923__A3 _0544_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_626 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_283 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5125__A2 net232 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_131_661 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_103_396 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_131_2086 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6873__A2 _3114_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_185_2728 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_130_193 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_57_1191 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4884__A1 _1279_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_218_743 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_245_562 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_233_702 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_218_787 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_232_201 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_217_275 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_6_582 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_232_212 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_232_223 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_217_Left_464 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_73_18 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6318__C _2638_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_109_1822 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_189_138 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_186_801 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_232_289 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6389__A1 _1061_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_88_659 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_201_621 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_200_2909 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6389__B2 _1109_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_197_160 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_186_823 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_158_514 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_158_547 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4939__A2 net212 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_197_193 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5061__A1 _1466_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_201_676 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_196_2868 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_56_523 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_236 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_139_772 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xclkbuf_leaf_105_i_clk clknet_4_5__leaf_i_clk clknet_leaf_105_i_clk vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_28_247 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_865 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_56_578 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_EDGE_ROW_226_Left_473 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_154_753 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_3_314 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_113_127 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_773 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_475 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3914__A3 _0549_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_114 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6270_ _2346_ net208 _2654_ _2655_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_51_294 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5116__A2 net218 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5221_ _1666_ _1669_ _0769_ _1670_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_4
XTAP_TAPCELL_ROW_149_2303 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_121_182 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4875__A1 _0823_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7612__C _1217_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5152_ _1600_ _1601_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XPHY_EDGE_ROW_235_Left_482 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
X_4103_ core_0.fetch.out_buffer_valid _0723_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XANTENNA__7813__A1 _1034_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5083_ _1482_ _1491_ _1502_ _1531_ _1532_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_0_223_212 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_208_297 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4034_ net215 net206 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__inv_2
XFILLER_0_79_604 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4744__S _1236_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_84_1516 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4642__A4 _1200_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_177_812 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_204_481 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_84 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_188_193 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5985_ _1603_ _1639_ _2375_ _2376_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_93_106 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_192_804 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_59_372 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_176_355 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7724_ _3813_ _0481_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_59_394 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4936_ net201 _1398_ _1390_ _1399_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
XPHY_EDGE_ROW_244_Left_491 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_47_556 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7655_ _1078_ _1072_ _1105_ _3761_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_4867_ _0844_ core_0.decode.i_imm_pass\[9\] _1305_ _1347_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_170_85 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_34_217 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6606_ net23 _1148_ _2953_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_7_664 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_144_241 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_144_252 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7586_ _3704_ _3705_ _3675_ _3706_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__5355__A2 _1527_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6552__A1 net118 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_31_882 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_4798_ core_0.fetch.out_buffer_data_pred _1241_ _1304_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_7_697 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_172_594 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6537_ _2909_ _0198_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_144_296 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5374__I _1809_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_30_401 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_160_767 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_120_609 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_113_650 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5107__A2 net185 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_95_1656 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_179_72 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_434 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6468_ _2286_ _1713_ net214 _1455_ _2638_ _2847_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai221_2
X_8207_ _0383_ clknet_leaf_12_i_clk net79 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_4
XANTENNA__6855__A2 _3108_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5419_ _1747_ _1855_ _1860_ _0129_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_1
Xoutput150 net150 o_mem_data[5] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
Xclkbuf_leaf_84_i_clk clknet_4_12__leaf_i_clk clknet_leaf_84_i_clk vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
Xoutput161 net161 o_req_addr[0] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_30_489 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6399_ _1088_ _2777_ _2779_ _2332_ _2780_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai211_2
Xoutput172 net172 o_req_addr[5] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput183 net183 sr_bus_addr[14] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
X_8138_ _0314_ clknet_leaf_100_i_clk core_0.execute.rf.reg_outputs\[2\]\[13\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xoutput194 net194 sr_bus_data_o[0] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_227_562 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_215_702 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7804__A1 _0776_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_8069_ _0245_ clknet_leaf_106_i_clk core_0.execute.rf.reg_outputs\[6\]\[8\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_2
Xclkbuf_leaf_99_i_clk clknet_4_7__leaf_i_clk clknet_leaf_99_i_clk vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__7280__A2 _3458_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_3_552 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4094__A2 _0530_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5291__A1 net72 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_180_2669 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_242_576 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_230_727 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_39_982 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7032__A2 _1620_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_179_171 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_179_182 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_214_34 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_85_629 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_97_489 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_22_i_clk clknet_4_8__leaf_i_clk clknet_leaf_22_i_clk vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_194_141 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_104_1763 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5594__A2 _1994_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_182_314 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_194_174 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_66_865 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_194_196 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_504 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_81_813 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_2_i_clk_I clknet_4_0__leaf_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xwire211 _1718_ net211 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
Xclkbuf_leaf_37_i_clk clknet_4_11__leaf_i_clk clknet_leaf_37_i_clk vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__5346__A2 _1789_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_230_55 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_133_2104 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_230_66 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_190_380 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_163_594 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_378 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_59_1220 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_61_570 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_150_244 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6846__A2 _3092_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_115_1892 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
Xload_slew216 _0648_ net216 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XTAP_TAPCELL_ROW_226_3223 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4321__A3 _0937_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_206_702 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_205_212 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_245_392 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_233_532 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6048__C _1432_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_144_2244 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_17_66 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4085__A2 _0524_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_88_412 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5282__A1 _1431_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7023__A2 _1939_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_48_309 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_220_259 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5034__A1 core_0.dec_l_reg_sel\[2\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_88_489 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_124_34 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_185_130 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_174_804 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_201_473 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5770_ _2170_ _1568_ _2171_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_29_545 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_8_417 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_237_3352 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_8_428 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_191 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_124_89 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_8_439 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_185_196 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4721_ core_0.fetch.out_buffer_data_instr\[15\] _1261_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_29_578 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_123_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7440_ _3547_ _3596_ _3597_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_4_601 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_83_194 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5337__A2 _1754_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4652_ _1197_ _1199_ _1200_ _1210_ _1211_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or4_1
XFILLER_0_44_559 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_3_100 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_155_2373 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_154_594 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput30 i_mem_data[3] net30 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput41 i_req_data[12] net41 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
X_7371_ _1389_ _3392_ _3539_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or2_1
Xinput52 i_req_data[22] net52 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4583_ _1156_ net150 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput63 i_req_data[3] net63 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_40_721 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_4_667 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6322_ _2700_ _2703_ _2704_ _2705_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_0_40_765 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_229_827 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6253_ core_0.decode.oc_alu_mode\[3\] _1620_ _2638_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__4848__A1 core_0.decode.i_imm_pass\[0\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5204_ _1558_ _1652_ _1653_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_228_359 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_58_84 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6184_ _2569_ _2570_ _2571_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_0_110_686 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_209_562 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5135_ _1580_ _1581_ _1582_ _1583_ _1584_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and4_2
XANTENNA__4538__I core_0.decode.oc_alu_mode\[12\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_224_510 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_90_1597 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_224_543 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7262__A2 _3391_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5066_ _1466_ net190 _1515_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__5273__A1 _1480_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_28_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4076__A2 _0578_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_0_500 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_224_587 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_211_204 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4017_ _0567_ _0523_ _0526_ core_0.execute.rf.reg_outputs\[2\]\[7\] _0645_ vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_2
XTAP_TAPCELL_ROW_0_511 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_205_790 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_36_941 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_67_629 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_79_489 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5369__I _1816_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_94_448 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5576__A2 _1172_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5968_ _2355_ _2358_ _2359_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_191_100 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_865 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_149_388 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_176_174 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_191_122 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_43_1032 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_118_731 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7707_ _1034_ _3801_ _3804_ _0473_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4919_ net185 _1382_ _1197_ _1383_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_0_192_667 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5899_ _1059_ _2004_ _2285_ _1107_ _2290_ _2291_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_0_74_172 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_152_509 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7638_ _0748_ _3729_ _3749_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6525__A1 core_0.ew_data\[15\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_35_559 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5328__A2 _1695_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_7_472 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_145_583 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_191_199 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_687 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_250 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7569_ core_0.execute.pc_high_buff_out\[2\] _3682_ _3690_ _3691_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__4000__A2 core_0.execute.rf.reg_outputs\[4\]\[8\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_132_244 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_210_3035 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_30_220 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_30_231 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_120_428 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_160_597 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_31_765 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_132_299 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6828__A2 _3086_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_8_611 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7252__C _1736_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5500__A2 _1929_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_54_1161 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7789__B1 _3802_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7912__CLK clknet_leaf_81_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_89_209 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_3_6_0_i_clk_I clknet_0_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_81_i_clk_I clknet_4_13__leaf_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_230_502 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_199_255 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_202_215 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_221_3164 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_199_277 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_242_395 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_199_288 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7005__A2 _3177_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_202_259 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_97_286 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_167_130 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5567__A2 _0739_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_128_517 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_193_2827 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_167_174 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_54_802 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_183_634 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4775__B1 _0881_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_65_1290 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_155_336 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_182_133 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_183_656 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_109_753 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7308__A3 _3467_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_155_369 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_182_144 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_14_679 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_81_632 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_241 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_54_857 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_93_492 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5319__A2 _1600_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_170_317 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6516__B2 net7 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_124_723 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_136_594 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_34_570 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_117_1921 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_232_3293 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_111_406 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_480 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6819__A2 _3086_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_226_819 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_119_45 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_28_98 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_234_863 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4058__A2 _0541_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6940_ _1227_ _1715_ _3160_ _1230_ _3161_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai211_2
XANTENNA__6506__C _2626_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_607 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_135_66 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6871_ core_0.execute.rf.reg_outputs\[1\]\[7\] _3114_ _3112_ _3118_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_240_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5007__A1 _1131_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_186_450 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5822_ _1633_ _2218_ _2219_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_4
XTAP_TAPCELL_ROW_33_911 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_29_320 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5558__A2 _1956_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6755__A1 _2967_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_640 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_157_2402 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_201_292 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_146_325 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_174_634 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_91_418 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4766__B1 _0881_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5753_ _2151_ _2153_ _2154_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_56_150 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_60_30 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_247 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_72_610 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_162_807 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_174_667 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_621 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4704_ core_0.fetch.out_buffer_data_instr\[9\] net69 _1246_ _1250_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_17_548 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_161_317 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_17_559 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5684_ _2078_ _2083_ _2084_ _2085_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_161_328 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_142 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5138__B _0779_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7423_ _3563_ net85 _3553_ _3582_ _3583_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_114_222 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4635_ core_0.de_jmp_pred _1193_ _1194_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__7180__A1 _1926_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_79_1459 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_114_244 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_4_453 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_130_704 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7354_ _3523_ _0401_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_142_575 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_754 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_102_417 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4566_ _1146_ core_0.fetch.current_req_branch_pred vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__5730__A2 _2123_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4533__A3 _1069_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_142_597 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_92_1615 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_8_97 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_69_72 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6305_ core_0.execute.alu_mul_div.div_cur\[9\] _1117_ _2689_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_228_101 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7285_ net74 _3462_ _3463_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_40_584 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5652__I _1576_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4497_ _1088_ _1062_ _1089_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_110_450 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_168_2531 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7935__CLK clknet_leaf_32_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6236_ _1379_ _2620_ _2621_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_110_472 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4297__A2 _0914_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5494__A1 _1451_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_244_627 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_216_329 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_228_189 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6167_ _2024_ _2552_ _1458_ _2554_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_85_60 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_103_i_clk_I clknet_4_5__leaf_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5118_ _1561_ _1566_ _1567_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_6098_ core_0.ew_data\[4\] _2486_ _2487_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_224_351 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4049__A2 _0523_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5246__A1 _1461_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_240_822 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5049_ core_0.execute.rf.reg_outputs\[6\]\[12\] _1435_ _1486_ core_0.execute.rf.reg_outputs\[5\]\[12\]
+ _1498_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_196_203 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3900__I _0526_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6994__A1 _2436_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_196_225 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_169_439 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_95_702 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_196_247 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_output106_I net106 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_67_448 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5549__A2 _1957_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6746__A1 _2946_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_165_612 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_179_2660 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_101_1722 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_54_109 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6432__B _2133_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_75_481 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_165_689 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_164_177 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_35_356 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_734 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_28_i_clk_I clknet_4_10__leaf_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_23_507 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_11_649 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5048__B _0779_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_180_659 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3980__A1 _0534_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7010__I2 _1929_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_16_570 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7171__A1 _1369_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_106_778 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_277 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_562 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_120_247 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_219_134 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_219_156 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_112_1851 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_112_1862 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5485__A1 _1364_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_234_104 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_158_Left_405 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_235_638 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_234_115 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_128_2047 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7710__C _1283_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_141_2203 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_231_833 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_243_693 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_188_726 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_236_98 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_215_395 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_188_737 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6985__A1 _1372_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_19_738 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5788__A2 _1953_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6326__C _2090_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_205_2970 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5230__C _1678_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_230_365 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_230_387 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_14_34 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_105_47 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_168_461 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_640 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_128_314 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5004__A4 core_0.decode.oc_alu_mode\[2\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_123_1991 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_167_Left_414 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_234_3322 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6342__B core_0.dec_mem_access vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_54_610 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_144_807 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_156_667 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_6_707 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_155_144 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_26_334 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_139_2176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_171_626 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_356 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_142 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3971__A1 net90 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_81_462 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_136_391 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_152_2332 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_30_77 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_124_564 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_170_169 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4420_ net79 _1024_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_3
XFILLER_0_112_737 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_124_597 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4351_ _0959_ _0967_ _0968_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_22_584 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_238_421 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_238_454 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7070_ core_0.execute.alu_mul_div.mul_res\[9\] _3177_ _3173_ _3281_ _3178_ _1585_
+ _3282_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_0_1_489 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_176_Left_423 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__7465__A2 net77 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4282_ core_0.fetch.prev_request_pc\[15\] _0827_ _0886_ core_0.fetch.prev_request_pc\[14\]
+ _0899_ _0900_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_0_190_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_245_3451 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6021_ _2408_ _2410_ _2411_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__4088__I _0709_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_222_800 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5228__A1 _1625_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_240_107 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7399__I net37 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_240_118 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_206_373 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7768__A3 _3842_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_163_2472 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6976__A1 _3175_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7972_ _0149_ clknet_leaf_46_i_clk core_0.execute.mem_stage_pc\[7\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_89_551 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_77_702 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_89_562 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_221_354 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6923_ net93 _3128_ _3139_ _3147_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_178_247 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4451__A2 _1045_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_185_Left_432 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__6728__A1 _2986_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_77_768 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6854_ _3106_ _3108_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_146_111 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_174_431 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5805_ _2183_ _2195_ _2196_ _2203_ _2204_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_6785_ _2951_ _3064_ _3068_ _0287_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_3997_ _0626_ net209 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__4551__I _1133_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5736_ _1714_ _1695_ _1696_ _2137_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_0_91_248 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_134_317 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_162_626 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_146_177 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_161_114 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_44_142 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_95_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_17_378 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5667_ _1803_ _1501_ _2068_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_60_635 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_495 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_44_197 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4618_ _1175_ core_0.execute.alu_flag_reg.o_d\[0\] _1176_ _1177_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_142_361 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7406_ _1357_ _1013_ _3546_ _3568_ _3569_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_4_261 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5598_ _1997_ _1998_ _1999_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_4
XANTENNA__5703__A2 _1637_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_13_540 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_60_679 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6900__A1 _2956_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input67_I i_req_data[7] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_13_562 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_102_236 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7337_ core_0.dec_alu_flags_ie _3495_ _3509_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_229_410 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_194_Left_441 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_13_584 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_102_247 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4549_ _0812_ _1031_ _1132_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or2_4
XFILLER_0_40_370 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_130_589 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_187_72 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7268_ _1431_ _1415_ _1736_ _2662_ _3448_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XANTENNA__8113__CLK clknet_leaf_111_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_217_627 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6219_ _1699_ _2133_ _2604_ _2605_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_4
XTAP_TAPCELL_ROW_51_1120 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_7199_ _3386_ _2334_ _3387_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_244_457 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5219__A1 _0771_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_240_652 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_212_365 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_16_708 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_212_376 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_185_718 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_67_212 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_95_521 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6719__A1 _2972_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_779 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_138_623 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_67_278 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_222_34 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6195__A2 _2249_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_126_807 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_138_667 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7392__A1 core_0.execute.sreg_irq_pc.o_d\[1\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_62_1260 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_152_103 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_24_796 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5942__A2 _2279_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_180_423 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_142 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_153_648 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_152_136 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_50_123 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7695__A2 _1095_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_106_597 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_133_383 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_121_578 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7447__A2 net74 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_101_291 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_235_446 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_207_137 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_222_107 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6407__B1 _2534_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_204_822 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4636__I core_0.dec_sreg_irt vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6958__A1 core_0.execute.alu_mul_div.mul_res\[0\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6958__B2 _1451_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_702 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_240_3392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_116_68 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_231_685 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_25_66 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5630__A1 _1715_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_735 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_58_223 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_88 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3920_ _0534_ _0535_ _0536_ core_0.execute.rf.reg_outputs\[6\]\[14\] _0555_ vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_0_25_99 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_59_768 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_169_781 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_199_2899 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_73_204 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_129_667 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_132_34 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7383__A1 _1357_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_621 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_156_453 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4197__A1 _0725_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_184_784 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_116_317 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_128_177 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6570_ core_0.dec_rf_ie\[5\] core_0.ew_reg_ie\[5\] _2201_ _2926_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_26_131 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_6_559 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_144_659 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5521_ _1948_ _0807_ _1949_ _1950_ _0141_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_27_698 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7135__A1 _2855_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_143_158 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_203_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6800__B _3072_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_54_495 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_171_478 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8240_ _0416_ clknet_leaf_41_i_clk core_0.execute.sreg_irq_pc.o_d\[12\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_14_348 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5452_ core_0.execute.alu_mul_div.div_cur\[11\] _1814_ _1817_ _1888_ _1889_ vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_41_156 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_76_1429 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8136__CLK clknet_leaf_103_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5697__A1 _1123_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4403_ _0959_ _0950_ _1010_ _1011_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or3_1
X_8171_ _0347_ clknet_leaf_87_i_clk net93 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_4
XFILLER_0_140_865 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_151_191 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5383_ _1748_ _1825_ _1829_ _0124_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_7122_ _3320_ _3316_ _3329_ _3330_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_0_112_589 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4334_ core_0.fetch.prev_request_pc\[9\] core_0.fetch.prev_request_pc\[8\] _0951_
+ _0952_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_0_10_543 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_157_20 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_226_413 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7053_ _2648_ _3265_ _3266_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_4265_ _0882_ _0883_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_66_51 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8286__CLK clknet_leaf_32_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_226_457 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6004_ _2202_ _2393_ _2394_ _0180_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4196_ _0724_ _0814_ _0815_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_87_1558 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7610__A2 _3675_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_10_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_179_556 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_221_151 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7955_ _0133_ clknet_leaf_19_i_clk core_0.execute.alu_mul_div.div_cur\[11\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_49_212 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4424__A2 _0970_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5621__A1 _1761_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6906_ net100 _3135_ _3124_ _3138_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_7886_ _0077_ clknet_leaf_81_i_clk core_0.decode.i_instr_l\[11\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_194_559 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_37_418 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_727 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_278 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_176_2630 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6837_ _0722_ _3098_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_108_807 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xclkbuf_4_4__f_i_clk clknet_3_2_0_i_clk clknet_4_4__leaf_i_clk vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_18_621 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7374__A1 _1953_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_135_604 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_181_209 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_364 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_80_708 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_190_732 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6768_ _2988_ _3043_ _3058_ _0280_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_80_719 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_17_142 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_135_648 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_190_754 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_782 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3935__A1 _0568_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_21_766 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_5719_ _1124_ _1585_ _2091_ _2092_ _2120_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai211_2
XANTENNA__7126__A1 _3189_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6699_ _2994_ _3000_ _3018_ _0251_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_190_798 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_143_670 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7677__A2 _1094_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_679 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_98_1687 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5688__A1 _1479_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_60_465 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output173_I net173 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_60_487 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_198_82 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7429__A2 net86 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4360__A1 _0970_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_217_413 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7541__B _1357_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6101__A2 _2260_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_245_766 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_232_416 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_217_34 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_204_107 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_125_2017 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5860__A1 _1382_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_123 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4456__I net71 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_29_855 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5996__B _0798_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_201_814 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_29_866 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_87_329 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4415__A2 core_0.fetch.prev_request_pc\[0\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_202_2940 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5612__A1 _1929_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4392__S _0959_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_96_863 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_212_195 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_107_1794 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_157_228 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_233_66 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_185_559 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_218_3125 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_95_373 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_535 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_138_453 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5287__I _1735_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_120_1950 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_172_209 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_237 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_138_486 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5915__A2 _1576_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_451 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8159__CLK clknet_leaf_88_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_64_782 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_102_37 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__3926__A1 _0534_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7716__B _3809_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_136_2146 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7117__A1 _1225_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_141_607 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_153_467 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_181_776 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_141_629 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_23_134 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6112__S _2293_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_106_372 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7668__A2 _1062_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_122_865 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5951__S _2342_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4351__A1 _0959_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_863 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_229_3265 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_71_1359 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_242_3421 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_235_243 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_208_457 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4050_ _0516_ core_0.execute.rf.reg_outputs\[3\]\[4\] net231 _0675_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
XTAP_TAPCELL_ROW_147_2275 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
Xinput6 i_core_int_sreg[14] net6 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_36_76 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_160_2431 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_204_663 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5603__A1 _1558_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_153_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4952_ _1400_ net216 _1410_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_7740_ _3821_ _0489_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_203_195 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_59_554 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_148_228 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_143_66 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3903_ _0517_ _0539_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_46_215 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_74_524 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7356__A1 _2646_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_86_384 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7671_ _1078_ _1080_ _3773_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_143_88 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4883_ core_0.decode.i_flush core_0.fetch.dbg_out core_0.fetch.flush_event_invalidate
+ _1355_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_86_395 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6622_ _2930_ core_0.ew_data\[5\] _2966_ _2967_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_4
XFILLER_0_6_301 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_62_708 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_82_1499 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_6_312 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_579 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_462 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_15_602 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_144_434 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_613 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3917__A1 net94 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_6_345 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6553_ _2209_ _2783_ _2917_ _0206_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__7108__A1 _3149_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_116_158 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_6_367 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7108__B2 _3209_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_131_106 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5504_ _1933_ _1936_ _1229_ _1937_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_171_2560 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_171_286 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6484_ net77 _2531_ _2862_ _2537_ _2863_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_131_128 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7659__A2 _1053_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_42_465 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8223_ _0399_ clknet_leaf_8_i_clk core_0.execute.alu_flag_reg.o_d\[1\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_2
X_5435_ _1233_ _1868_ _1874_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4342__A1 _0827_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_77_50 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8154_ _0330_ clknet_leaf_95_i_clk core_0.execute.rf.reg_outputs\[1\]\[13\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_2
X_5366_ _1809_ _1814_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_58_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_77_72 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4893__A2 _1305_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4317_ net67 core_0.fetch.out_buffer_data_instr\[7\] _0725_ _0935_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_7105_ _2778_ _3313_ _3314_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_8085_ _0261_ clknet_leaf_108_i_clk core_0.execute.rf.reg_outputs\[5\]\[8\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_2
X_5297_ _1419_ _1745_ _0122_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__7292__B1 _3399_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7036_ _1371_ _3249_ _3250_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4248_ _0865_ _0866_ _0867_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_241_202 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_242_747 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_198_128 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4179_ core_0.execute.alu_mul_div.i_div _0798_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_241_246 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_93_82 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_97_627 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_241_279 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7595__A1 core_0.execute.pc_high_out\[5\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6398__A2 _2778_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6705__B _3016_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_182_Right_182 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_26_825 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_7938_ _0116_ clknet_leaf_41_i_clk core_0.execute.sreg_priv_control.o_d\[10\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_78_863 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_167_537 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_77_362 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5070__A2 net205 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_37_204 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7869_ _0061_ clknet_leaf_63_i_clk core_0.fetch.prev_request_pc\[12\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_46_1063 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7347__A1 _3510_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8301__CLK clknet_leaf_12_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_154_209 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_150 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_14_Right_14 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_163_721 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_203_69 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_172 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_80_516 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_46_782 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_527 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XPHY_EDGE_ROW_122_Left_369 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_135_489 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_213_3066 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_162_286 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_60_240 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_60_251 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA_output98_I net98 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_487 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_865 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_60_295 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_137 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4333__A1 core_0.fetch.prev_request_pc\[7\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_131_2087 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_185_2729 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_57_1192 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6666__I _2998_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4884__A2 _0727_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_218_733 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_245_530 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_23_Right_23 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__5570__I _1283_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6086__A1 core_0.decode.oc_alu_mode\[11\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_131_Left_378 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_6_583 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5833__A1 net136 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4186__I net156 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_109_1823 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_224_3195 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_232_268 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_220_419 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_87_115 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_198_662 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6389__A2 _1701_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_241_780 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87_137 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4914__I core_0.dec_sreg_irt vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_200_143 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5061__A2 _0597_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_200_154 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_32_Right_32 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_201_699 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_196_2869 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7338__A1 _1172_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_84_855 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_95_192 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_200_198 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_22_34 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_126_401 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_56_568 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_140_Left_387 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_22_45 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6010__A1 net81 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_153_220 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6010__B2 _2245_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_153_242 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_189_18 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_114_607 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_181_562 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_36_281 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_52_741 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_153_264 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_154_798 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_141_415 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4572__A1 core_0.ew_data\[0\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_113_117 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_24_454 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_76_i_clk_I clknet_4_13__leaf_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_465 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_12_605 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_113_139 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_11_104 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_12_649 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6313__A2 _2695_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_137 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_121_150 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5220_ _0771_ _0773_ _1667_ _1668_ _1669_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai31_4
XFILLER_0_228_519 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_41_Right_41 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_149_2304 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_20_660 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4875__A2 _1321_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6576__I core_0.ew_mem_access vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5151_ _1599_ _1600_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_236_541 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4102_ _0721_ _0722_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_47_53 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_209_788 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5082_ _1520_ _1525_ _1530_ _1531_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_0_138_77 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4033_ _0652_ _0657_ _0659_ _0660_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_0_223_257 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_211_408 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_79_627 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_211_419 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_78_115 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_189_662 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7577__A1 core_0.execute.pc_high_buff_out\[3\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_84_1517 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_188_172 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_231_290 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_50_Right_50 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_59_340 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_3_i_clk clknet_4_2__leaf_i_clk clknet_leaf_3_i_clk vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_94_619 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5984_ _1689_ _1665_ _1677_ _1603_ _2375_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_87_660 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7723_ net190 core_0.decode.i_imm_pass\[6\] _1946_ _3813_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_59_384 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4935_ _0731_ _1398_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_74_321 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_170_53 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_191_337 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_35_719 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7654_ _1102_ _3760_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_191_348 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_632 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4866_ _1346_ _0090_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_34_207 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6605_ _2936_ _2951_ _2952_ _0223_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_34_229 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4797_ _1301_ _1303_ _0064_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_7585_ core_0.execute.pc_high_buff_out\[4\] _3682_ _3705_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6552__A2 _1985_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_31_883 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_105_629 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_172_584 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6536_ net125 _2482_ _2906_ _2909_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_15_454 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_42_251 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_465 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_560 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_113_640 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_42_273 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_95_1657 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6467_ _1713_ net214 _2846_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6304__A2 _2332_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7501__A1 core_0.execute.sreg_scratch.o_d\[2\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_30_446 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_219_508 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8206_ _0382_ clknet_leaf_129_i_clk core_0.execute.alu_mul_div.div_res\[15\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_30_457 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_88_93 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_101_835 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_112_161 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xoutput140 net140 o_mem_data[10] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
X_5418_ core_0.execute.alu_mul_div.div_cur\[6\] _1838_ _1816_ _1859_ _1860_ vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__7803__C _1133_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput151 net151 o_mem_data[6] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
X_6398_ _1433_ _2778_ _2779_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xoutput162 net162 o_req_addr[10] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
Xoutput173 net173 o_req_addr[6] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
Xoutput184 net184 sr_bus_addr[15] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
X_8137_ _0313_ clknet_leaf_99_i_clk core_0.execute.rf.reg_outputs\[2\]\[12\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5349_ core_0.execute.alu_mul_div.div_cur\[13\] _1528_ _1529_ _1797_ vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_2
Xoutput195 net195 sr_bus_data_o[10] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_10_170 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3903__I _0517_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6068__A1 _2403_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_195_72 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7804__A2 _1134_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_215_714 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8068_ _0244_ clknet_leaf_107_i_clk core_0.execute.rf.reg_outputs\[6\]\[7\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_227_585 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4618__A2 core_0.execute.alu_flag_reg.o_d\[0\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output136_I net136 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_214_224 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_199_426 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7019_ _3222_ _3181_ _3234_ _0355_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__4174__S0 _0769_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_215_769 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_3_553 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_230_706 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_104 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_97_413 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5291__A2 _0810_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_202_419 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_97_424 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_168_802 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_223_780 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_186_109 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7568__A1 _3682_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_39_983 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_179_150 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_69_159 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_195_632 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_107 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6240__A1 _2356_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_513 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_167_356 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_78_693 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_38_535 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_104_1764 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_194_164 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_855 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_93_652 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_423 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_25_207 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_92_151 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7266__B _1395_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xwire212 net213 net212 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_230_34 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7841__CLK clknet_leaf_67_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_80_335 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_81_858 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_163_562 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_92_195 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_34_741 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_133_2105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4554__A1 _1131_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_763 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_191_2799 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_59_1221 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_150_234 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_402 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_103_150 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_150_289 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_131_492 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_115_1893 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4857__A2 _1341_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4909__I _1373_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_226_3224 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4321__A4 _0938_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_218_563 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_245_360 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_205_224 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_144_2245 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_108_69 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_205_257 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4085__A3 _0527_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_88_402 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5282__A2 _1729_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_177_109 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_88_457 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_158_301 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_198_481 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_158_312 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_213_290 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_201_430 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_186_654 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5034__A2 core_0.dec_l_reg_sel\[1\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_682 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_185_142 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_29_524 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_158_367 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_33_66 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_56_321 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_173_304 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_237_3353 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_56_332 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6782__A2 _3065_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_29_557 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_652 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_127_710 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_185_186 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4720_ _1259_ _1237_ _1260_ _0030_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_33_99 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_527 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_56_387 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4651_ _1209_ net192 _1210_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_83_184 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_140_34 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5475__I core_0.execute.alu_mul_div.cbit\[0\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_142_713 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_25_741 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_116_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xinput20 i_mem_ack net20 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_155_2374 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
Xinput31 i_mem_data[4] net31 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4582_ core_0.ew_data\[5\] net157 _1156_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_24_240 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7370_ core_0.execute.irq_en _1389_ _3538_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xinput42 i_req_data[13] net42 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_24_251 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput53 i_req_data[23] net53 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xinput64 i_req_data[4] net64 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_4_679 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6321_ _2372_ _2642_ _2704_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_12_457 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6298__A1 _1107_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6252_ _1756_ _1592_ _2637_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_122_492 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_0_852 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5203_ net217 _1650_ _1651_ _1652_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XANTENNA__4848__A2 _1307_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5424__B _1841_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6183_ core_0.execute.alu_mul_div.div_cur\[6\] _2279_ _2570_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__7247__B1 _2571_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5134_ core_0.execute.rf.reg_outputs\[1\]\[9\] net218 _1486_ core_0.execute.rf.reg_outputs\[5\]\[9\]
+ core_0.execute.rf.reg_outputs\[6\]\[9\] _1435_ _1583_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XTAP_TAPCELL_ROW_90_1587 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_224_500 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_90_1598 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7798__A1 _1120_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_236_382 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5065_ _0641_ _0646_ _0647_ _1459_ _1514_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai31_4
X_4016_ _0533_ _0541_ _0543_ core_0.execute.rf.reg_outputs\[5\]\[7\] _0644_ vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_0_79_413 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_0_501 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_74_84 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_0_512 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_189_492 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_177_632 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_36_942 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_181_30 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_107 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_181_63 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5967_ _2356_ _2357_ _2358_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_48_855 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_59_192 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_90_72 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6773__A2 _3041_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_181_96 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4784__A1 _1290_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7706_ core_0.dec_mem_we _1053_ _3804_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4918_ net178 _1382_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_4
XTAP_TAPCELL_ROW_43_1033 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_47_376 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5898_ _2286_ _1603_ _1653_ _1686_ _2289_ _2290_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai221_2
XFILLER_0_63_836 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7637_ _3732_ _3747_ _3748_ _0459_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_191_167 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_133_702 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_35_549 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_462 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_63_858 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_90_644 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5385__I _1765_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_145_562 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4849_ _0851_ _1306_ _1337_ _0082_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__6525__A2 _1985_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_117_275 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_132_201 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4536__A1 _1121_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5584__I0 core_0.dec_mem_we vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7568_ _3682_ _3688_ _3689_ _3690_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_0_31_711 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4000__A3 _0520_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_210_3036 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6519_ net78 _2531_ _2896_ _2537_ _2897_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_7499_ core_0.execute.sreg_scratch.o_d\[1\] _3641_ _3516_ _3643_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_30_243 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_690 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_8_612 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_101_632 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_113_492 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_219_349 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_30_298 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_234_308 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_54_1162 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_234_319 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_104_i_clk clknet_4_5__leaf_i_clk clknet_leaf_104_i_clk vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_227_360 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_215_511 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7789__A1 core_0.decode.i_instr_l\[13\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7789__B2 core_0.decode.i_instr_l\[10\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_243_842 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_227_393 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_199_212 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_24_i_clk_I clknet_4_8__leaf_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_215_566 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6461__A1 _1121_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_203_728 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_225_34 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_230_536 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_221_3165 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_202_227 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_119_i_clk clknet_4_6__leaf_i_clk clknet_leaf_119_i_clk vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_225_67 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6213__A1 _2286_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_85_416 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_211_772 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6213__B2 _1686_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_167_142 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6764__A2 _3049_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_195_484 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_109_710 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_193_2828 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_155_326 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_156_849 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_167_186 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_65_1291 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_66_663 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4775__B2 net172 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_365 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_505 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_685 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_241_66 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_26_527 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_387 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5509__B _1941_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_241_88 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6516__A2 _2579_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_53_346 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7713__A1 core_0.decode.i_imm_pass\[1\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4527__A1 _1114_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_53_368 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_123_212 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_688 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_117_1911 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_117_1922 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_232_3294 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_34_582 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_110_37 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_0_104 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_1_627 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_276 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_21_298 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_206_522 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6854__I _3106_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_233_352 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6452__A1 _1380_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4058__A3 _0543_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4374__I net73 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6870_ _2972_ _3107_ _3117_ _0323_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_159_632 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_48_107 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6204__A1 _2018_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5007__A2 _1455_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_202_772 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5821_ core_0.execute.rf.reg_outputs\[1\]\[4\] _1615_ _2218_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_233_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_33_912 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6755__A2 _3042_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_201_282 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_83_i_clk clknet_4_12__leaf_i_clk clknet_leaf_83_i_clk vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__4766__B2 net168 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5752_ _1715_ _1631_ _2152_ _2153_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_158_197 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_57_685 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_45_836 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_44_313 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_387 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_57_696 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_60_53 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4703_ _1249_ _0024_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_44_324 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_45_858 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_115_702 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_127_562 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_151_88 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5683_ _1993_ _1995_ _2084_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__7704__A1 _3786_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_4_410 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4518__A1 _1107_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7422_ _3547_ _1968_ _3582_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4634_ core_0.dec_jump_cond_code\[3\] _1185_ _1188_ _1191_ _1192_ _1193_ vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai221_4
XFILLER_0_60_839 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xclkbuf_leaf_98_i_clk clknet_4_7__leaf_i_clk clknet_leaf_98_i_clk vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__7180__A2 _3373_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_13_722 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4565_ _0727_ _0947_ _1145_ _1146_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XANTENNA__5191__A1 _1596_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7353_ _1217_ _3521_ _3522_ _3523_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and3_1
XTAP_TAPCELL_ROW_92_1616 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6304_ core_0.execute.alu_mul_div.div_res\[9\] _2332_ _2279_ _2688_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_40_563 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7284_ _1742_ _3454_ _3462_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4496_ core_0.execute.alu_mul_div.i_mul _1088_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
Xclkbuf_leaf_21_i_clk clknet_4_8__leaf_i_clk clknet_leaf_21_i_clk vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XPHY_EDGE_ROW_4_Right_4 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_100_92 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_168_2532 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6235_ net86 _2531_ _2619_ _2537_ _2620_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_12_298 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_682 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5494__A2 _1926_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6166_ _2024_ _2552_ _2553_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_85_72 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_176_85 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_225_842 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5117_ _1562_ _1563_ _1564_ _1565_ _1566_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and4_2
X_6097_ _2201_ _2486_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XANTENNA_clone1_I net222 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_36_i_clk clknet_4_11__leaf_i_clk clknet_leaf_36_i_clk vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__4049__A3 _0526_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5246__A2 net204 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_224_363 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5048_ _0789_ core_0.execute.rf.reg_outputs\[4\]\[12\] _0779_ _1497_ vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA_input12_I i_core_int_sreg[5] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6994__A2 _3181_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_67_405 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_79_265 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_79_276 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_427 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_95_736 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_149_142 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_179_2661 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6999_ _3153_ _3215_ _1366_ _3216_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__6746__A2 _3042_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_95_769 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_220_591 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_101_1723 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_164_123 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_192_454 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_47_184 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_11_639 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_152_329 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4509__A1 _1037_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7010__I3 _1631_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_51_828 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3980__A2 _0542_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7171__A2 _1227_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_63_699 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8192__CLK clknet_leaf_129_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5182__A1 _1446_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_160_384 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output80_I net80 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_219_102 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_120_259 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_112_1852 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6682__A1 _2972_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_128_2048 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_215_330 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_215_352 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_236_66 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_203_503 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_188_705 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5511__C _1841_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_141_2204 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_230_311 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_242_171 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6985__A2 _1367_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_19_739 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_205_2971 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_67_1320 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4996__A1 core_0.dec_l_reg_sel\[2\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_405 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_85_224 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_156_602 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6623__B _1978_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6737__A2 _3020_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4922__I _1385_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4748__A1 net58 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_123_1992 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_155_112 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5945__B1 _2250_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_234_3323 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_27_836 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_94_780 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_696 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5239__B _1061_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_858 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_139_2177 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_53_132 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_595 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_30_34 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3971__A2 _0578_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_42_839 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_54_699 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_121_69 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_152_2333 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_112_705 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7454__B _3545_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5173__A1 _1553_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_349 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_201_80 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_151_384 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4350_ core_0.fetch.prev_request_pc\[14\] _0956_ _0967_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__4920__A1 _1196_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_238_444 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4281_ _0887_ _0897_ _0898_ _0899_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_120_782 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6020_ _2300_ _2409_ _2410_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or2_1
XTAP_TAPCELL_ROW_245_3452 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input4_I i_core_int_sreg[12] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_219_680 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_183_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_225_138 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_207_842 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_234_650 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5228__A2 _1676_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_42 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_234_683 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_222_823 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7971_ _0148_ clknet_leaf_38_i_clk core_0.execute.mem_stage_pc\[6\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_163_2473 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_233_171 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_221_322 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6976__A2 _3189_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_233_193 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_221_333 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8065__CLK clknet_leaf_111_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4987__A1 _0770_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6922_ _2992_ _3130_ _3146_ _0346_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_221_388 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_187_760 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_193_207 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6853_ _3106_ _3107_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XANTENNA__6728__A2 _3022_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_202_591 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_159_484 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_63 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6025__S _1603_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5804_ _1987_ _2183_ _2203_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_147_646 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6784_ core_0.execute.rf.reg_outputs\[3\]\[2\] _3065_ _3057_ _3068_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_119_348 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3996_ _0619_ _0624_ _0625_ _0626_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_0_91_216 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_135_808 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_9_568 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_57_482 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_45_644 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5735_ _2090_ _2114_ _2135_ _2136_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_4
XFILLER_0_161_104 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_162_638 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_45_666 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_368 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7902__CLK clknet_leaf_68_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5666_ _1803_ _1500_ _2067_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_45_699 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_88_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5164__A1 _1446_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7405_ _1357_ core_0.execute.mem_stage_pc\[4\] _3568_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_32_349 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_4_251 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4617_ core_0.dec_jump_cond_code\[0\] _1176_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_2
X_5597_ _1479_ _1931_ _1998_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__6900__A2 _3129_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_13_552 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_130_524 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_142_384 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_130_535 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4911__A1 _1369_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7336_ _3494_ _3496_ _3508_ _1950_ _0398_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_4548_ core_0.decode.oc_alu_mode\[3\] _1131_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_0_229_422 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_40_382 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_229_455 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7267_ _2690_ _3391_ _3447_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4479_ _1069_ _1071_ _1072_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_4
XANTENNA__5467__A2 _1838_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6664__A1 core_0.ew_reg_ie\[6\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6218_ _2432_ _2603_ _2293_ _2604_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_51_1121 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_7198_ _1209_ _3386_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_244_469 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6149_ _2532_ _2533_ _2535_ _2536_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__6416__A1 _2576_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5219__A2 _0768_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_327 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_231_119 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_212_311 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_79_Right_79 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__4978__A1 _1381_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_240_664 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_169_248 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_240_686 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_16_709 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_67_224 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6443__B _1114_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6719__A2 _3021_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_67_246 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_95_555 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_178_782 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_184_229 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_55_419 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_82_205 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_48_471 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7392__A2 _3543_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_165_454 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_82_238 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_62_1261 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_75_290 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_153_627 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_222_79 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_24_797 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_106_521 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_180_435 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_91_772 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3953__A2 _0530_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_839 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_50_102 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_180_457 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_63_496 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_88_Right_88 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_134_863 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7274__B net73 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_51_647 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5155__A1 _0782_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_161_660 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_349 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_239_208 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_160_170 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4902__A1 _1367_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_121_546 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4410__C _0877_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_208_606 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6655__B2 net25 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_235_414 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_196_Right_196 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_73_1390 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4917__I _1380_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4130__A2 _0743_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8088__CLK clknet_leaf_104_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_216_661 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_97_Right_97 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_222_119 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6407__B2 net4 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_216_683 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_243_480 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_216_694 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6958__A2 _3177_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7080__A1 _3149_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4969__A1 _1381_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_240_3393 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_58_202 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5630__A2 _1934_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_231_697 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_175_207 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_203_399 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_129_613 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_58_257 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_706 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_169_793 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_39_460 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_67_780 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7383__A2 net72 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4197__A2 net38 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_17_Left_264 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_73_238 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_132_57 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5394__A1 _1233_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_66 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_6_527 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_128_189 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_171_424 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_41_88 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5520_ _1051_ _1950_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_183_295 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_260 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7135__A2 _3181_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_81_282 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_42_647 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7184__B core_0.execute.alu_mul_div.div_res\[11\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
X_5451_ _1375_ _1886_ _1887_ _1822_ _1888_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_152_671 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_76_1419 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_112_524 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4402_ core_0.fetch.prev_request_pc\[4\] _1009_ core_0.fetch.prev_request_pc\[5\]
+ _1010_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__5697__A2 _1934_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6894__A1 _2940_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_140_855 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8170_ _0346_ clknet_leaf_84_i_clk net92 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_2
X_5382_ core_0.execute.alu_mul_div.div_cur\[1\] _1814_ _1817_ _1828_ _1829_ vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_100_708 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7121_ _2797_ _3328_ _3329_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_4333_ core_0.fetch.prev_request_pc\[7\] core_0.fetch.prev_request_pc\[6\] _0950_
+ _0951_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_0_238_241 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1_276 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_10_566 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6646__B2 net22 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4264_ core_0.fetch.pc_flush_override core_0.decode.i_flush _0882_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_7052_ _3261_ _1451_ _3263_ _3264_ _3265_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XPHY_EDGE_ROW_26_Left_273 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_226_436 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_66 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_66_41 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_157_65 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6003_ core_0.ew_data\[2\] _2209_ _2394_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_EDGE_ROW_163_Right_163 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__4121__A2 _0735_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4827__I _1305_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4195_ core_0.fetch.out_buffer_data_instr\[0\] _0814_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xcore0_220 o_mem_addr_high[7] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_0_207_672 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_87_1559 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_96_308 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_210_804 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7954_ _0132_ clknet_leaf_19_i_clk core_0.execute.alu_mul_div.div_cur\[10\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_2
XANTENNA__5621__A2 _1613_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_77_533 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6905_ _2967_ _3129_ _3137_ _0338_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_194_527 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_166_218 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7885_ _0076_ clknet_leaf_50_i_clk core_0.decode.i_instr_l\[10\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_77_566 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_35_Left_282 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
X_6836_ _2981_ _3086_ _3097_ _0309_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_175_741 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_176_2620 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_77_599 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7374__A2 _3540_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_18_633 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4188__A2 net20 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_45_430 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6767_ core_0.execute.rf.reg_outputs\[4\]\[11\] _3049_ _3057_ _3058_ vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3979_ _0568_ core_0.execute.rf.reg_outputs\[3\]\[10\] _0549_ _0610_ vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_0_45_452 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_772 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_162_435 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_174_295 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5718_ _1124_ _2053_ _2091_ _2092_ _2119_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai211_2
XANTENNA__7806__C _1279_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_162_457 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_21_767 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6698_ core_0.execute.rf.reg_outputs\[6\]\[14\] _2998_ _3016_ _3018_ vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_134_159 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_33_636 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_115_340 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_116_863 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5137__A1 core_0.execute.rf.reg_outputs\[2\]\[8\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_32_135 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5649_ _2046_ _2049_ _2050_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_103_513 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5393__I _1809_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_32_146 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3906__I _0541_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_98_1688 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6885__A1 _2992_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_319 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_41_680 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7319_ net78 _3487_ _3384_ _3493_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XPHY_EDGE_ROW_44_Left_291 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_130_387 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8299_ _0475_ clknet_leaf_16_i_clk net178 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_4
XFILLER_0_245_712 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_187_2760 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_229_274 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_244_200 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_130_Right_130 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_125_2007 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_125_2018 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_244_288 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5860__A2 net186 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_217_68 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_99_146 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7062__A1 _1909_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_29_856 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_213_675 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_202_2941 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5612__A2 _1683_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_197_398 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_185_538 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_wire215_I _0660_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_107_1795 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_138_410 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4472__I core_0.decode.i_instr_l\[0\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_178_590 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_218_3126 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_28_419 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_588 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_95_385 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_4_6__f_i_clk_I clknet_3_3_0_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4405__C _0877_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7365__A2 _3533_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_120_1951 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5376__A1 core_0.execute.alu_mul_div.div_cur\[0\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_64_750 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_138_498 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3926__A2 _0542_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_136_2147 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_181_766 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_125_159 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_422 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5128__A1 _1482_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_140_107 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_180_287 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_384 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6876__A1 _2983_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_133_170 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_122_855 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_32_691 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_121_376 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_229_3255 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6628__A1 _2930_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_236_723 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_229_3266 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_242_3411 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_242_3422 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_235_255 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_235_277 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_147_2276 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
Xinput7 i_core_int_sreg[15] net7 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA_clkbuf_leaf_72_i_clk_I clknet_4_13__leaf_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7053__A1 _2648_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_160_2432 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_203_130 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_87_820 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_203_163 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_188_365 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5603__A2 _1652_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_691 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_188_376 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_87_842 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4951_ _1301_ _1409_ _0112_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__6083__B _1456_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_176_527 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_188_387 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_47_706 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_129_410 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_146_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_74_503 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3902_ _0522_ _0528_ _0531_ _0537_ _0538_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai211_4
XFILLER_0_19_419 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7670_ _3771_ _3772_ _0468_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4882_ _0876_ _1136_ _0727_ _0881_ _0098_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai31_1
XANTENNA__7356__A2 _2684_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6621_ _2929_ _2964_ _2965_ _2966_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_0_46_249 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8103__CLK clknet_leaf_94_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_117_627 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_290 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_7_836 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_74_569 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_116_104 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_55_750 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_116_115 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_172_733 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_184_593 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_116_126 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_6_335 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_858 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_55_772 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_156_295 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_171_221 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_474 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3917__A2 _0521_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6552_ net118 _1985_ _2917_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_15_625 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_144_457 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5503_ _1908_ _1613_ _1935_ _1936_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_54_293 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_171_276 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_232_Right_232 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
X_6483_ _2447_ _2860_ _2861_ _2862_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
XTAP_TAPCELL_ROW_171_2561 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_8222_ _0398_ clknet_leaf_16_i_clk core_0.execute.alu_flag_reg.o_d\[0\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_2
X_5434_ _1375_ _1872_ _1873_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_140_663 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_842 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4342__A2 _0959_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_8153_ _0329_ clknet_leaf_96_i_clk core_0.execute.rf.reg_outputs\[1\]\[12\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_2_585 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5365_ core_0.execute.alu_mul_div.div_cur\[1\] _1812_ _1813_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_100_527 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_112_387 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6619__A1 net25 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7104_ _3311_ _3312_ _3313_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_227_723 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4316_ _0929_ _0933_ _0934_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_4
X_8084_ _0260_ clknet_leaf_109_i_clk core_0.execute.rf.reg_outputs\[5\]\[7\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_2
X_5296_ _1731_ _1737_ _1744_ _1745_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_227_756 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7292__A1 net75 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_226_244 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7035_ _3202_ _3248_ _1366_ _3249_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4247_ net65 core_0.fetch.out_buffer_data_instr\[5\] _0725_ _0866_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_227_789 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_242_726 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_226_288 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_198_107 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5842__A2 _1444_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4178_ core_0.ew_submit _0757_ _0765_ _0796_ _0797_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai22_2
XFILLER_0_93_61 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7044__A1 _1592_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_96_116 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_179_343 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_210_601 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7595__A2 _3673_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7937_ _0115_ clknet_leaf_41_i_clk core_0.execute.sreg_priv_control.o_d\[9\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_26_826 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_195_836 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_89_190 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_77_352 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_210_667 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_93_823 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7868_ _0060_ clknet_leaf_63_i_clk core_0.fetch.prev_request_pc\[11\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_37_216 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_46_1064 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_37_249 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6819_ _2940_ _3086_ _3088_ _0301_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_107_104 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6721__B _3031_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7799_ _3861_ _3862_ _3863_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_135_424 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_18_452 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_163_744 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_282 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_73_591 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_122_107 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6307__B1 _2690_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_213_3067 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_103_310 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6858__A1 _2946_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_104_855 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5905__I0 _1721_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_103_343 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4333__A2 core_0.fetch.prev_request_pc\[6\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_131_2088 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7271__C _1735_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7807__B1 _3866_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_57_1193 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_228_34 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6168__B _1456_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_218_767 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7283__A1 _1414_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6086__A2 _2466_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7283__B2 _1431_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_205_406 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_6_584 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5833__A2 _2209_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_109_1824 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_232_247 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_224_3196 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_213_472 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87_127 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_244_66 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_69_842 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_244_77 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_200_100 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5597__A1 _1479_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_158_527 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5061__A3 _0602_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_196_2859 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_95_160 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_96_683 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_138_251 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_28_249 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_56_558 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_83_333 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_83_344 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4930__I _1393_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6010__A2 _2268_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8276__CLK clknet_leaf_26_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_37_772 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_154_766 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_24_411 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_71_539 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_399 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_126_468 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_107_660 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_141_405 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_19_i_clk_I clknet_4_8__leaf_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_153_276 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4572__A2 net157 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_444 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_839 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_3_338 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6849__A1 _2994_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_106_181 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7510__A2 _3641_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_110_803 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_122_663 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_149_2305 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_208_200 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_20_683 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5150_ _1467_ net202 _1598_ _1599_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_4
XFILLER_0_236_520 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6078__B _1480_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_138_34 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7274__A1 net87 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4101_ net71 _0721_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_3
X_5081_ _1526_ _1527_ _1528_ _1529_ _1530_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_0_236_575 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_47_65 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_223_203 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_236_597 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_224_737 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4032_ _0658_ _0659_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__inv_1
XANTENNA__6806__B _3072_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7026__A1 _1620_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_2_34 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7577__A2 _3682_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_84_1518 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_204_483 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_204_494 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_78_149 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5588__A1 _1711_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_177_836 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5983_ _2373_ _2374_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_0_63_86 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_59_352 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_63_97 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_177_858 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7722_ _3812_ _0480_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_86_160 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4934_ core_0.execute.sreg_data_page _1394_ _1397_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__7329__A2 _2265_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_192_839 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_19_238 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7653_ _3758_ _3759_ _0464_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_157_571 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_90_804 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4865_ _0843_ core_0.decode.i_imm_pass\[8\] _1305_ _1346_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_28_750 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6604_ core_0.execute.rf.reg_outputs\[7\]\[2\] _2941_ _1978_ _2952_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_15_400 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7584_ _3676_ _3702_ _3703_ _3704_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_62_539 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_145_766 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4796_ core_0.fetch.prev_request_pc\[15\] net225 _0880_ net167 _1303_ vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_0_27_282 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_15_422 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_7_677 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_105_619 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_31_884 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6535_ _2908_ _0197_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_7_699 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_104_107 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_144_276 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_241 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_132_438 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_179_30 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_70_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_95_1647 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6466_ _1059_ _1993_ _2845_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_70_594 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_95_1658 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7501__A2 _3641_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_179_85 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8205_ _0381_ clknet_leaf_2_i_clk core_0.execute.alu_mul_div.div_res\[14\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__7372__B _1395_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5512__A1 _1841_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5417_ _1857_ _1858_ _1822_ _1859_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
Xoutput130 net130 o_mem_addr[8] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_100_313 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_112_173 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_113_696 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput141 net141 o_mem_data[11] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
X_6397_ core_0.execute.alu_mul_div.mul_res\[12\] _2778_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__inv_2
XANTENNA_clkbuf_4_12__f_i_clk_I clknet_3_6_0_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput152 net152 o_mem_data[7] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_101_858 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xoutput163 net163 o_req_addr[11] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_11_672 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput174 net174 o_req_addr[7] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
X_8136_ _0312_ clknet_leaf_103_i_clk core_0.execute.rf.reg_outputs\[2\]\[11\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_10_160 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5348_ core_0.execute.alu_mul_div.div_cur\[11\] _1752_ _1788_ _1792_ _1795_ _1796_
+ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XANTENNA_input42_I i_req_data[13] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput185 net185 sr_bus_addr[1] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
Xoutput196 net196 sr_bus_data_o[11] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA__7265__A1 _3409_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_100_379 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8067_ _0243_ clknet_leaf_111_i_clk core_0.execute.rf.reg_outputs\[6\]\[6\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_2
XANTENNA__4079__A1 _0533_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5279_ _1727_ _0798_ _1432_ _1728_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_199_405 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7018_ _3189_ _3233_ _3234_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__8149__CLK clknet_leaf_107_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4174__S1 _0768_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_3_543 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6716__B _3016_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7017__A1 _1631_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_3_554 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_195_600 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_39_984 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_69_138 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_222_280 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_97_469 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_179_184 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_210_442 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_66_801 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_78_661 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_194_121 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_78_683 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_194_143 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_214_69 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_77_171 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_155_508 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_183_817 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_104_1765 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_183_839 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_19_772 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_25_219 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_837 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_93_697 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4003__A1 _0517_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_92_174 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xwire213 _0689_ net213 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_108_457 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_136_777 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_591 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_34_731 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5067__B _1459_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_20_i_clk_I clknet_4_8__leaf_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_133_2106 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5751__A1 _1683_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4554__A2 _1134_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_59_1222 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_104_641 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_61_594 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_0_308 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_238_807 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5503__A1 _1908_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_131_482 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5581__I _1983_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_239_66 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_115_1894 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_246_840 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_226_3225 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_218_531 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7256__A1 _3384_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_218_597 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_206_737 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_108_26 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_233_534 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_144_2235 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4865__I0 _0843_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_144_2246 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5530__B _1217_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_205_269 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4085__A4 core_0.execute.rf.reg_outputs\[2\]\[1\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4490__A1 core_0.decode.i_instr_l\[6\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_88_447 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_201_442 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_159_858 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_185_121 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5034__A3 core_0.dec_l_reg_sel\[0\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4242__A1 _0851_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_186_677 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_694 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_185_154 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_237_3354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5990__A1 _2123_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_84_664 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_173_338 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5990__B2 _1721_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4650_ core_0.dec_sreg_store _1209_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_126_243 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6080__C _1600_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput10 i_core_int_sreg[3] net10 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
Xinput21 i_mem_data[0] net21 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_3_102 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5742__A1 _1558_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_141_202 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_155_2375 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_4581_ _1155_ net149 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput32 i_mem_data[5] net32 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput43 i_req_data[14] net43 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xinput54 i_req_data[24] net54 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_109_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_135 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_403 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6320_ _2287_ _2056_ _2058_ _1690_ _2702_ _2703_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai221_2
XFILLER_0_142_769 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput65 i_req_data[5] net65 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_6251_ _1107_ _2634_ _2635_ _2636_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_228_317 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5202_ net95 _1446_ _1651_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_0_149_66 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_0_864 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6182_ core_0.execute.alu_mul_div.div_res\[6\] _1114_ _2566_ _2568_ _1432_ _2569_
+ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_0_149_88 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7247__A1 _1430_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_110_699 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5133_ core_0.execute.rf.reg_outputs\[7\]\[9\] net232 _1443_ core_0.execute.rf.reg_outputs\[3\]\[9\]
+ _1582_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_TAPCELL_ROW_90_1588 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_5064_ _1466_ net191 _1513_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_0_74_41 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_52 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5273__A3 _1721_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4015_ _0567_ core_0.execute.rf.reg_outputs\[3\]\[7\] _0548_ _0643_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_2
XTAP_TAPCELL_ROW_0_502 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_0_513 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4481__A1 _1066_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_220_751 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_36_943 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_177_644 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_220_762 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_9_Left_256 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_47_300 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5966_ _2271_ _2342_ _2354_ _2357_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_0_192_614 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_165_828 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7705_ _3800_ _3803_ _1284_ _0472_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_177_699 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_191_102 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4917_ _1380_ _1381_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XTAP_TAPCELL_ROW_43_1023 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_75_664 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_43_1034 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_5897_ _1456_ _2288_ _1652_ _2289_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_192_658 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_601 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_118_755 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7636_ core_0.execute.pc_high_buff_out\[4\] _3731_ _1216_ _3748_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_191_146 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_174 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_75_697 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_191_157 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_145_552 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4848_ core_0.decode.i_imm_pass\[0\] _1307_ _1337_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_28_580 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_28_591 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_118_788 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_416 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_160_500 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_172_371 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7567_ core_0.execute.pc_high_out\[1\] core_0.execute.pc_high_out\[0\] core_0.execute.pc_high_out\[2\]
+ _3689_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__5733__A1 _2113_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4536__A2 _1053_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_117_287 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4779_ core_0.fetch.prev_request_pc\[7\] _1285_ _0881_ net174 _1294_ vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_0_43_550 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5584__I1 net159 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_82 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6518_ _2447_ _2894_ _2895_ _2896_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_15_274 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_210_3037 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_120_408 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7498_ _0720_ _3640_ _3642_ _0426_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_70_391 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7486__A1 net106 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6449_ _2447_ _2827_ _2828_ _2829_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_113_482 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_8_613 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_101_644 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_101_655 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7238__A1 _1742_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_54_1163 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_8119_ _0295_ clknet_leaf_103_i_clk core_0.execute.rf.reg_outputs\[3\]\[10\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_101_699 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7789__A2 _3786_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_227_383 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_243_854 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_203_718 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_230_515 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_242_375 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_221_3166 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_199_279 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_202_239 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_98_778 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_85_406 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_195_430 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7410__A1 _1357_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6213__A2 _1758_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6960__I core_0.execute.alu_mul_div.mul_res\[1\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_195_452 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_211_784 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_168_699 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_210_294 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_195_496 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4775__A2 _1285_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_193_2829 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6181__B _0798_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5972__A1 _1059_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_182_113 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_65_1292 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_183_647 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_108_210 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_163 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_81_612 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_182_135 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_314 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_164_861 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_182_168 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7713__A2 _1064_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_81_656 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5724__A1 _1819_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4527__A2 _1053_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_117_1912 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_151_533 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_80_177 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_232_3295 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_80_188 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_34_594 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_110_49 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_111_408 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_123_279 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8314__CLK clknet_leaf_76_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6524__I0 _0553_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_104_482 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_0_138 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xclkbuf_leaf_2_i_clk clknet_4_0__leaf_i_clk clknet_leaf_2_i_clk vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_131_290 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_237_125 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7229__A1 net81 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_28_34 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_28_45 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_218_372 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_119_69 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_233_331 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_234_865 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5255__A3 _1517_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4463__A1 _1041_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_178_408 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_199_780 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_88_244 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_88_277 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7401__A1 _3563_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_159_644 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5820_ _2202_ _2216_ _2217_ _0172_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_159_655 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4215__A1 _0823_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_33_913 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_215_90 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5751_ _1683_ _1637_ _2152_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__4766__A2 _1285_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_56_141 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_146_338 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_226_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_60_32 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_174_658 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4702_ core_0.fetch.out_buffer_data_instr\[8\] net68 _1246_ _1249_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_72_612 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_174_669 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_84_483 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_56_185 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_494 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5682_ _2074_ _2075_ _2082_ _2083_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA__6507__A3 _2884_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_115_714 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7704__A2 _3788_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_13_670 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_60_98 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_807 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_142_511 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7421_ _1283_ _3581_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_44_358 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_72_667 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4518__A2 _1053_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4633_ _1173_ core_0.execute.alu_flag_reg.o_d\[3\] _1181_ _1192_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_0_25_550 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_154_382 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_4_444 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_115_769 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7352_ core_0.execute.alu_flag_reg.o_d\[3\] _3510_ _3522_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__or2_1
X_4564_ _0727_ _1144_ _1145_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__5191__A2 _1624_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_30 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_69_41 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_40_531 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6303_ _1114_ _2686_ _2687_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__7468__A1 _3581_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_12_244 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_92_1617 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_123_780 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_7283_ _1414_ core_0.execute.sreg_irq_pc.o_d\[11\] _1420_ _1431_ _1736_ _3461_ vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi221_2
X_4495_ _1087_ _0010_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_69_96 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6234_ _2447_ _2617_ _2618_ _2619_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_40_597 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_168_2533 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6691__A2 _3006_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6165_ _2465_ _2016_ _2029_ _2552_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__7142__S _1372_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_85_62 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_209_372 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_237_692 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5116_ core_0.execute.rf.reg_outputs\[1\]\[11\] net218 _1486_ core_0.execute.rf.reg_outputs\[5\]\[11\]
+ core_0.execute.rf.reg_outputs\[6\]\[11\] _1435_ _1565_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi222_2
XFILLER_0_176_97 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6096_ _2346_ net204 _2484_ _2485_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_33_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7640__A1 core_0.execute.pc_high_buff_out\[5\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4049__A4 core_0.execute.rf.reg_outputs\[2\]\[4\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
X_5047_ core_0.execute.rf.reg_outputs\[1\]\[12\] net218 _1496_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_79_222 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4454__A1 _1046_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_169_419 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_67_417 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_177_430 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_95_748 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6998_ _2001_ _2005_ _1929_ _1665_ core_0.execute.alu_mul_div.cbit\[0\] _1228_ _3215_
+ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux4_2
XTAP_TAPCELL_ROW_179_2662 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_94_247 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_138_839 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_149_176 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_164_102 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_192_422 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_101_1724 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_5949_ core_0.dec_sreg_irt _2340_ _2341_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_48_675 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_137_338 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_483 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_192_466 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_118_552 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_192_488 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_122 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_714 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_145_360 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_62_144 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7619_ net194 _3733_ _3734_ _3735_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__5706__A1 _1123_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_7_282 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3980__A3 _0544_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_133_533 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_161_842 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_62_177 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7171__A3 _1364_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_106_769 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_16_594 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_177_Right_177 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_31_531 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_105_279 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7459__A1 _3563_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_31_542 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_31_553 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_114_791 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6131__A1 _1831_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output73_I net73 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_112_1853 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4142__B1 _0549_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6682__A2 _2999_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_234_117 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_234_128 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_128_2049 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_236_34 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_216_865 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5080__B _1460_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7631__A1 net203 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_203_515 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_141_2205 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_187_205 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_242_183 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_187_216 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_67_1321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_205_2972 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_187_227 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4996__A2 core_0.dec_l_reg_sel\[1\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6904__B _3124_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_428 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_86_737 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_98_597 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6198__A1 _1378_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_168_452 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4748__A2 _1241_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_195_282 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_14_69 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_183_422 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_123_1993 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_128_349 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_156_658 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_234_3324 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_38_174 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4143__C _0534_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_139_2178 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_42_807 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_54_667 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__7698__A1 _1055_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5158__C1 _1606_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_124_522 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_306 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_170_149 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_152_2334 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_41_339 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5173__A2 _1613_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6370__A1 _2749_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_151_352 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_78_1450 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_34_391 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_144_Right_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_111_238 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_22_575 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_22_597 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4280_ core_0.fetch.prev_request_pc\[13\] _0830_ _0886_ core_0.fetch.prev_request_pc\[14\]
+ _0898_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai22_1
XTAP_TAPCELL_ROW_245_3453 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4684__A1 net38 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_207_854 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_146_34 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_176_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4385__I net86 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7622__A1 _0736_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7970_ _0147_ clknet_leaf_40_i_clk core_0.execute.mem_stage_pc\[5\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_163_2463 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_163_2474 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_222_835 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_206_397 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6921_ net92 _3135_ _3139_ _3146_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_178_216 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4987__A2 _0778_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_77_726 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6189__A1 _2202_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_76_214 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6852_ core_0.ew_reg_ie\[1\] _2934_ _3106_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_0_187_772 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_76_258 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5803_ _2201_ _2202_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_174_411 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_159_496 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4739__A2 _1238_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6783_ _2946_ _3064_ _3067_ _0286_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_3995_ net103 _0578_ _0625_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_45_612 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_147_658 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_44_100 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5734_ _1698_ _2134_ _2135_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_162_606 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_280 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_99_Left_346 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
Xclkbuf_leaf_103_i_clk clknet_4_5__leaf_i_clk clknet_leaf_103_i_clk vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_146_168 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_174_477 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_45_656 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_431 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_115_500 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_134_319 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7689__A1 _3786_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_60_604 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5665_ _2063_ _2065_ _2066_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__3962__A3 _0518_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_143_842 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_44_177 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7404_ _1980_ _3567_ _0407_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__6041__S _1482_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4616_ core_0.dec_jump_cond_code\[1\] _1175_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA_clkbuf_leaf_67_i_clk_I clknet_4_15__leaf_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6361__A1 _1686_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5596_ _1765_ _1665_ _1997_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_0_25_380 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6361__B2 _1752_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_130_514 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_103_739 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_111_Right_111 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
X_7335_ net194 _3495_ _3507_ _3496_ _3508_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__4911__A2 _1231_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4547_ _1130_ _0003_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xclkbuf_leaf_118_i_clk clknet_4_6__leaf_i_clk clknet_leaf_118_i_clk vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_102_238 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_130_569 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7266_ _3442_ _3446_ _1395_ _0390_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_111_772 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4478_ _1038_ _1039_ _1071_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_0_96_72 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6217_ _2602_ _2498_ _2102_ _2603_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__6664__A2 _2934_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_217_629 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_229_489 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7197_ _3382_ _3383_ _3384_ _3385_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_244_426 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4675__A1 _1227_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_51_1122 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6148_ core_0.execute.pc_high_buff_out\[6\] _2249_ _2534_ net13 _2535_ vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__7613__A1 _1209_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_213_813 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6079_ net223 _1597_ _2468_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_224_161 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4427__A1 _0883_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_169_205 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_240_632 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_206_37 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4978__A2 _0553_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_726 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_737 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6216__S _1625_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_178_750 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_240_698 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_68_759 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_246_Right_246 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_49_1095 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5927__A1 _2300_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_165_422 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_177_282 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_36_623 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_483 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_62_1251 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_82_228 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_222_69 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_62_1262 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_165_488 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_24_798 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_24_807 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_63_464 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_118_382 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_91_784 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_23_328 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6352__A1 _2626_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50_125 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5155__A2 _0767_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_133_352 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_51_659 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_90_294 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_16_391 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_133_385 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4902__A2 _1231_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_121_558 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5790__S _2190_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6104__A1 net83 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6104__B2 _2245_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6655__A2 core_0.ew_data\[13\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_82_i_clk clknet_4_13__leaf_i_clk clknet_leaf_82_i_clk vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_TAPCELL_ROW_73_1391 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6407__A2 _2579_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7604__A1 _3663_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4418__A1 net80 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_243_492 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_231_632 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_116_26 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_215_194 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_97_i_clk clknet_4_7__leaf_i_clk clknet_leaf_97_i_clk vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_98_350 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4969__A2 _0592_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_240_3394 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5091__A1 net93 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_203_367 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_86_523 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_98_383 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_169_750 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_58_247 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_213_Right_213 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_58_269 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_20_i_clk clknet_4_8__leaf_i_clk clknet_leaf_20_i_clk vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_168_282 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_184_731 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6040__B1 _1999_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_144_617 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_183_263 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7465__B _3540_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_143_127 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_125_842 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_26_177 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xclkbuf_leaf_35_i_clk clknet_4_11__leaf_i_clk clknet_leaf_35_i_clk vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_5450_ _1374_ _1880_ _1887_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__6343__A1 _2346_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5146__A2 _1557_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_112_503 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_42_659 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_112_514 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4401_ _0948_ _0949_ _1009_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__6894__A2 _3129_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5381_ _1233_ _1818_ _1827_ _1822_ _1828_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_239_710 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7120_ _3326_ _3327_ _3328_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4332_ _0903_ _0909_ _0948_ _0949_ _0950_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_0_10_523 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_239_765 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6646__A2 core_0.ew_data\[10\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7051_ _1224_ _3215_ _1222_ _3264_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_4263_ _0881_ net177 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XANTENNA__4657__A1 _1172_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8032__CLK clknet_leaf_53_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6002_ _2346_ net221 _2392_ _2393_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_4194_ core_0.decode.input_valid _0812_ _0813_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_0_66_86 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4409__A1 _0835_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_173_10 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7953_ _0131_ clknet_leaf_4_i_clk core_0.execute.alu_mul_div.div_cur\[9\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_221_142 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6904_ net99 _3135_ _3124_ _3137_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_7884_ _0075_ clknet_leaf_51_i_clk core_0.decode.i_instr_l\[9\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_65_707 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_159_271 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5909__A1 _1559_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6835_ core_0.execute.rf.reg_outputs\[2\]\[8\] _3092_ _3083_ _3097_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_9_322 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_159_282 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_176_2621 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_77_589 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_147_433 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_119_135 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_175_753 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6766_ _1963_ _3057_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA__6582__A1 net155 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3978_ _0534_ _0535_ _0536_ core_0.execute.rf.reg_outputs\[6\]\[10\] _0609_ vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_0_135_628 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_656 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_175_797 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_190_734 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_18_667 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5717_ _2116_ _2117_ _1554_ _2118_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_73_762 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_45_464 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_18_678 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3935__A3 _0549_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6697_ _2992_ _3000_ _3017_ _0250_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_45_486 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_21_768 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_115_330 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_72_283 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6334__A1 _2360_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5137__A2 _1438_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5648_ _2036_ _2038_ _2048_ _2049_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_98_1689 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6885__A2 _3108_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_103_547 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5579_ _1982_ _0166_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4896__A1 _0804_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7318_ _3409_ _3488_ _3489_ _3491_ _3492_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai22_2
XFILLER_0_229_220 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8298_ _0474_ clknet_leaf_48_i_clk core_0.dec_mem_access vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__dffq_2
X_7249_ _3409_ _3431_ _3432_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_187_2761 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output159_I net159 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_229_286 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_204_109 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_125_2008 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_99_114 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_225_492 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_213_632 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7062__A2 _1585_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_29_857 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5073__A1 net94 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_240_451 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_202_2931 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_240_473 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_240_484 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_202_2942 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_68_556 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_96_865 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_107_1796 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_218_3127 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_198_2890 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_166_753 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_120_1952 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_55_239 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5376__A2 _1814_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_125_116 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_107_842 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3926__A3 _0544_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_136_2148 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_23_103 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_497 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6325__A1 _2123_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5128__A2 _1576_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_106_352 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_456 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6876__A2 _3107_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8055__CLK clknet_leaf_104_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_31_180 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_20_865 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6629__B _1978_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_229_3256 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5533__B _1217_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6628__A2 core_0.ew_data\[6\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4639__A1 net185 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_235_212 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_242_3412 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_36_34 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_147_2277 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
Xinput8 i_core_int_sreg[1] net8 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_clkbuf_leaf_15_i_clk_I clknet_4_8__leaf_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_216_481 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_189_834 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_78_309 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_160_2433 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_188_333 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_203_142 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5064__A1 _1466_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_188_355 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4950_ core_0.execute.sreg_priv_control.o_d\[6\] _1394_ _1408_ _1391_ _1409_ vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__6800__A2 _3070_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4811__A1 core_0.decode.i_instr_l\[4\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3901_ _0534_ _0535_ _0536_ core_0.execute.rf.reg_outputs\[6\]\[15\] _0537_ vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_0_19_409 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_129_422 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4881_ _0827_ _1321_ _1354_ _0097_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__5695__S _1554_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_139_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6620_ net32 _1149_ _2965_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_46_239 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_129_466 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_156_263 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_6_314 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7195__B _1736_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6551_ _2916_ _0205_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_61_209 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_144_436 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_172_745 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_6_347 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_27_486 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5502_ _1908_ _1934_ _1935_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_144_469 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_172_778 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_15_648 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_70_732 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_592 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6482_ core_0.execute.sreg_priv_control.o_d\[14\] _1386_ _2577_ core_0.execute.sreg_irq_pc.o_d\[14\]
+ _2861_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_42_434 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_171_2562 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_8221_ _0397_ clknet_leaf_35_i_clk net78 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_4
XANTENNA__6867__A2 _3114_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5433_ _1790_ _1788_ _1872_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_112_333 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_140_642 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4878__A1 core_0.decode.i_imm_pass\[14\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_8152_ _0328_ clknet_leaf_102_i_clk core_0.execute.rf.reg_outputs\[1\]\[11\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5364_ _1811_ _1812_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_22_191 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_597 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_239_562 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_227_702 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7103_ _1222_ _3216_ _3312_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_112_399 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4315_ _0917_ _0928_ _0930_ _0932_ _0933_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or4_2
XANTENNA__7816__A1 _1098_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_8083_ _0259_ clknet_leaf_114_i_clk core_0.execute.rf.reg_outputs\[5\]\[6\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_77_74 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_10_375 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5295_ _1741_ _1743_ _0731_ _1744_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_168_98 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_226_234 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7034_ _3245_ _3247_ _1229_ _3248_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__7292__A2 _3398_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4246_ net66 core_0.fetch.out_buffer_data_instr\[6\] _0724_ _0865_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_227_768 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_199_609 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_214_418 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_93_40 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_93_51 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4177_ _0766_ _0795_ _0796_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_207_492 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_179_311 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_182_2691 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7044__A2 _3209_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_97_629 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5055__A1 _0630_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4573__I _1151_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_96_128 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7936_ _0114_ clknet_leaf_34_i_clk core_0.execute.sreg_priv_control.o_d\[8\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_139_208 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_222_495 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_26_827 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_77_342 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_78_865 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_194_325 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_195_859 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7867_ _0059_ clknet_leaf_59_i_clk core_0.fetch.prev_request_pc\[10\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_46_1065 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_182_509 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_77_397 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_606 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6818_ core_0.execute.rf.reg_outputs\[2\]\[0\] _3087_ _3083_ _3088_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__5358__A2 _1713_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_148_786 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_65_559 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7798_ _1120_ _3838_ _3859_ _3862_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_135_414 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_190_520 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_196 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_138 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6749_ core_0.execute.rf.reg_outputs\[4\]\[3\] _3043_ _3045_ _3048_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__4522__B _1078_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_45_261 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_570 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_162_255 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6307__B2 _2360_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_61_754 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_213_3068 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_190_597 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_116_683 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_150_439 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6858__A2 _3107_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_489 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_60_297 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4333__A3 _0950_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5530__A2 _1957_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_131_697 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_103_399 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_131_2089 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_218_713 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7807__A1 core_0.decode.i_instr_l\[15\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_57_1194 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7807__B2 core_0.decode.i_instr_l\[12\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_217_212 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7915__CLK clknet_leaf_119_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_217_256 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_70_1350 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_245_576 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5294__A1 net72 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_205_418 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_6_585 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_189_108 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_109_1825 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_224_3197 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_232_259 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_198_642 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_201_602 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_201_613 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5597__A2 _1931_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_84_802 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_96_662 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_201_668 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_138_241 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_239 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_113_38 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5349__A2 _1528_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_43_209 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_81_1490 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_154_745 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_126_447 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_153_244 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_4_807 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_24_423 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_153_255 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_107_672 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_694 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_52_787 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6849__A2 _3087_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_117 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_51_297 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_139 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5521__A2 _0807_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_149_2306 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_209_702 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4658__I _0722_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_47_22 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4100_ _0720_ net194 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__inv_4
XFILLER_0_236_543 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5080_ _0570_ _0575_ _1460_ _0579_ _1529_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai211_4
XFILLER_0_236_565 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5285__A1 _1195_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6482__B1 _2577_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4031_ net100 _0577_ _0658_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__7026__A2 _3178_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_189_642 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_79_629 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_154_34 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_204_451 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_204_Left_451 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__5037__A1 _0782_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_189_664 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_204_473 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_84_1519 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_188_152 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6785__A1 _2951_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5982_ _1623_ _1594_ _1558_ _2373_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__5588__A2 _1719_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_63_76 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_149_528 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_231_292 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_188_174 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_176_325 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4933_ _1396_ _0107_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_7721_ net189 core_0.decode.i_imm_pass\[5\] _1946_ _3812_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_192_807 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6822__B _3083_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_47_526 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_75_835 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_86_172 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_129_230 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4864_ _0833_ _1321_ _1345_ _0089_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_7652_ core_0.dec_mem_long _1032_ _1217_ _3759_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_6603_ _2930_ core_0.ew_data\[2\] _2950_ _2951_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_4
XANTENNA__5438__B _1841_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7583_ core_0.execute.pc_high_out\[4\] _3695_ _3703_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or2_1
X_4795_ _1301_ _1302_ _0063_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_7_656 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4012__A2 core_0.execute.rf.reg_outputs\[4\]\[7\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_15_412 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_55_581 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6534_ net124 _2440_ _2906_ _2908_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_144_266 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_31_885 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_6_177 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_160_737 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_213_Left_460 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_43_776 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_125_480 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6465_ _2090_ _2843_ _1699_ _2844_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_179_53 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_489 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_95_1648 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_42_297 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8204_ _0380_ clknet_leaf_1_i_clk core_0.execute.alu_mul_div.div_res\[13\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_101_815 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5416_ _1233_ _1850_ _1858_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xoutput120 net120 o_mem_addr[13] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_30_448 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput131 net131 o_mem_addr[9] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
X_6396_ _2765_ _2768_ _2776_ _2777_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_4
XANTENNA__5512__A2 _1719_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput142 net142 o_mem_data[12] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_63_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xoutput153 net153 o_mem_data[8] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
X_8135_ _0311_ clknet_leaf_104_i_clk core_0.execute.rf.reg_outputs\[2\]\[10\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xoutput164 net164 o_req_addr[12] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
X_5347_ _1793_ _1794_ _1795_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
Xoutput175 net175 o_req_addr[8] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_227_510 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_684 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput186 net186 sr_bus_addr[2] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_239_381 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput197 net197 sr_bus_data_o[12] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XTAP_TAPCELL_ROW_184_2720 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_8066_ _0242_ clknet_leaf_112_i_clk core_0.execute.rf.reg_outputs\[6\]\[5\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_10_194 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5278_ core_0.execute.alu_mul_div.div_res\[0\] _1727_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__4079__A2 _0541_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5276__A1 core_0.execute.alu_mul_div.i_mul vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input35_I i_mem_data[8] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_215_727 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7017_ _1631_ _3209_ _3231_ _3232_ _3233_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_4229_ _0842_ _0843_ _0844_ _0847_ _0848_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor4_2
XFILLER_0_242_524 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_214_215 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_3_544 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7017__A2 _3209_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5028__A1 _1457_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_168_804 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_39_985 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6776__A1 _2996_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_214_37 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_210_454 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7919_ _0010_ clknet_4_3__leaf_i_clk core_0.decode.oc_alu_mode\[7\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_194_133 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_104_1755 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_104_1766 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_77_183 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_183_829 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6528__A1 _1729_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_182_317 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_194_177 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_92_131 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_135_200 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_148_594 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_182_339 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_25_209 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_108_447 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xwire214 _1540_ net214 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_18_283 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_133_2107 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_163_586 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5751__A2 _1637_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_61_562 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_59_1223 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5503__A2 _1613_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_237_318 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_103_185 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_115_1895 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_218_521 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_226_3226 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5267__A1 _1714_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_233_524 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_205_226 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_205_237 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_108_49 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_144_2236 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_233_557 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4427__B _1029_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_88_415 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5019__A1 net88 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4490__A2 core_0.decode.i_instr_l\[4\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_198_450 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_220_229 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_213_270 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_640 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8243__CLK clknet_leaf_43_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_198_483 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_124_37 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_161 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_174_807 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4242__A2 _0854_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_186_689 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_237_3355 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6519__A1 net78 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_29_559 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_127_712 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6519__B2 _2537_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_83_142 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_204_81 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_EDGE_ROW_62_Left_309 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_83_175 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_127_767 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_182_862 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_37_592 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_197 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xinput11 i_core_int_sreg[4] net11 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_114_406 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput22 i_mem_data[10] net22 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_4580_ core_0.ew_data\[4\] net157 _1155_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_TAPCELL_ROW_155_2376 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5742__A2 _1652_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_142_737 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_154_597 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xinput33 i_mem_data[6] net33 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput44 i_req_data[15] net44 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xinput55 i_req_data[25] net55 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput66 i_req_data[6] net66 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_24_286 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_40_746 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_122_450 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_448 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6250_ _2047_ _2161_ _2635_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6542__I1 _2611_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5201_ core_0.execute.rf.reg_outputs\[2\]\[1\] _1438_ _1648_ _0769_ _1649_ _1650_
+ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi221_4
X_6181_ _1433_ _2567_ _0798_ _2568_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_110_667 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_481 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_110_678 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5132_ _0789_ core_0.execute.rf.reg_outputs\[4\]\[9\] _0779_ _1581_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XPHY_EDGE_ROW_71_Left_318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__5258__A1 _1695_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_90_1589 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_236_384 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_224_524 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5063_ _1508_ _1509_ _1510_ _1511_ _1512_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_0_224_535 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4014_ _0533_ _0523_ _0526_ core_0.execute.rf.reg_outputs\[6\]\[7\] _0642_ vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_0_224_579 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_212_719 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_0_503 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_0_514 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_79_448 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6758__A1 core_0.execute.rf.reg_outputs\[4\]\[7\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5012__I _1460_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_220_741 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_36_944 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_181_43 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_149_347 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_176_133 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5965_ core_0.dec_sreg_load core_0.dec_sreg_jal_over _2356_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_0_47_312 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_75_621 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5430__A1 _1233_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_47_323 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_183 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_632 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_87_492 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7704_ _3786_ _3788_ _3802_ _3799_ _3803_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai31_1
X_4916_ _1379_ _1380_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XPHY_EDGE_ROW_80_Left_327 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_164_317 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_176_177 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5896_ _2287_ _1603_ _2288_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_118_723 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_158_Right_158 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_43_1024 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_47_367 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3992__A1 _0565_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_118_745 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_145_531 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7635_ net204 _3733_ _3746_ _3747_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__7183__A1 _2714_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4847_ _1334_ _1336_ _0081_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_173_862 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_117_255 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_145_564 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_145_575 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4778_ _1290_ _1293_ _0055_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_7566_ core_0.execute.pc_high_out\[2\] core_0.execute.pc_high_out\[1\] core_0.execute.pc_high_out\[0\]
+ _3688_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and3_1
XANTENNA__5733__A2 _2122_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6930__A1 _1221_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_145_597 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_702 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_43_562 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7383__B _3546_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_132_247 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6517_ core_0.execute.sreg_priv_control.o_d\[15\] _1386_ _2577_ core_0.execute.sreg_irq_pc.o_d\[15\]
+ _2895_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_TAPCELL_ROW_210_3027 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_190_2790 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_210_3038 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_30_212 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7497_ core_0.execute.sreg_scratch.o_d\[0\] _3641_ _3516_ _3642_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_31_757 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6448_ core_0.execute.sreg_priv_control.o_d\[13\] _1386_ _2577_ core_0.execute.sreg_irq_pc.o_d\[13\]
+ _2828_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_TAPCELL_ROW_8_603 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_100_100 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_8_614 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_246_104 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_267 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_30_278 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6379_ _2244_ _2760_ _2761_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_100_155 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_11_492 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8118_ _0294_ clknet_leaf_108_i_clk core_0.execute.rf.reg_outputs\[3\]\[9\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_54_1164 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_100_177 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5249__A1 _1695_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6727__B _3031_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_215_513 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8049_ _0225_ clknet_leaf_114_i_clk core_0.execute.rf.reg_outputs\[7\]\[4\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_215_546 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_221_3167 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_225_58 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_225_69 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_119_Left_366 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_167_122 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_168_645 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_156_807 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_168_667 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_210_251 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5421__A1 _1374_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_128_509 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_195_464 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4761__I _1051_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_155_306 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_183_626 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_131 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_155_328 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_125_Right_125 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_65_1293 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5078__B _1461_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3983__A1 net89 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_136_531 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_80_101 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7174__A1 _3261_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_93_484 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_108_233 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5185__B1 _1436_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_136_586 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_136_597 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6921__A1 net92 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_117_1913 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4932__B1 _1394_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_584 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_232_3296 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_21_201 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_21_212 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_104_450 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1_629 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_128_Left_375 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_104_472 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_132_781 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7721__I0 net189 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5488__A1 _1230_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_104_494 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_237_137 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_790 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_246_682 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_218_384 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_206_524 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_233_343 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4999__B1 _1443_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_88_201 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_233_376 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4463__A2 _1048_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_233_387 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_34 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_89_757 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_137_Left_384 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_89_768 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_202_741 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7401__A2 net81 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_44_89 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_159_667 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4215__A2 _0827_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_33_903 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_33_914 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_57_632 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4671__I _1226_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_492 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5750_ _1715_ _1631_ _2151_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_29_345 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_146_317 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_158_177 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_228 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4701_ _1248_ _0023_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_173_136 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5681_ _2079_ _2081_ _2082_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__7165__A1 _1369_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_121_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_219_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_71_123 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7704__A3 _3802_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_154_350 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7420_ _1980_ _3580_ _0410_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_4632_ core_0.dec_jump_cond_code\[3\] _1190_ _1191_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_13_671 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_115_726 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_154_372 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_182_681 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5715__A2 _2092_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6912__A1 _2981_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_142_523 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_702 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_25_573 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_34 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_114_236 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_71_189 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7351_ net213 _3502_ _3518_ _3520_ _3510_ _3521_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai221_2
XFILLER_0_114_247 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_EDGE_ROW_146_Left_393 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_170_865 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4563_ core_0.fetch.prev_req_branch_pred _1144_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_142_567 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_130_718 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6302_ _2281_ _2684_ _2685_ _2686_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_7282_ _2752_ _3391_ _3460_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4494_ _1061_ _1062_ _1064_ _1086_ _1087_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_TAPCELL_ROW_92_1618 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_229_616 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5479__A1 _1909_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6233_ core_0.execute.sreg_priv_control.o_d\[8\] _1386_ _2577_ core_0.execute.sreg_irq_pc.o_d\[8\]
+ _2618_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_100_72 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_168_2523 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_229_649 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_168_2534 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_110_464 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6164_ core_0.decode.oc_alu_mode\[4\] _2550_ _2551_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5115_ core_0.execute.rf.reg_outputs\[7\]\[11\] net232 _1443_ core_0.execute.rf.reg_outputs\[3\]\[11\]
+ _1564_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_6095_ _2458_ _2483_ core_0.dec_mem_access _2484_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_236_192 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_227_Right_227 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
X_5046_ _1493_ _1494_ _1495_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__7640__A2 _3731_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_26_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_79_212 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4454__A2 _1048_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_63_i_clk_I clknet_4_15__leaf_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_224_387 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_212_527 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_212_538 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_149_133 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_94_215 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_138_807 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6997_ _3198_ _3205_ _3213_ _3214_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XANTENNA__5403__A1 _1375_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_179_2663 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_165_626 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5948_ net79 _2268_ _2339_ _2245_ _2340_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_47_142 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_101_1725 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_164_125 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_164_136 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7156__A1 _1369_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_62_101 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_63_624 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5879_ _2243_ _2271_ _2272_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_192_478 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_161_810 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7618_ _0739_ _3733_ _3734_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5167__B1 _1434_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_105_203 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_106_726 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5706__A2 _1676_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_106_737 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_118_597 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6903__A1 _2961_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_62_156 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_173_692 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_133_545 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output189_I net189 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7549_ _3672_ _3673_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_31_521 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4390__A1 core_0.fetch.prev_request_pc\[6\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7459__A2 net76 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_120_239 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_219_126 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6131__A2 _2516_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_112_1854 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4142__A1 core_0.ew_reg_ie\[6\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4142__B2 core_0.ew_reg_ie\[7\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_234_107 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_228_671 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4756__I _1051_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6176__C _2562_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_215_354 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_98_510 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_188_718 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_141_2206 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_203_527 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6985__A4 _3202_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_67_1311 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_231_858 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_67_1322 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_205_2973 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4996__A3 core_0.dec_l_reg_sel\[0\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_230_379 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_105_39 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7395__A1 _1357_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_14_37 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_39_632 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_120 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_128_317 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_156_626 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_123_1983 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5945__A2 _2254_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4424__C _0877_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_123_1994 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_234_3325 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_94_782 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7147__A1 _1719_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_66_484 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_109_553 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_337 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_139_2179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5158__B1 _1605_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_81_454 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_121_38 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7698__A2 _1094_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_121_49 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_10_630 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_163_180 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_152_2335 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_151_342 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_152_865 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6370__A2 _2750_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_381 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_22_521 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_78_1451 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_112_729 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4381__A1 core_0.fetch.prev_request_pc\[9\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50_863 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_716 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_280 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_34 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4867__S _1305_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_120_773 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_238_457 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_39_89 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_245_3454 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4684__A2 _1238_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5881__A1 _1729_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_206_321 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_218_192 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_163_2464 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5698__S _1554_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_206_387 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_169_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6920_ _2990_ _3130_ _3145_ _0345_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_89_1580 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_221_357 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_18_730 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6851_ _2996_ _3087_ _3105_ _0316_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_162_34 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5497__I net97 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7386__A1 _1980_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_193_209 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5802_ _1984_ _2201_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_146_103 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3994_ _0620_ _0621_ _0622_ _0623_ _0624_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_4
X_6782_ core_0.execute.rf.reg_outputs\[3\]\[1\] _3065_ _3057_ _3067_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__5936__A2 _2299_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_119_328 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_29_142 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_57_462 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_91_207 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_304 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5733_ _2113_ _2122_ _2129_ _2132_ _2133_ _2134_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XANTENNA__7138__A1 _1915_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_17_348 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_154_Left_401 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__7689__A2 _3788_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5664_ _2051_ _2054_ _2064_ _2065_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_161_139 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_44_167 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5446__B _1817_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7403_ core_0.execute.sreg_irq_pc.o_d\[3\] _3543_ _3566_ _3567_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4615_ core_0.dec_jump_cond_code\[1\] core_0.dec_jump_cond_code\[0\] core_0.execute.alu_flag_reg.o_d\[2\]
+ _1174_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_5595_ _1993_ _1995_ _1996_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_115_578 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4372__A1 _0965_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_102_206 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7334_ _2854_ _2886_ _2887_ _3506_ _3507_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor4_4
X_4546_ core_0.decode.oc_alu_mode\[13\] _1062_ _1064_ _1129_ _1130_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_102_228 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_130_537 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_229_435 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7265_ _3409_ _3445_ _3446_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__7310__A1 _0964_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4477_ _1066_ _1068_ _1069_ _1070_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_0_111_784 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6216_ _2097_ _2095_ _1625_ _2602_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_7196_ _1051_ _1392_ _3384_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_0_216_107 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_51_1123 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4675__A2 _1230_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5872__A1 net186 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6147_ _2260_ _2534_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XPHY_EDGE_ROW_163_Left_410 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_224_140 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7613__A2 _2249_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6078_ _2300_ _1560_ _1480_ _2467_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_224_151 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_240_611 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_225_696 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_224_173 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6791__I _1963_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5029_ _1467_ net187 _1478_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_213_858 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_197_526 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_200_508 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_68_749 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8304__CLK clknet_leaf_76_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_95_535 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_184_209 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output104_I net104 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_177_261 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_49_1096 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_83_708 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_165_412 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_1_i_clk clknet_4_2__leaf_i_clk clknet_leaf_1_i_clk vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__5927__A2 _1624_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_222_37 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_62_1252 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_36_635 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_153_629 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_24_799 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_51_605 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_133_320 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_216_3099 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_23_318 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_50_104 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_134_865 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_50_115 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_381 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_121_504 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6031__I _2009_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5075__C _1461_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_32_863 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7301__A1 net76 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6104__A2 _2268_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_102_773 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4115__A1 core_0.execute.pc_high_out\[2\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5863__A1 net186 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_235_438 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_207_129 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_73_1392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4419__C _0963_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_204_803 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6915__B _3139_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_231_622 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4418__A2 _0883_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_203_346 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_116_49 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_240_3395 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5091__A2 _1492_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_98_362 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_58_215 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7368__A1 core_0.execute.alu_flag_reg.o_d\[4\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_231_699 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_98_395 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_175_209 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_196_581 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5110__I _1558_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5918__A2 _2309_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6040__A1 _1665_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_129_648 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_183_220 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_129_659 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_27_613 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_132_37 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6650__B _2984_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_184_776 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_82_741 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_82_752 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_240 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_212_70 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_82_796 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_clkbuf_leaf_11_i_clk_I clknet_4_9__leaf_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6343__A2 net195 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7540__A1 _3663_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4400_ net83 _1008_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__inv_2
XANTENNA__4354__A1 _0847_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5380_ _1232_ _1826_ _1827_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_152_695 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1_212 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_112_537 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_671 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_151_194 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4331_ core_0.fetch.prev_request_pc\[2\] core_0.fetch.prev_request_pc\[1\] core_0.fetch.prev_request_pc\[0\]
+ _0949_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_4
X_7050_ _1224_ _3262_ _3263_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or2_1
X_4262_ _0880_ _0881_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_120_581 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6001_ _2359_ _2391_ _2346_ _2392_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_226_438 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_66_43 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4193_ _0754_ _0756_ _0811_ _0812_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and3_4
XFILLER_0_157_78 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_66_76 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4409__A2 _0947_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_234_493 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7952_ _0130_ clknet_leaf_4_i_clk core_0.execute.alu_mul_div.div_cur\[8\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_2
XANTENNA__5082__A2 _1525_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6903_ _2961_ _3129_ _3136_ _0337_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_82_75 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7883_ _0074_ clknet_leaf_83_i_clk core_0.decode.i_instr_l\[8\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_106_60 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_71 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_248 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_175_710 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6834_ _2977_ _3086_ _3096_ _0308_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_77_568 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5909__A2 _1689_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_15_80 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_719 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_176_2622 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_147_445 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_613 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_345 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_92_527 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7656__B _1037_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6765_ _2986_ _3043_ _3056_ _0279_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_119_158 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_175_776 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5955__I core_0.dec_mem_access vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3977_ _0605_ _0594_ _0606_ _0607_ _0608_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai211_4
XANTENNA__6582__A2 _2190_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5716_ _1124_ _1568_ _2091_ _2092_ _2117_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_0_72_240 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_251 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6696_ core_0.execute.rf.reg_outputs\[6\]\[13\] _3006_ _3016_ _3017_ vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_93_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_134_139 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_73_785 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_21_769 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_116_865 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_32_115 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5647_ _2047_ _2041_ _2048_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__6334__A2 _2716_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_5_562 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_32_137 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_60_457 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_143_684 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_142_172 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_143_695 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_863 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_479 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5578_ core_0.execute.trap_flag _0177_ _1982_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA_input65_I i_req_data[5] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_103_559 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4896__A2 _1221_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7391__B _3545_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7317_ _3409_ _3490_ _3491_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5690__I net211 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4529_ _1037_ _1090_ _1116_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_13_395 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_8297_ _0473_ clknet_leaf_46_i_clk core_0.dec_mem_we vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__6098__A1 core_0.ew_data\[4\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_187_2751 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_7248_ _2539_ _3430_ _3431_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_187_2762 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5845__A1 _2236_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4648__A2 _0731_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_244_235 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7179_ _1748_ _3374_ _0375_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_125_2009 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_213_600 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7598__A1 core_0.execute.pc_high_out\[6\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_198_802 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6735__B _3031_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_148 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6270__A1 _2346_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_212_143 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_201_806 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_29_858 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5073__A2 _0521_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_197_345 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_202_2932 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_213_699 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_157_209 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_212_187 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_95_332 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_96_855 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_95_343 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_178_570 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_107_1797 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_56_719 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_218_3128 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_198_2891 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_55_207 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_516 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_120_1953 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_181_702 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_193_562 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7770__A1 _1136_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4584__A1 core_0.ew_data\[6\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_443 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_165_286 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_36_465 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_24_627 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_136_2149 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7522__A1 _0615_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_23_126 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4336__A1 core_0.fetch.prev_request_pc\[11\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7994__CLK clknet_leaf_89_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_75_1410 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_161_492 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5814__B _2183_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_855 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6089__A1 core_0.execute.alu_mul_div.i_mul vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_236_703 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_229_3257 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_208_427 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4639__A2 net178 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_242_3413 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_236_758 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_235_224 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_235_235 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5105__I _1553_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_235_257 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_235_268 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_223_419 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_102_i_clk clknet_4_7__leaf_i_clk clknet_leaf_102_i_clk vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_TAPCELL_ROW_147_2278 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7589__A1 _3673_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput9 i_core_int_sreg[2] net9 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_243_290 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_160_2434 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_99_660 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6261__A1 _2626_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5064__A2 net191 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_203_154 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_86_1550 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_86_321 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_176_518 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_546 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_leaf_117_i_clk clknet_4_4__leaf_i_clk clknet_leaf_117_i_clk vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__4811__A2 _1307_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_47_708 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_52_34 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3900_ _0526_ _0536_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_52_45 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4880_ core_0.decode.i_imm_pass\[15\] _1341_ _1354_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_86_376 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_129_434 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_74_527 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_223_80 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7761__A1 _1038_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_184_573 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_117_629 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_129_489 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_156_275 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6550_ net117 _2752_ _2906_ _2916_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_27_454 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_6_337 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5501_ net99 _1629_ _1492_ _1934_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_6481_ core_0.execute.sreg_scratch.o_d\[14\] _2579_ _2534_ net6 _2860_ vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_0_201_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_171_2563 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_8220_ _0396_ clknet_leaf_33_i_clk net77 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_4
XANTENNA__4327__A1 _0877_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_42_457 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5432_ _1747_ _1866_ _1871_ _0131_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_0_124_172 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_140_632 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_112_345 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4878__A2 _1341_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_8151_ _0327_ clknet_leaf_102_i_clk core_0.execute.rf.reg_outputs\[1\]\[10\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5363_ _1374_ _1809_ _1810_ _1811_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_0_10_310 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_112_378 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7277__B1 _3399_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7102_ _1225_ _3309_ _3310_ _1372_ _3311_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_4314_ _0902_ _0915_ _0931_ _0932_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_77_64 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8082_ _0258_ clknet_leaf_114_i_clk core_0.execute.rf.reg_outputs\[5\]\[5\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_2
X_5294_ net72 _1742_ _1735_ _1743_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__5827__A1 net135 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_226_213 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_387 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4245_ _0820_ _0863_ _0864_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7033_ _1226_ _1613_ _3246_ _3247_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_226_257 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4176_ _0786_ _0791_ _0792_ _0771_ _0794_ _0795_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XTAP_TAPCELL_ROW_182_2692 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_184_98 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_96_107 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5055__A2 _0635_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6252__A1 _1756_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7935_ _0113_ clknet_leaf_32_i_clk core_0.execute.sreg_priv_control.o_d\[7\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_195_816 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_26_828 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_78_855 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_179_378 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_89_192 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7866_ _0058_ clknet_leaf_63_i_clk core_0.fetch.prev_request_pc\[9\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_148_732 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6004__A1 _2202_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_92_302 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_46_1066 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6817_ _3085_ _3087_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_9_142 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_93_858 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_163_702 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_175_562 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7797_ _1096_ _3778_ _3860_ _3861_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
Xclkbuf_leaf_81_i_clk clknet_4_13__leaf_i_clk clknet_leaf_81_i_clk vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_190_510 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_454 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_190_532 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6748_ _2951_ _3042_ _3047_ _0271_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__4522__C _1064_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_402 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_163_768 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_273 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_190_576 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_60_210 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_33_435 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6679_ core_0.execute.rf.reg_outputs\[6\]\[5\] _3006_ _3004_ _3008_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_61_744 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7504__A1 net212 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_115_150 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_213_3069 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_60_243 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_766 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_96_i_clk clknet_4_6__leaf_i_clk clknet_leaf_96_i_clk vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_20_107 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output171_I net171 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_131_2079 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7807__A2 _3788_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_57_1195 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_245_544 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_70_1351 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5294__A2 _1742_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_232_205 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_217_279 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_6_586 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_109_1815 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_232_227 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_109_1826 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_224_3198 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_34_i_clk clknet_4_11__leaf_i_clk clknet_leaf_34_i_clk vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_241_761 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_197_120 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6243__A1 _2026_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_241_772 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_198_654 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_100_Left_347 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_197_142 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_68_310 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_186_827 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_158_518 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_197_164 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6794__A2 _3070_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_197_197 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_185_337 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_185_348 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_387 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__7296__B _1395_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_49_i_clk clknet_4_12__leaf_i_clk clknet_leaf_49_i_clk vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__5349__A3 _1529_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_37 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_166_573 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_81_1480 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4557__A1 _1065_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_153_212 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_71_519 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_640 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_273 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_52_733 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_457 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_24_479 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_134_492 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5544__B _1964_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_121_142 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_652 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_20_685 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_208_224 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_138_69 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6482__A1 core_0.execute.sreg_priv_control.o_d\[14\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
X_4030_ _0653_ _0654_ _0655_ _0656_ _0657_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_4
XPHY_EDGE_ROW_10_Right_10 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_223_216 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5824__A4 _2215_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_223_227 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_79_608 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_79_619 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_139_Right_139 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__6234__A1 _2447_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_188_120 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_78_107 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5037__A2 _0767_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_2_69 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_231_260 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5981_ _2369_ _2371_ _2372_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_151_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6785__A2 _3064_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_63_66 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7720_ _3811_ _0479_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4796__A1 core_0.fetch.prev_request_pc\[15\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4932_ net194 _1391_ _1394_ core_0.execute.sreg_priv_control.o_d\[0\] _1395_ _1396_
+ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_0_19_207 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_376 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_176_359 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_87_696 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_129_242 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7651_ _1132_ _1102_ _3758_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_4863_ core_0.decode.i_imm_pass\[7\] _1341_ _1345_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_75_858 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_145_702 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_157_562 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_170_34 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_200_691 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6602_ _2929_ _2948_ _2949_ _2950_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_0_6_101 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_184_370 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_172_521 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_184_381 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7582_ core_0.execute.pc_high_out\[4\] _3695_ _3702_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_144_223 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4794_ core_0.fetch.prev_request_pc\[14\] net225 _0880_ net166 _1302_ vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_0_90_839 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_103_50 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_144_234 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_7_668 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6533_ _2907_ _0196_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_42_210 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_103_72 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_144_256 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_31_886 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_15_457 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6464_ _2121_ _2842_ _2096_ _2118_ _2294_ _2123_ _2843_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux4_4
XFILLER_0_113_632 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_125_492 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_95_1649 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_8203_ _0379_ clknet_leaf_2_i_clk core_0.execute.alu_mul_div.div_res\[12\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_179_76 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput110 net110 o_instr_long_addr[2] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
X_5415_ _1374_ _1856_ _1857_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6170__B1 _2022_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput121 net121 o_mem_addr[14] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
X_6395_ _1107_ _2769_ _2771_ _2775_ _2776_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XFILLER_0_88_85 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xoutput132 net132 o_mem_addr_high[0] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
Xoutput143 net143 o_mem_data[13] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_246_308 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput154 net154 o_mem_data[9] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
X_8134_ _0310_ clknet_leaf_105_i_clk core_0.execute.rf.reg_outputs\[2\]\[9\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xoutput165 net165 o_req_addr[13] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
X_5346_ core_0.execute.alu_mul_div.div_cur\[10\] _1789_ _1794_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xoutput176 net176 o_req_addr[9] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_56_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xoutput187 net187 sr_bus_addr[3] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_10_173 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_696 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_184_2721 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
Xoutput198 net198 sr_bus_data_o[13] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_227_533 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_195_53 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8065_ _0241_ clknet_leaf_111_i_clk core_0.execute.rf.reg_outputs\[6\]\[4\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5277_ _1433_ _1724_ _1725_ _0799_ _1726_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai211_4
XFILLER_0_215_706 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4079__A3 _0543_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5276__A2 core_0.execute.alu_mul_div.mul_res\[0\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
X_7016_ _3224_ _3230_ _3175_ _3232_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4228_ _0726_ _0845_ _0846_ _0847_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_199_418 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input28_I i_mem_data[1] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_3_545 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_4159_ core_0.dec_l_reg_sel\[1\] core_0.dec_l_reg_sel\[0\] _0778_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_97_405 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_106_Right_106 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__5028__A2 _1458_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6225__A1 _2608_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_223_772 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_39_975 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_179_142 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_39_986 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_78_630 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6776__A2 _3043_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4787__A1 core_0.fetch.prev_request_pc\[11\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7918_ _0009_ clknet_leaf_120_i_clk core_0.decode.oc_alu_mode\[6\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_4
XANTENNA__4787__B2 net163 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_167_348 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_93_611 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_144_90 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_527 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_104_1756 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5629__B _2018_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7849_ _0042_ clknet_leaf_64_i_clk core_0.fetch.out_buffer_data_instr\[26\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_195_2850 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6528__A2 _2190_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_65_346 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_19_763 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_53_508 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_817 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_135_212 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_80_305 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_81_839 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_93_699 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_230_37 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4003__A3 _0549_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5200__A2 _1444_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8195__CLK clknet_leaf_2_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xwire215 _0660_ net215 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_92_187 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_151_716 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_133_2108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_190_384 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_150_226 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_254 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_59_1224 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_58_i_clk_I clknet_4_14__leaf_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_265 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output96_I net96 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_799 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_103_142 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_131_462 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6700__A2 _2998_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5083__C _1531_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_115_1896 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_226_3227 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_218_533 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4695__S _1241_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5267__A2 _1715_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_206_717 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_218_588 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_245_374 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_205_216 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_144_2237 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_214_761 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4427__C _0963_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5019__A2 _0521_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_201_411 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_186_613 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6923__B _3139_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_241_591 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_213_282 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_198_473 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6767__A2 _3049_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4778__A1 _1290_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_201_444 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_69_674 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_84_611 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4242__A3 _0857_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_836 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_68_173 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_324 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_858 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_127_702 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_139_562 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_237_3356 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6519__A2 _2531_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7716__A1 _1196_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_126_223 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7192__A2 _3372_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_72_839 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_140_37 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_210 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput12 i_core_int_sreg[5] net12 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__4250__I0 net60 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput23 i_mem_data[11] net23 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_155_2377 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
Xinput34 i_mem_data[7] net34 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_25_766 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput45 i_req_data[16] net45 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_24_243 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_254 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xinput56 i_req_data[26] net56 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4950__B2 _1391_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput67 i_req_data[7] net67 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__4669__I _1224_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_208_Right_208 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_122_484 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5200_ _0700_ _1444_ _1446_ _1649_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_209_500 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6180_ core_0.execute.alu_mul_div.mul_res\[6\] _2567_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_0_237_842 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_199_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_58_77 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5131_ core_0.execute.rf.reg_outputs\[2\]\[9\] _1438_ _1580_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_236_330 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_236_341 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6455__A1 _2356_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5258__A2 _1696_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5062_ _1460_ net180 _1511_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or2_2
XFILLER_0_236_374 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_165_34 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_224_547 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_4013_ _0638_ _0594_ _0639_ _0640_ _0641_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai211_4
XANTENNA__8068__CLK clknet_leaf_107_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6207__A1 core_0.decode.oc_alu_mode\[11\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_0_504 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_211_208 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_189_440 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_0_515 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6833__B _3083_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6758__A2 _3049_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_189_484 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_176_101 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4769__A1 _1284_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_36_945 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_90_31 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5964_ _2271_ _2342_ _2354_ _2355_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_87_471 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_53 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7703_ _3773_ _3801_ _3802_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_4915_ _1378_ _1379_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_47_335 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_181_88 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5895_ core_0.decode.oc_alu_mode\[2\] _2287_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_4
XANTENNA__7707__A1 _1034_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_43_1025 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_74_132 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_192_649 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_157_370 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_7634_ _0743_ _3729_ _3746_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_35_508 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3992__A2 _0541_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_63_828 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4846_ _1280_ net44 _1170_ _1335_ _1336_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_0_191_148 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_75_699 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_16_711 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_7_454 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_62_327 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5194__A1 _1481_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7565_ _3673_ _3686_ _3687_ _1950_ _0448_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_4777_ core_0.fetch.prev_request_pc\[6\] _1285_ _0881_ net173 _1293_ vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_0_132_204 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_160_524 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6516_ core_0.execute.sreg_scratch.o_d\[15\] _2579_ _2534_ net7 _2894_ vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__4941__A1 _1301_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_210_3028 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_7496_ _3639_ _3641_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XTAP_TAPCELL_ROW_190_2791 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6447_ core_0.execute.sreg_scratch.o_d\[13\] _2579_ _2534_ net5 _2827_ vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_0_30_235 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_31_769 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_3_682 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_8_604 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6694__A1 _2990_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6378_ _2753_ _2759_ _2760_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_228_831 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_11_471 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8117_ _0293_ clknet_leaf_108_i_clk core_0.execute.rf.reg_outputs\[3\]\[8\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_227_330 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5329_ core_0.execute.alu_mul_div.div_cur\[5\] _1715_ _1763_ _1775_ _1776_ _1777_
+ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XTAP_TAPCELL_ROW_54_1165 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_227_352 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_227_363 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_8048_ _0224_ clknet_leaf_119_i_clk core_0.execute.rf.reg_outputs\[7\]\[3\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_output134_I net134 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_199_259 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_230_517 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_221_3168 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_242_399 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6749__A2 _3043_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_211_731 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_167_112 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5957__B1 _2257_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_210_241 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_168_657 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_39_836 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_39_858 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_109_702 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_182_104 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_167_189 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_65_1294 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_81_603 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_136_521 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_38_379 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3983__A2 _0578_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_182_148 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_636 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_93_496 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6921__A2 _3135_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_80_157 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_117_1914 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4932__A1 net194 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_574 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_151_557 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_232_3297 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7721__I1 core_0.decode.i_imm_pass\[5\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6685__A1 core_0.execute.rf.reg_outputs\[6\]\[8\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_131_292 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_219_820 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_232_Left_479 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_219_842 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_234_801 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6437__A1 _1061_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_206_514 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6437__B2 _1109_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_245_182 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4999__A1 _0769_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4999__B2 core_0.execute.rf.reg_outputs\[3\]\[0\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4463__A3 _1056_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_233_399 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6653__B _2984_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_158_123 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_159_646 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_202_764 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7928__CLK clknet_leaf_129_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_97_780 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_241_Left_488 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__4215__A3 _0830_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_186_454 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_33_904 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_9_708 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_482 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_202_797 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_201_296 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4700_ core_0.fetch.out_buffer_data_instr\[7\] net67 _1246_ _1248_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_45_828 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_56_154 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_60_45 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5680_ _2080_ _2070_ _2081_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_139_392 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7165__A2 _1227_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_72_625 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_127_543 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4631_ core_0.dec_jump_cond_code\[2\] _1189_ _1190_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6373__B1 _2534_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_13_672 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_71_135 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7915__D _0006_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_114_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6912__A2 _3129_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_114_226 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_154_395 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4923__A1 _1209_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7350_ _1458_ _1990_ _2886_ _1549_ _3519_ _3520_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai221_2
XFILLER_0_108_790 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5716__C _2092_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4562_ _1143_ _0005_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_4_457 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_52_371 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_130_708 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6301_ _2280_ core_0.execute.alu_mul_div.mul_res\[9\] _2685_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_142_579 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7281_ _3456_ _3459_ _1395_ _0392_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_69_65 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_92_1619 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_4493_ _1077_ _1079_ _1081_ _1085_ _1086_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_2
XANTENNA__5479__A2 _1585_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6232_ core_0.execute.sreg_scratch.o_d\[8\] _2579_ _2534_ net15 _2617_ vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_40_588 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_110_443 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_168_2524 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_110_454 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6163_ _2022_ _2548_ _2550_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_209_352 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5114_ _0789_ core_0.execute.rf.reg_outputs\[4\]\[11\] _0779_ _1563_ vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__5451__C _1822_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6094_ _2360_ _2482_ _2483_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_EDGE_ROW_191_Right_191 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__6979__A2 _3193_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_85_97 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_224_333 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5100__A1 _1543_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5045_ core_0.execute.rf.reg_outputs\[7\]\[12\] net232 _1443_ core_0.execute.rf.reg_outputs\[3\]\[12\]
+ _1494_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_109_82 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_224_355 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_196_207 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_79_224 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_196_229 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_19_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_79_257 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_419 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6996_ _1222_ _2436_ _3204_ _3213_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_1
XANTENNA__6600__A1 net22 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_220_583 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_165_616 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_179_2664 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_5947_ _2335_ _2336_ _2337_ _2338_ _2339_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_0_164_104 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_101_1726 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_164_115 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_192_2820 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3965__A2 _0594_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_839 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7156__A2 _1227_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5878_ core_0.dec_sreg_jal_over _2270_ _2271_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_146_863 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_705 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7617_ _3729_ _3733_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
Xclkbuf_4_7__f_i_clk clknet_3_3_0_i_clk clknet_4_7__leaf_i_clk vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__5167__B2 core_0.execute.rf.reg_outputs\[6\]\[7\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
X_4829_ _1280_ _1252_ _1323_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_133_524 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6903__A2 _3129_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_172_181 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7548_ _1955_ _3671_ _3672_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_0_16_574 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_133_557 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_133_568 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4390__A2 _0950_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7479_ _3626_ _3628_ _3629_ _1217_ _0420_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_160_387 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_31_566 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4102__I _0721_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_219_138 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_112_1855 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_101_487 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_216_823 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5890__A2 _1476_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_215_311 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7092__A1 core_0.execute.alu_mul_div.mul_res\[11\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_231_804 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_141_2207 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_230_303 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_231_837 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_67_1312 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6473__B _1457_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_205_2974 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_168_410 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4772__I _1283_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_780 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_168_454 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_195_262 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_39_644 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_211_594 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_155_104 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_38_132 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_123_1984 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_183_424 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_234_3315 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_38_154 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_94_772 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_109_521 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_149_690 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_183_435 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_234_3326 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7147__A2 _3209_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_93_271 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_171_608 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_422 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5158__A1 core_0.execute.rf.reg_outputs\[5\]\[6\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_53_124 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_658 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_170_107 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5158__B2 core_0.execute.rf.reg_outputs\[7\]\[6\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_30_37 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_109_598 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_124_524 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_152_833 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_41_308 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_136_395 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_10_631 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_152_2336 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_124_568 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_201_72 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_34_393 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_78_1452 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_1_416 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_111_218 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_438 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6658__B2 net26 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_10_728 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_120_741 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_292 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5330__A1 core_0.execute.alu_mul_div.div_cur\[5\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_219_650 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6367__C _1114_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_245_3455 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5881__A2 _2244_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5979__S _1558_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3892__A1 _0517_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_234_642 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7083__A1 _3177_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_34 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_222_804 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_234_664 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_55_56 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_163_2465 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_221_314 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6830__A1 _2967_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_221_325 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_89_1581 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_89_555 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4682__I _1236_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_89_566 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_159_410 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_49_408 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_18_731 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6850_ core_0.execute.rf.reg_outputs\[2\]\[15\] _3085_ _3098_ _3105_ vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_76_238 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5801_ _2200_ _0170_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__8106__CLK clknet_leaf_94_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5397__A1 core_0.execute.alu_mul_div.div_cur\[4\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_231_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XPHY_EDGE_ROW_8_Right_8 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
X_6781_ _2940_ _3064_ _3066_ _0285_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_3993_ _0517_ _0524_ _0527_ core_0.execute.rf.reg_outputs\[2\]\[9\] _0623_ vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_0_85_750 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_186_284 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_147_649 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5732_ _1765_ _2088_ _2133_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_4
XFILLER_0_174_457 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_18_839 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7138__A2 _1549_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_128_863 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5727__B _1689_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5149__A1 _1467_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5663_ _2058_ _2059_ _2064_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_127_384 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8256__CLK clknet_leaf_32_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_4_210 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6897__A1 net96 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7402_ net212 _3544_ _3545_ _3565_ _3566_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_4614_ core_0.dec_jump_cond_code\[2\] _1173_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_0_60_639 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5594_ _1702_ _1994_ _1995_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_111_50 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_4_243 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_170_663 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_842 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7333_ _2777_ _3497_ _3498_ _3505_ _3506_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or4_2
XFILLER_0_111_72 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4545_ _1127_ _1128_ _1129_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5018__I _1466_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_102_218 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_130_527 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6649__B2 net23 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7264_ _3443_ _3444_ _3445_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_40_374 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_111_741 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_96_41 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4476_ core_0.decode.i_instr_l\[3\] core_0.decode.i_instr_l\[2\] _1069_ vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_4
X_6215_ _2591_ _2593_ _2597_ _2600_ _2601_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai211_2
XPHY_EDGE_ROW_39_Right_39 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
X_7195_ _1024_ _1741_ _1736_ _3383_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_6146_ core_0.execute.sreg_priv_control.o_d\[6\] _1385_ _2254_ core_0.execute.sreg_scratch.o_d\[6\]
+ _2533_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_TAPCELL_ROW_51_1124 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3883__A1 _0518_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_29_90 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7074__A1 _1372_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6077_ _2013_ _2015_ _2465_ _2466_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_127_2040 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5085__B1 _1443_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6821__A1 _2946_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5028_ _1457_ _1458_ _1474_ _1476_ _1477_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA_input10_I i_core_int_sreg[3] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_206_39 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_240_667 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_67_216 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5388__A1 _1375_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_138_627 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6979_ core_0.execute.alu_mul_div.mul_res\[2\] _3193_ _3197_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_EDGE_ROW_48_Right_48 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_49_1097 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_177_273 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_48_441 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_177_295 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_137_137 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3938__A2 _0530_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_193_766 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_192_243 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_485 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4060__A1 _0567_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_62_1253 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_91_720 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_422 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_75_282 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_153_619 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_36_647 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_180_416 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_118_384 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_106_535 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_263 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_63_488 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_134_855 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5560__A1 _0972_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4363__A2 _0942_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_133_376 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_160_162 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_43_190 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_161_696 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7344__S _3502_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_31_352 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_EDGE_ROW_57_Right_57 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__5312__A1 _1515_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_8_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_73_1393 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7065__A1 _1224_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_216_653 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_204_815 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_243_461 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_204_826 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_99_842 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_188_527 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_240_3396 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_169_730 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_59_739 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_66_Right_66 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__7368__A2 _3510_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_230_177 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_86_547 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_168_251 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_169_785 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_128_104 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_196_593 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_772 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_73_208 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_184_744 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4051__A1 core_0.execute.rf.reg_outputs\[7\]\[4\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_156_457 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_183_243 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_625 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_658 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_137_682 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_143_129 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_42_617 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_26_168 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_842 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4354__A2 _0947_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_112_527 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_124_387 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_EDGE_ROW_75_Right_75 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
X_4330_ core_0.fetch.prev_request_pc\[3\] _0948_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_10_503 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_547 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4677__I _1232_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4261_ _0722_ _0879_ _0880_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_4
XANTENNA__6500__B1 _2594_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_120_593 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6000_ _2360_ _2390_ _2391_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5854__A2 net192 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_157_57 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_input2_I i_core_int_sreg[10] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_66_55 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4192_ _0810_ _0811_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_0_181_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5606__A2 _1476_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6803__A1 _2986_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_206_174 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7951_ _0129_ clknet_leaf_4_i_clk core_0.execute.alu_mul_div.div_cur\[7\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_206_185 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_206_196 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_84_Right_84 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_82_43 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_222_667 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7002__B _3175_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6902_ net98 _3135_ _3124_ _3136_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_221_155 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7882_ _0073_ clknet_leaf_85_i_clk core_0.decode.i_instr_l\[7\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_49_216 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__7359__A2 _3526_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_194_519 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_159_240 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6833_ core_0.execute.rf.reg_outputs\[2\]\[7\] _3092_ _3083_ _3096_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_65_709 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_147_413 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_176_2623 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_58_772 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6764_ core_0.execute.rf.reg_outputs\[4\]\[10\] _3049_ _3045_ _3056_ vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__4042__A1 core_0.execute.rf.reg_outputs\[7\]\[5\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_18_625 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3976_ _0565_ core_0.execute.rf.reg_outputs\[4\]\[10\] _0520_ _0607_ vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_0_174_243 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_422 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_18_647 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_45_433 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5715_ _2091_ _2092_ _2115_ _2116_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_134_107 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_18_669 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6695_ _1963_ _3016_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_190_758 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_21_759 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_116_855 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_31_80 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5646_ _2040_ _2047_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_72_274 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_86_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XPHY_EDGE_ROW_93_Right_93 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_131_836 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_130_313 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5577_ _1981_ _0177_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_13_352 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_131_858 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_198_86 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_672 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7819__B1 _3758_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7316_ _1400_ core_0.execute.sreg_irq_pc.o_d\[15\] _1428_ _1430_ _3490_ vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_4528_ _1034_ _1113_ _1115_ _0008_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_8296_ _0472_ clknet_leaf_87_i_clk core_0.dec_used_operands\[1\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_40_171 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input58_I i_req_data[28] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_130_379 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7295__A1 _3409_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6098__A2 _2486_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_193 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7247_ _1430_ _1408_ _2571_ _3390_ _3430_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_TAPCELL_ROW_187_2752 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_4459_ core_0.decode.oc_alu_mode\[1\] _1053_ _1054_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_217_417 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_229_288 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4648__A3 _1206_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_229_299 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7178_ _1231_ _3373_ core_0.execute.alu_mul_div.div_res\[8\] _3374_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_244_247 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7047__A1 _1224_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_13_Left_260 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
X_6129_ _1601_ _1624_ _2318_ _2517_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_99_116 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_99_138 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_213_634 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_197_313 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_240_431 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_29_859 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6270__A2 net208 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_202_2933 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_185_508 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_212_177 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_212_199 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_107_1798 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_218_3129 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6022__A2 _1683_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_198_2892 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_95_377 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_539 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_138_457 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_411 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_120_1954 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_36_433 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_166_799 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4584__A2 net157 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_107_822 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_119_693 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_136_2139 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_23_105 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_128_i_clk_I clknet_4_0__leaf_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_23_116 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7522__A2 _3640_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_180_279 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_138 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_161_460 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4698__S _1246_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_161_471 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_190 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_387 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_20_801 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_75_1411 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_32_683 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_121_368 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7286__A1 net74 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6089__A2 core_0.execute.alu_mul_div.mul_res\[4\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_229_3258 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_235_203 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5836__A2 _1444_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4639__A3 _1197_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_236_737 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_242_3414 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_147_2279 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5049__B1 _1486_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_160_2435 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_189_858 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_204_667 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_86_1540 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_99_683 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_182_Left_429 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_207_93 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_231_486 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_59_558 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7757__B _1284_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_156_221 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6013__A2 _2342_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7210__A1 _0810_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_86_399 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_157_766 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_39_271 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_39_282 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_422 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_55_753 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_116_107 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_156_287 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_15_606 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5500_ _1908_ _1929_ _1932_ _1933_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_42_403 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_617 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6480_ _1898_ _1117_ _2857_ _2858_ _2859_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_0_70_734 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_82_594 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7513__A2 _3646_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5431_ core_0.execute.alu_mul_div.div_cur\[8\] _1838_ _1816_ _1870_ _1871_ vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XTAP_TAPCELL_ROW_171_2564 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4327__A2 _0944_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_191_Left_438 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_2_511 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_469 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_180_791 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_113_858 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_97_1680 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_8150_ _0326_ clknet_leaf_106_i_clk core_0.execute.rf.reg_outputs\[1\]\[9\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_140_655 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_23_683 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5362_ core_0.execute.alu_mul_div.comp _0801_ _1810_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_0_22_171 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7277__A1 net73 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7101_ _1224_ _3262_ _3310_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_239_553 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4313_ core_0.fetch.prev_request_pc\[0\] _0851_ _0931_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_8081_ _0257_ clknet_leaf_114_i_clk core_0.execute.rf.reg_outputs\[5\]\[4\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_2
X_5293_ _1172_ _1739_ _1742_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_4
Xclkbuf_leaf_0_i_clk clknet_4_0__leaf_i_clk clknet_leaf_0_i_clk vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_7032_ _1226_ _1620_ _3246_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5827__A2 _2209_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_226_225 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4244_ _0834_ _0839_ _0848_ _0862_ _0863_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_0_242_718 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_226_269 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_242_729 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4175_ _0789_ _0793_ _0794_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_241_206 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_207_461 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_93_86 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_182_2693 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6252__A2 _1592_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_222_453 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_179_346 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7934_ _0112_ clknet_leaf_32_i_clk core_0.execute.sreg_priv_control.o_d\[6\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5031__I _1479_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_195_828 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_91 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_26_829 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_7865_ _0057_ clknet_leaf_59_i_clk core_0.fetch.prev_request_pc\[8\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_194_327 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_37_208 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_77_377 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7201__A1 _1414_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6816_ _3085_ _3086_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_203_18 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_92_314 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_46_1067 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4015__A1 _0567_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_65_539 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7796_ _3834_ _3860_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_148_777 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7752__A2 _1062_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_147_276 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6747_ core_0.execute.rf.reg_outputs\[4\]\[2\] _3043_ _3045_ _3047_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__5763__A1 _1756_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_175_596 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_3959_ _0584_ _0589_ _0591_ _0592_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_4
XFILLER_0_190_544 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_46_786 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_572 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6678_ _2961_ _2999_ _3007_ _0241_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_61_734 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7504__A2 _3640_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5629_ _1761_ _2019_ _2018_ _2030_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_103_335 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7268__A1 _1431_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_131_699 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output164_I net164 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_8279_ _0455_ clknet_leaf_27_i_clk core_0.execute.pc_high_buff_out\[0\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_2
XTAP_TAPCELL_ROW_57_1196 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_218_737 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5818__A2 _2215_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_228_37 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_245_556 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_70_1352 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_6_587 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7421__I _1283_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_109_1816 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_244_14 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_224_3199 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_213_431 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_54_i_clk_I clknet_4_11__leaf_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7440__A1 _3547_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6243__A2 _2034_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_213_464 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_201_604 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_69_823 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4254__A1 _0869_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_213_486 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_355 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_84_804 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_96_664 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_wire213_I _0689_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_138_210 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_200_158 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_96_686 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_113_18 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_139_766 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7743__A2 _1062_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_49 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_138_276 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_81_1481 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4557__A2 _1043_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_138_298 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_153_224 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_285 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_153_268 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_3_308 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5506__A1 _1367_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_51_244 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6554__I0 net119 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_12_609 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_121_121 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7259__A1 net85 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_110_839 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_20_664 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_121_198 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_236_512 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_138_37 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_208_236 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6656__B _2984_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6482__A2 _1386_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_217_792 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_223_239 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_37 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_78_119 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5980_ _1601_ _2370_ _2371_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_189_677 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_59_322 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_177_828 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_59_344 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4931_ _0722_ _0731_ _1395_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_0_63_89 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_87_664 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_144_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_7650_ _1279_ _1945_ _1031_ _0463_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_4862_ _0901_ _1306_ _1344_ _0088_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__5719__C _2092_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_86_174 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_86_185 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_731 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6601_ net29 _1149_ _2949_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_90_807 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_117_427 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7581_ _3673_ _3700_ _3701_ _1950_ _0450_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_7_636 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4793_ _1283_ _1301_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_6532_ net123 _2390_ _2906_ _2907_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_103_62 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_103_84 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_31_887 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_70_531 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_391 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_132_419 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_103_95 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_113_611 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7498__A1 _0720_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6463_ _2125_ _2128_ _2842_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_179_33 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_778 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_42_255 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_469 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_70_564 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_842 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_8202_ _0378_ clknet_leaf_1_i_clk core_0.execute.alu_mul_div.div_res\[11\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_179_55 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_2_330 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5414_ core_0.execute.alu_mul_div.div_cur\[7\] _1758_ _1780_ _1856_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__xor3_1
Xoutput100 net100 dbg_r0[6] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XANTENNA__6170__A1 core_0.decode.oc_alu_mode\[7\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput111 net111 o_instr_long_addr[3] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
X_6394_ _2300_ _1560_ _2642_ _2773_ _2774_ _2775_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai32_2
Xoutput122 net122 o_mem_addr[15] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA__6170__B2 core_0.decode.oc_alu_mode\[6\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput133 net133 o_mem_addr_high[1] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
X_8133_ _0309_ clknet_leaf_106_i_clk core_0.execute.rf.reg_outputs\[2\]\[8\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_88_97 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_101_839 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput144 net144 o_mem_data[14] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
X_5345_ core_0.execute.alu_mul_div.div_cur\[11\] _1752_ _1793_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__nor2_1
Xoutput155 net155 o_mem_long vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA__4720__A2 _1237_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput166 net166 o_req_addr[14] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
Xoutput177 net177 o_req_ppl_submit vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_239_372 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput188 net188 sr_bus_addr[4] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA_clkbuf_4_5__f_i_clk_I clknet_3_2_0_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_8064_ _0240_ clknet_leaf_94_i_clk core_0.execute.rf.reg_outputs\[6\]\[3\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_184_2722 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
Xoutput199 net199 sr_bus_data_o[14] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_10_185 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5276_ core_0.execute.alu_mul_div.i_mul core_0.execute.alu_mul_div.mul_res\[0\] _1725_
+ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_195_65 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_49_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_7015_ _3224_ _3230_ _3231_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__7834__CLK clknet_leaf_81_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4227_ _0726_ net61 _0846_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_214_217 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_3_546 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_4158_ _0768_ _0776_ _0777_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_69_108 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_97_417 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7422__A1 _3547_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_223_784 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_39_976 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_4089_ core_0.execute.rf.reg_outputs\[1\]\[0\] _0710_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_0_179_154 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_168_839 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_179_165 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_195_625 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7397__B _3516_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7917_ _0008_ clknet_4_3__leaf_i_clk core_0.execute.alu_mul_div.i_div vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5984__A1 _1689_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4814__B _1313_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_104_1757 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_7848_ _0041_ clknet_leaf_66_i_clk core_0.fetch.out_buffer_data_instr\[25\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_195_2851 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_194_168 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_148_574 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_230 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5736__A1 _1714_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_92_155 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_191_842 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_93_689 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7779_ core_0.dec_rf_ie\[3\] _3766_ _3833_ _3850_ _3851_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_80_317 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4105__I _0724_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_18_263 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_136_769 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_46_583 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_723 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_274 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_745 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_133_2109 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_34_767 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_33_244 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_6_691 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_59_1225 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_150_238 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_277 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_61_586 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6161__A1 _2010_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_103_154 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output89_I net89 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_116_i_clk clknet_4_4__leaf_i_clk clknet_leaf_116_i_clk vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_131_496 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4711__A2 _1237_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_115_1897 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_226_3228 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_108_18 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_233_537 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_144_2238 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_233_559 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_88_406 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4227__A1 _0726_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_214_795 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_213_261 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_159_839 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_213_294 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_201_434 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_83_1510 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_68_152 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_601 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_686 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4216__S _0723_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4242__A4 _0860_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_56_314 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_69_697 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_201_489 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_68_185 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_237_3357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_185_179 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7716__A2 _0514_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_83_133 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_84_656 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_204_72 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_72_807 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_84_667 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_154_522 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_182_842 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_83_166 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_127_769 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_83_188 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_181_352 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xinput13 i_core_int_sreg[6] net13 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_155_2367 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_25_745 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_617 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_531 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput24 i_mem_data[12] net24 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_155_2378 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
Xinput35 i_mem_data[8] net35 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__5555__B _1964_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput46 i_req_data[17] net46 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
Xinput57 i_req_data[27] net57 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__4950__A2 _1394_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput68 i_req_data[8] net68 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_40_715 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_428 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_597 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6152__A1 _1378_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_122_452 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_172_Right_172 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_150_794 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_34 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5130_ net103 _1492_ _1579_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_110_669 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_209_534 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5061_ _1466_ _0597_ _0602_ _0603_ _1510_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or4_4
Xclkbuf_leaf_80_i_clk clknet_4_13__leaf_i_clk clknet_leaf_80_i_clk vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__4466__A1 _1059_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_224_537 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4012_ _0532_ core_0.execute.rf.reg_outputs\[4\]\[7\] _0519_ _0640_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_0_205_751 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6207__A2 _2592_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_0_505 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_79_417 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7404__A1 _1980_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_0_516 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_220_710 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_205_784 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_95_i_clk clknet_4_7__leaf_i_clk clknet_leaf_95_i_clk vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_TAPCELL_ROW_36_946 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_149_327 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5963_ _2352_ _2353_ _2354_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_177_636 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_220_754 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_87_450 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7702_ _1085_ _1098_ _3762_ _3787_ _3801_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and4_1
X_4914_ core_0.dec_sreg_irt _1378_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_181_67 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_192_606 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_74_100 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5894_ core_0.decode.oc_alu_mode\[7\] _2286_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_3
XFILLER_0_59_185 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_74_111 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_114_50 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_191_105 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_47_347 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_43_1026 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_7633_ _3732_ _3744_ _3745_ _0458_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__5718__A1 _1124_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4845_ _0726_ _1261_ _1335_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_191_138 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3992__A3 _0543_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_7_422 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_173_842 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_28_572 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_317 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_177 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7564_ core_0.execute.pc_high_out\[1\] _3672_ _3687_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_90_648 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5194__A2 _1451_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4776_ _1290_ _1292_ _0054_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_117_279 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_7_488 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_99_63 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6515_ core_0.execute.alu_mul_div.div_cur\[15\] _1117_ _2890_ _2892_ _2893_ vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_4
X_7495_ _3639_ _3640_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_43_564 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_126_791 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_31_715 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_266 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_210_3029 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_190_2792 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_113_430 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_125_290 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_160_558 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_33_i_clk clknet_4_10__leaf_i_clk clknet_leaf_33_i_clk vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_130_82 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6446_ _2785_ _2759_ _2792_ _2826_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__6143__A1 _2202_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_70_383 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_rebuffer13_I net232 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_141_772 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_30_247 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_113_474 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_8_605 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6694__A2 _3000_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_101_636 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6377_ _1380_ _2757_ _2758_ _2759_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_2_193 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8116_ _0292_ clknet_leaf_108_i_clk core_0.execute.rf.reg_outputs\[3\]\[7\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_11_483 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5328_ core_0.execute.alu_mul_div.div_cur\[4\] _1695_ _1776_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA_input40_I i_req_data[11] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_54_1155 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_54_1166 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_48_i_clk clknet_4_12__leaf_i_clk clknet_leaf_48_i_clk vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__7643__A1 net206 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_8047_ _0223_ clknet_leaf_117_i_clk core_0.execute.rf.reg_outputs\[7\]\[2\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5259_ _1701_ _1702_ _1708_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__4457__A1 _1051_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_243_846 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_242_323 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_199_216 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_202_209 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_98_737 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_221_3169 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_211_743 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_195_422 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8162__CLK clknet_leaf_89_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5957__B2 core_0.execute.pc_high_out\[2\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_211_776 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_195_444 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_38_303 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_325 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_195_488 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_195_499 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_65_1295 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_38_369 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_65_166 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_626 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_164_853 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_109_769 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5185__A2 _1615_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_123_216 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_117_1915 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_80_169 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4932__A2 _1391_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_232_3298 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_61_372 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_22_737 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6134__A1 core_0.execute.alu_mul_div.i_mul vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6685__A2 _3006_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_238_629 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_131_282 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_5_Left_252 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_237_139 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_28_37 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_246_662 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7634__A1 _0743_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6437__A2 _1702_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_100_691 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_206_559 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_199_772 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_214_592 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_158_102 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_69 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5948__A1 net79 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5948__B2 _2245_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6070__B1 _2113_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_4_11__f_i_clk_I clknet_3_5_0_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_202_776 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_201_264 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4215__A4 _0833_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_33_905 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_29_314 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_241_Right_241 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_151_26 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_29_347 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_139_360 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_127_511 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_155_820 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_167_691 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_57_689 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_155_842 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_60_57 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_44_317 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7165__A3 _1230_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_44_328 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_115_706 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4630_ core_0.execute.alu_flag_reg.o_d\[1\] core_0.execute.alu_flag_reg.o_d\[0\]
+ _1181_ _1189_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_154_341 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_127_566 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_170_801 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_142_503 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6373__B2 net3 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_13_673 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_170_823 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_4_414 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4561_ _1137_ _1062_ _1064_ _1142_ _1143_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_107_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6300_ _2626_ _2672_ _2683_ _2684_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_4
X_7280_ _3409_ _3458_ _3459_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6125__A1 _1690_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_8_69 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6125__B2 _1631_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_100_30 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4492_ _1082_ _1084_ _1085_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_123_772 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_247 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_100_41 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6231_ _2542_ _2585_ _2616_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_40_567 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_110_411 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_88 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_168_2525 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_228_139 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6162_ _2022_ _2548_ _2549_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_176_34 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7625__A1 _3732_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5113_ core_0.execute.rf.reg_outputs\[2\]\[11\] _1438_ _1562_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_236_150 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6093_ _1117_ _2480_ _2481_ _2482_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_4
XFILLER_0_85_76 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5044_ core_0.execute.rf.reg_outputs\[2\]\[12\] _1438_ _1493_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5100__A2 _1548_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6844__B _3098_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_109_94 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_224_367 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_205_570 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_79_247 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_189_282 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_177_422 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6995_ core_0.execute.alu_mul_div.mul_res\[4\] _3212_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__6061__B1 _2264_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_48_634 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_94_239 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5946_ core_0.execute.pc_high_buff_out\[1\] _2249_ _2260_ net8 _2338_ vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_192_403 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_179_2665 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_75_431 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4611__A1 net155 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_118_500 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_47_144 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_36_807 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_48_667 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_101_1727 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_8_731 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5877_ core_0.dec_sreg_irt _1732_ _2269_ _2270_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XTAP_TAPCELL_ROW_192_2821 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_35_306 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7156__A3 _1364_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_75_486 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_118_544 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_145_341 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7616_ _3731_ _3732_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_62_114 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_145_352 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4828_ core_0.decode.i_instr_l\[11\] _1321_ _1322_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5167__A2 _1615_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6364__A1 _1107_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6364__B2 _1121_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_161_834 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_172_171 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7547_ _3637_ _3669_ _3670_ _3671_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4759_ core_0.decode.i_flush _1279_ _0813_ _1281_ _1282_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__nor4_2
XFILLER_0_172_193 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_160_344 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_597 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6116__A1 _1457_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_31_534 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7478_ net194 _1398_ _3628_ _3629_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_31_545 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4127__B1 _0745_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6667__A2 _3000_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_113_271 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6429_ _2808_ _2729_ _2102_ _2809_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_101_422 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_113_282 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4678__A1 _0804_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_112_1856 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_227_150 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_243_610 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_243_632 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_216_857 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7092__A2 _3300_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6754__B _3045_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_203_507 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_188_709 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_141_2208 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_67_1313 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4850__A1 core_0.decode.i_imm_pass\[1\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_205_2975 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_58_409 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_206 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_228 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_156_606 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_195_252 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_94_751 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_123_1985 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_155_116 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_453 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_234_3316 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_137_842 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_38_177 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_26_317 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_183_469 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_152_801 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5158__A2 _1604_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_26_339 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_136 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_124_514 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_170_119 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_163_160 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_191_480 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_10_632 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_81_478 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_489 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_152_2337 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8058__CLK clknet_leaf_99_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_78_1453 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_201_84 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_772 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_50_865 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6658__A2 core_0.ew_data\[14\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5866__B1 _2258_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_58 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_120_775 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5330__A2 _1715_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_245_3456 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7607__A1 core_0.execute.pc_high_out\[7\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_219_695 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3892__A2 _0524_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_146_37 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_206_345 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_55_46 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5094__A1 net94 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_206_367 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_89_512 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_163_2466 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_234_687 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6830__A2 _3086_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_79 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7479__C _1217_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_178_208 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_89_1582 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4841__A1 _0726_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_221_337 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_187_720 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_226_92 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_221_348 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_18_732 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_59_Left_306 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_77_718 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_159_422 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_159_433 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_202_551 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_34 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5800_ net132 _2199_ _2190_ _2200_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_6780_ core_0.execute.rf.reg_outputs\[3\]\[0\] _3065_ _3057_ _3066_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__6594__A1 net36 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3992_ _0565_ _0541_ _0543_ core_0.execute.rf.reg_outputs\[5\]\[9\] _0622_ vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_4
XANTENNA__5397__A2 _1812_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_174_403 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_71_67 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7791__B1 _3802_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_159_488 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_807 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5731_ _2130_ _2131_ _2113_ _2132_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_85_762 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_91_209 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_174_447 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_224_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_84_261 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_57_486 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_45_648 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6346__A1 _2113_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5662_ _2051_ _2054_ _2063_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__5149__A2 _1196_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_127_352 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__7543__B1 _1398_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_4_200 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_723 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_158 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_142_311 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4613_ _0811_ _1172_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_7401_ _3563_ net81 _3553_ _3564_ _3565_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_115_536 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6897__A2 _3130_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_182_491 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_4_222 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_72_489 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5593_ _1491_ _1994_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_4
XFILLER_0_154_193 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_174_2595 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_25_372 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_5_767 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7332_ _2646_ _2684_ _3504_ _3505_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
XPHY_EDGE_ROW_68_Left_315 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
X_4544_ _1049_ _1112_ _1128_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_40_331 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_4_288 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_556 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7263_ _1400_ core_0.execute.sreg_irq_pc.o_d\[8\] _1412_ _1430_ _3444_ vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__6649__A2 core_0.ew_data\[11\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_13_578 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4475_ _1067_ _1035_ _1068_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_0_96_31 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_187_66 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6214_ _1059_ _2018_ _2598_ _1620_ _2599_ _2600_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_0_96_64 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5462__C _1748_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_229_459 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_209_3020 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5321__A2 _1552_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7194_ net79 _1739_ _1740_ _3382_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_0_187_88 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6145_ core_0.execute.pc_high_out\[6\] _2257_ _2264_ core_0.execute.sreg_irq_pc.o_d\[6\]
+ _2532_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_TAPCELL_ROW_51_1125 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3883__A2 core_0.dec_r_reg_sel\[1\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_237_492 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_225_632 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7074__A2 _1224_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_31_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6076_ _1999_ _2009_ _2465_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or2_1
XTAP_TAPCELL_ROW_127_2041 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_224_142 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5969__I _2356_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_197_506 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6821__A2 _3086_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5027_ _1470_ _1471_ _1475_ _1476_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XPHY_EDGE_ROW_77_Left_324 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_197_528 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4832__A1 core_0.decode.i_instr_l\[12\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_178_731 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_221_860 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6034__B1 _2423_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_95_559 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6585__A1 core_0.ew_reg_ie\[7\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6978_ core_0.execute.alu_mul_div.mul_res\[2\] _3193_ _3196_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_49_1098 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_119_820 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_0_70 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_82_209 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5929_ _1819_ _1665_ _2320_ _2321_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_119_842 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_76_784 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_62_1254 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4060__A2 core_0.execute.rf.reg_outputs\[3\]\[3\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_134_801 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6337__A1 _2718_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_659 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_75_294 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_136 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_63_456 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_91_776 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_138_2170 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_173_480 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_180_439 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_output194_I net194 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_8_594 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6888__A2 _3106_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_86_Left_333 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_51_629 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_133_333 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4899__A1 _1231_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_161_664 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_16_394 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5560__A2 _1957_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_32_865 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6749__B _3045_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_133_388 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_160_174 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_114_591 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_102_753 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6468__C _2638_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_235_418 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_73_1383 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_73_1394 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_216_621 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_95_Left_342 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_215_142 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6273__B1 _2534_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_231_602 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_124_i_clk_I clknet_4_1__leaf_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_116_18 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_240_3397 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_169_742 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_86_515 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_98_375 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_129_606 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_211_370 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_168_263 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_784 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4051__A2 _0529_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_26_103 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4224__S _0824_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_82_732 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_352 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_147 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_143_119 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_137_694 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_183_299 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_23_790 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6879__A2 _3114_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_82_787 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_54_489 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_124_333 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5119__I _1567_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5000__A1 net88 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_151_130 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_35_692 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_41_139 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_2_715 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5551__A2 _1957_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_49_i_clk_I clknet_4_12__leaf_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6659__B _2984_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_151_174 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_239_702 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_2_737 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4958__I _1381_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4260_ _0875_ _0878_ _0879_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__5282__C _1195_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6500__A1 _1059_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5303__A2 _1713_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6500__B2 _2815_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_66_34 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5854__A3 _1199_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_226_429 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4191_ _0809_ _0810_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_157_69 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_219_492 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5789__I _2189_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_234_451 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_207_676 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_206_142 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_174_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6803__A2 _3065_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7950_ _0128_ clknet_leaf_4_i_clk core_0.execute.alu_mul_div.div_cur\[6\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_173_46 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6901_ _3128_ _3135_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
X_7881_ _0072_ clknet_leaf_52_i_clk core_0.decode.i_instr_l\[6\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_4
XFILLER_0_89_375 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_77_537 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6832_ _2972_ _3086_ _3095_ _0307_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_82_99 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_77_559 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8223__CLK clknet_leaf_8_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4417__I1 _0860_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_9_314 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_106_95 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_176_2624 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_64_209 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6763_ _2983_ _3042_ _3055_ _0278_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_3975_ core_0.execute.rf.reg_outputs\[7\]\[10\] _0530_ _0606_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_92_529 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_147_447 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4042__A2 _0529_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_73_710 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_570 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_412 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5714_ _1714_ _1501_ _2115_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6319__A1 _1109_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_128_661 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_17_136 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_73_754 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6694_ _2990_ _3000_ _3015_ _0249_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__4361__C _0963_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_122_50 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_128_683 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_456 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_72_242 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_17_158 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_73_776 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5645_ _2036_ _2038_ _2046_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_143_642 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_72_297 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_215_3090 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_142_152 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_103_517 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5576_ _1051_ _1172_ _1981_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__5542__A2 _1957_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_143_697 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_14_865 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_5_597 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_342 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_142_174 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_79_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_130_325 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5473__B _1841_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7315_ _2893_ _3393_ _3489_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_4527_ _1114_ _1053_ _1115_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__7819__A1 _1461_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_8295_ _0471_ clknet_leaf_88_i_clk core_0.dec_used_operands\[0\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_229_212 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7295__A2 _3471_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7246_ net84 _3398_ _3399_ _3428_ _3429_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_4458_ _1052_ _1053_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XTAP_TAPCELL_ROW_187_2753 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_245_716 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_229_278 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7177_ _1369_ _3372_ _3373_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
X_4389_ _0996_ _0966_ _0998_ _0999_ _0877_ net175 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XANTENNA__7047__A2 _1909_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6128_ _2300_ _2515_ _2516_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_0_99_106 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_213_602 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_198_804 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_198_815 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6059_ _2447_ _2448_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_198_826 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4805__A1 _1039_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_96_802 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_213_679 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_212_145 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_202_2934 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6007__B1 _2264_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6558__A1 net121 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_107_1799 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_178_594 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_198_2893 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_55_209 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_83_518 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4552__B _1132_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3947__I _0580_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_64_710 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_120_1955 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_153_417 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_165_277 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_834 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_165_299 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_91_562 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_275 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_798 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_118_193 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_51_426 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_134_664 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_17_692 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6730__A1 _2988_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_121_303 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5533__A2 _1957_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_50_i_clk_I clknet_4_12__leaf_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6479__B _1432_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4592__I0 core_0.ew_data\[2\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_75_1412 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_32_695 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_161 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_229_3259 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5297__A1 _1419_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_242_3415 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_216_451 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_36_37 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_189_804 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4219__S _0724_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_216_473 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6797__A1 _2977_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_207_50 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_160_2436 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_207_72 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_203_156 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_86_1541 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_203_167 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_99_695 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_188_369 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6549__A1 _2576_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_74_507 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_169_594 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7210__A2 _1734_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_250 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_55_710 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4024__A2 core_0.execute.rf.reg_outputs\[4\]\[6\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_129_469 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5277__C _0799_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_6_317 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_765 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_172_737 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_184_597 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_171_236 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_478 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_629 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5430_ _1233_ _1861_ _1869_ _1822_ _1870_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XTAP_TAPCELL_ROW_171_2565 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_140_612 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_124_174 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6572__I1 core_0.ew_reg_ie\[6\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_2_523 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4688__I _1236_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_97_1681 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_5361_ _1749_ _1808_ _1809_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_4
XFILLER_0_140_667 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_23_695 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4312_ _0905_ _0908_ _0911_ _0916_ _0930_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_7100_ _1230_ _1913_ _3308_ _3309_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__7277__A2 _3398_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_8080_ _0256_ clknet_leaf_118_i_clk core_0.execute.rf.reg_outputs\[5\]\[3\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5292_ _1739_ _1740_ _1741_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__5288__A1 _1414_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7031_ _1908_ _1631_ _3244_ _3245_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4243_ _0816_ _0819_ _0861_ _0862_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_0_120_391 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_10_389 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4174_ core_0.ew_reg_ie\[0\] core_0.ew_reg_ie\[1\] core_0.ew_reg_ie\[2\] core_0.ew_reg_ie\[3\]
+ _0769_ _0768_ _0793_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_184_34 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_93_43 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_124_2000 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_182_2694 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_117_61 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7933_ _0111_ clknet_leaf_25_i_clk core_0.execute.sreg_priv_control.o_d\[5\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_96_109 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_117_72 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_195_818 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_26_819 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5460__A1 _1822_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7864_ _0056_ clknet_leaf_60_i_clk core_0.fetch.prev_request_pc\[7\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_194_317 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_148_734 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_65_507 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_187_391 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6815_ core_0.ew_reg_ie\[2\] _2934_ _3085_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_2
XANTENNA__7201__A2 core_0.execute.sreg_irq_pc.o_d\[1\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_46_710 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_46_1068 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_9_133 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5212__A1 _0771_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7795_ _1049_ _1139_ _1092_ _1037_ _3781_ _3859_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XPHY_EDGE_ROW_186_Right_186 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_42_80 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6746_ _2946_ _3042_ _3046_ _0270_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__5763__A2 _1592_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3958_ _0590_ _0578_ _0591_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_163_737 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_163_748 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_702 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_562 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_162_247 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3889_ _0518_ _0525_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__inv_3
X_6677_ core_0.execute.rf.reg_outputs\[6\]\[4\] _3006_ _3004_ _3007_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_73_595 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_804 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_150_409 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_234 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_3_4_0_i_clk clknet_0_i_clk clknet_3_4_0_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_5628_ _2027_ _2028_ _2029_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_5_361 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6712__A1 _2956_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input70_I i_req_data_valid vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_103_314 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8119__CLK clknet_leaf_103_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_130_111 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_20_109 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_103_347 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5559_ core_0.execute.mem_stage_pc\[13\] _1955_ _1964_ _1975_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_41_470 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_130_177 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_8278_ _0454_ clknet_leaf_26_i_clk core_0.execute.pc_high_out\[7\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5931__B _1559_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_57_1197 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output157_I net157 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7229_ net81 _3400_ net82 _3414_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_217_248 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_70_1353 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_6_588 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_232_229 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_109_1817 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_198_634 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_198_667 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_186_807 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6762__B _3045_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_213_476 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4254__A2 _0870_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_312 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5451__A1 _1375_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_200_104 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_186_829 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_200_115 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_200_137 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_95_142 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_139_734 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_710 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5203__A1 net217 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_83_348 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_153_Right_153 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__6951__A1 _1088_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_126_428 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_138_288 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_154_737 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_166_597 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_64_551 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_81_1482 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_193_394 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_37_776 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_119_480 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_253 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_713 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_153_247 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_181_556 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_51_201 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_212 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_107_664 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_24_448 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_134_461 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_686 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6554__I1 _2825_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_110_807 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_122_667 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_632 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4317__I0 net67 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_208_204 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_236_524 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_209_738 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_102_391 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6429__S _2102_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_47_69 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_223_207 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_223_218 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_154_37 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_231_240 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7431__A2 _3543_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_189_667 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87_632 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_231_273 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_99_492 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_204_498 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4930_ _1393_ _1394_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_188_177 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_EDGE_ROW_32_Left_279 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_176_317 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_231_295 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5993__A2 _2383_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_209 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_75_827 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5288__B _1736_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_234_92 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4861_ core_0.decode.i_imm_pass\[6\] _1341_ _1344_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__7195__A1 _1024_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_185_862 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_129_244 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_157_553 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_200_671 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_137_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6600_ net22 _1148_ _2948_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_157_575 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_184_361 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4792_ _1290_ _1300_ _0062_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_28_754 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_120_Right_120 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
X_7580_ core_0.execute.pc_high_out\[3\] _3672_ _3701_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_43_702 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_55_562 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6531_ _2189_ _2906_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_27_264 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_404 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_27_286 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_31_888 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4412__S _0959_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7498__A2 _3640_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_43_768 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6462_ _2090_ _2547_ _2841_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_179_45 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_212_3060 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_70_576 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8201_ _0377_ clknet_leaf_2_i_clk core_0.execute.alu_mul_div.div_res\[10\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5413_ core_0.execute.alu_mul_div.div_cur\[7\] _1811_ _1855_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__nor2_1
Xoutput101 net101 dbg_r0[7] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_0_42_289 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_41_Left_288 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
X_6393_ _2062_ _2066_ _2071_ _2774_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_179_78 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput112 net112 o_instr_long_addr[4] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA__7723__S _1946_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_179_89 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput123 net123 o_mem_addr[1] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_23_492 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_632 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput134 net134 o_mem_addr_high[2] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
X_8132_ _0308_ clknet_leaf_111_i_clk core_0.execute.rf.reg_outputs\[2\]\[7\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5344_ _1790_ _1791_ _1792_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_140_475 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput145 net145 o_mem_data[15] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_10_120 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_100_317 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput156 net156 o_mem_req vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_100_339 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xoutput167 net167 o_req_addr[15] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_11_676 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_130_2070 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
Xoutput178 net178 sr_bus_addr[0] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
Xoutput189 net189 sr_bus_addr[5] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
X_8063_ _0239_ clknet_leaf_109_i_clk core_0.execute.rf.reg_outputs\[6\]\[2\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5275_ _1451_ _1456_ _1692_ _1723_ _1724_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XTAP_TAPCELL_ROW_184_2723 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_4226_ core_0.fetch.out_buffer_data_instr\[30\] _0845_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__inv_1
X_7014_ _3229_ _3230_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_199_409 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4157_ _0775_ _0776_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XTAP_TAPCELL_ROW_3_547 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_179_100 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_207_292 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_223_763 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_50_Left_297 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__7678__B _1078_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4088_ _0709_ net201 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__inv_4
XFILLER_0_168_807 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_39_977 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_222_273 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7916_ _0007_ clknet_leaf_121_i_clk core_0.decode.oc_alu_mode\[4\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_4
XFILLER_0_78_654 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5984__A2 _1665_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_194_125 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_77_142 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_210_457 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3995__A1 net103 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7847_ _0040_ clknet_leaf_66_i_clk core_0.fetch.out_buffer_data_instr\[24\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_104_1758 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_195_2852 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_92_123 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_220 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_191_832 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5736__A2 _1695_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_136_737 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_148_597 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7778_ _1315_ _3847_ _3850_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_18_242 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_439 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6729_ core_0.execute.rf.reg_outputs\[5\]\[11\] _3027_ _3031_ _3036_ vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xwire217 _1645_ net217 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_163_556 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4830__B _1170_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_212 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_163_578 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_116_461 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7489__A2 _1398_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6536__I1 _2482_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_59_1215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7733__I0 net180 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_59_1226 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_21_418 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_667 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_131_486 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_115_1887 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_115_1898 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_226_3229 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3960__I _0592_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7110__A1 _2778_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5153__S _1601_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_245_332 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5121__B1 net218 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5672__A1 _1702_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_205_229 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_144_2239 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_226_590 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_222_Right_222 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_214_741 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7413__A2 _3542_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_198_442 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_241_571 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4227__A2 net61 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5424__A1 core_0.execute.alu_mul_div.div_cur\[8\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_632 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_241_593 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_198_486 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_185_103 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_83_1511 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5975__A2 _2284_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_201_457 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7177__A1 _1369_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_139_553 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_237_3358 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_166_350 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_127_715 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_166_361 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6924__A1 _2994_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_84_679 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_71_318 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_126_247 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_182_865 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_64_370 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xinput14 i_core_int_sreg[7] net14 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_155_2368 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
Xinput25 i_mem_data[13] net25 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_141_206 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput36 i_mem_data[9] net36 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_80_863 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput47 i_req_data[18] net47 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_40_705 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput58 i_req_data[28] net58 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_3_139 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_12_407 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput69 i_req_data[9] net69 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_94_1640 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_150_773 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6667__B _2984_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_209_502 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_20_473 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3910__A1 _0539_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7101__A1 _1224_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_236_321 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5060_ _1460_ net179 _1509_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or2_2
XANTENNA__7652__A2 _1032_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_236_387 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_224_527 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4011_ core_0.execute.rf.reg_outputs\[7\]\[7\] _0529_ _0639_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4466__A2 _1053_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_74_34 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_165_58 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_165_69 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_205_763 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_0_506 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_0_517 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5415__A1 _1374_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_220_733 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_177_626 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5962_ _1195_ core_0.execute.sreg_irq_pc.o_d\[2\] _2353_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_36_947 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5966__A2 _2342_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_220_766 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_176_125 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7701_ core_0.dec_used_operands\[1\] _3766_ _3800_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_177_659 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_47_304 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4913_ _1375_ _1363_ _1376_ _1377_ _0106_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_0_87_473 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7168__A1 _1369_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_87_484 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_158_851 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5893_ _2004_ _2284_ _2285_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_176_158 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7632_ core_0.execute.pc_high_buff_out\[3\] _3731_ _1216_ _3745_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_43_1027 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5179__B1 _1437_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5718__A2 _2053_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_114_73 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_118_737 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4844_ core_0.decode.i_instr_l\[15\] _1307_ _1334_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6915__A1 net89 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_145_512 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_90_605 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_145_523 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_118_759 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_145_556 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7563_ net201 _3670_ _3685_ _3686_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_74_189 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_99_20 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4775_ core_0.fetch.prev_request_pc\[5\] _1285_ _0881_ net172 _1292_ vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_0_99_31 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_212 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6514_ _2891_ _0798_ _1432_ _2892_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_7494_ _1430_ _0810_ _2579_ _3639_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and3_2
XFILLER_0_132_228 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_99_86 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_130_61 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_190_2793 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_15_278 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_373 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6445_ _1798_ _2279_ _2823_ _2824_ _2825_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai22_4
XFILLER_0_141_751 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7340__A1 net201 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_790 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_clkbuf_leaf_97_i_clk_I clknet_4_7__leaf_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_8_606 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_113_486 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_228_800 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6376_ _1379_ core_0.execute.sreg_irq_pc.o_d\[11\] _2758_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_2_172 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_440 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_61_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_246_118 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_101_659 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_140_294 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8115_ _0291_ clknet_leaf_111_i_clk core_0.execute.rf.reg_outputs\[3\]\[6\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_2
XANTENNA__3901__A1 _0534_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5327_ _1766_ _1773_ _1774_ _1775_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_4
XTAP_TAPCELL_ROW_54_1156 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_239_192 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7951__CLK clknet_leaf_4_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_8046_ _0222_ clknet_leaf_117_i_clk core_0.execute.rf.reg_outputs\[7\]\[1\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5258_ _1695_ _1696_ _1703_ _1704_ _1706_ _1707_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai221_4
XANTENNA_input33_I i_mem_data[6] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4457__A2 _1032_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4209_ core_0.fetch.out_buffer_data_instr\[29\] _0828_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_243_858 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5189_ _1482_ _1637_ _1638_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_199_228 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_242_379 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_221_3159 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8307__CLK clknet_leaf_76_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4317__S _0725_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_195_412 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5957__A2 _2250_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_195_434 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3968__A1 _0533_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7159__A1 _1227_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_210_287 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6532__S _2906_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_182_117 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_19_540 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_65_1296 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_108_214 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6906__A1 net100 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_108_225 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_562 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_616 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_175_191 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_108_247 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_164_865 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_124_707 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5148__S _1596_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_74_690 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4393__A1 net85 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5375__C _1822_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_62_863 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_117_1916 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_116_280 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_151_559 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_232_3299 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_104_442 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_132_751 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6134__A2 core_0.execute.alu_mul_div.mul_res\[5\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_104_464 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_131_272 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7162__I core_0.execute.alu_mul_div.div_res\[3\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7634__A2 _3729_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_28_49 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_100_681 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_218_376 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_218_387 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_206_527 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_234_847 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_233_335 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_233_368 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_221_508 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_89_749 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7398__A1 _3543_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_44_37 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_199_784 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_159_626 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5948__A2 _2268_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_97_760 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_215_72 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_33_906 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_84_410 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_96_281 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_29_337 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_123 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_174_629 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_186_489 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_EDGE_ROW_106_Left_353 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_151_38 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_127_523 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_127_534 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_487 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_127_545 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_182_640 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_182_651 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_56_189 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_115 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6373__A2 _2579_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_13_663 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_65_690 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_115_718 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7570__A1 _3675_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_127_578 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_154_364 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_182_673 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_37_392 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_13_674 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_142_515 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4384__A1 _0991_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4560_ _1138_ _1141_ _1142_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_clkbuf_leaf_119_i_clk_I clknet_4_6__leaf_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4923__A3 _1386_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_502 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_37 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_181_194 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_142_559 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4491_ _1083_ _1084_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_40_535 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6125__A2 _2010_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_45 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7322__A1 _1209_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6230_ _2576_ _2614_ _2615_ _0185_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_122_283 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_228_107 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4687__A2 _1237_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_168_2526 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_115_Left_362 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
X_6161_ _2010_ _2463_ _2154_ _2548_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5112_ net90 _1492_ _1561_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_0_85_44 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6092_ core_0.execute.alu_mul_div.div_cur\[4\] _1432_ _2481_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_224_313 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5043_ _1446_ _1492_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_225_858 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_109_62 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_100_i_clk clknet_4_7__leaf_i_clk clknet_leaf_100_i_clk vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_192_34 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7389__A1 _3547_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_196_209 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_192_89 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6994_ _2436_ _3181_ _3211_ _0353_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_125_50 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_94_207 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_149_125 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6061__B2 core_0.execute.sreg_irq_pc.o_d\[4\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_124_Left_371 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_220_563 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_410 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_149_158 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5945_ core_0.execute.sreg_scratch.o_d\[1\] _2254_ _2250_ core_0.execute.sreg_irq_flags.o_d\[1\]
+ _2337_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_TAPCELL_ROW_179_2655 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_179_2666 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_115_i_clk clknet_4_4__leaf_i_clk clknet_leaf_115_i_clk vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_177_489 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_101_1728 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_118_512 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_192_2811 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_48_679 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5876_ _2245_ _2267_ _2268_ net72 core_0.dec_sreg_irt _2269_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XTAP_TAPCELL_ROW_192_2822 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_63_616 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_146_843 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7615_ _3729_ _3730_ _1953_ _3731_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XANTENNA__7156__A4 _3358_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_146_865 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4827_ _1305_ _1321_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA__7561__A1 core_0.execute.pc_high_buff_out\[1\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_62_126 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_435 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_718 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_118_589 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4375__A1 _0892_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_62_148 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7546_ _1209_ _2257_ _3670_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_44_863 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_133_537 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4758_ _0727_ _1168_ _1280_ _1281_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_70_170 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7477_ _3627_ _3628_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_4689_ core_0.fetch.out_buffer_data_instr\[2\] net60 _1241_ _1242_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_31_557 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_133_Left_380 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_141_570 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_31_568 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6428_ _2116_ _2124_ _1625_ _2808_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_3_492 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_219_118 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4678__A2 _1233_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5875__A1 core_0.dec_sreg_jal_over vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6359_ core_0.decode.oc_alu_mode\[3\] _1620_ _2741_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_2
XTAP_TAPCELL_ROW_112_1857 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_101_489 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6419__A3 _2695_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5627__A1 _2010_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_8029_ _0206_ clknet_leaf_51_i_clk net118 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_242_121 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_215_357 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_203_519 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_98_524 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_141_2209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_231_839 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_187_209 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_67_1314 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4850__A2 _1307_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_205_2976 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_168_401 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_230_349 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_196_732 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_168_423 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6052__A1 core_0.dec_mem_access vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_78_292 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_134 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_109_501 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_123_1986 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_234_3317 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_93_251 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_183_448 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_476 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_94_785 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_93_273 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_136_331 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_148_191 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_163_150 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4366__A1 _0965_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_163_172 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_120_i_clk_I clknet_4_3__leaf_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_136_397 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_191_492 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_10_633 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_152_2338 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7304__A1 _2859_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_384 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_78_1443 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_105_762 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_78_1454 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_50_855 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_120_710 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_94_i_clk clknet_4_7__leaf_i_clk clknet_leaf_94_i_clk vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_22_579 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_91_1610 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5866__A1 core_0.execute.pc_high_out\[0\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_120_765 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5866__B2 net106 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_120_798 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_245_3457 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_219_674 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_218_173 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_207_836 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3892__A3 _0527_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6291__A1 _1121_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5094__A2 _1492_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_163_2467 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_233_187 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_199_570 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_89_1583 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_45_i_clk_I clknet_4_9__leaf_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_32_i_clk clknet_4_10__leaf_i_clk clknet_leaf_32_i_clk vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_TAPCELL_ROW_18_733 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_230_861 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_186_220 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_162_37 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3991_ _0517_ core_0.execute.rf.reg_outputs\[3\]\[9\] net231 _0621_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_2
XANTENNA__7791__A1 core_0.decode.i_instr_l\[14\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_85_741 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_147_629 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_29_134 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7791__B2 core_0.decode.i_instr_l\[11\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_174_415 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_186_286 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5730_ _1689_ _2123_ _2131_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_45_616 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_104 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_128_865 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5661_ _2045_ _2050_ _2061_ _2062_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_4
Xclkbuf_leaf_47_i_clk clknet_4_12__leaf_i_clk clknet_leaf_47_i_clk vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_5_702 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_217_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_115_504 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__7543__B2 core_0.execute.sreg_irq_flags.o_d\[4\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_72_457 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_7400_ _3547_ _1961_ _3564_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_60_608 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8002__CLK clknet_leaf_48_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4612_ _1171_ net122 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_26_863 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_212 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_182_481 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5592_ _1713_ net214 _1993_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_0_111_30 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_174_2596 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_170_643 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7331_ _3499_ _3500_ _3501_ _3503_ _3504_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor4_2
XFILLER_0_40_310 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_384 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_13_524 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_53_693 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4543_ _1037_ _1092_ _1127_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_25_395 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_130_518 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5516__S _1946_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_111_96 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4109__A1 net19 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7262_ _2652_ _3391_ _3443_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4474_ core_0.decode.i_instr_l\[5\] _1067_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__inv_1
XANTENNA__5857__A1 net186 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6213_ _2286_ _1758_ _2155_ _1686_ _2599_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_0_40_387 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7016__B _3175_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_110_242 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7193_ _2891_ _3381_ _3357_ _0382_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_209_3021 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7731__S _1946_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6144_ _2268_ _2531_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_110_297 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5609__A1 _1693_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_51_1126 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6855__B _3098_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6347__S _1625_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6075_ core_0.decode.oc_alu_mode\[4\] _2461_ _2463_ _2464_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__nand3_1
XTAP_TAPCELL_ROW_127_2031 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6282__A1 _2133_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_127_2042 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_213_817 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5026_ core_0.dec_alu_carry_en core_0.execute.alu_flag_reg.o_d\[1\] _1475_ vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_24_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_169_209 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_240_636 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4832__A2 _1321_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_212_349 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_45_80 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6034__A1 _1121_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_177_220 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7231__B1 _3399_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6034__B2 _1107_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_138_607 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_193_702 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6977_ _3175_ _2322_ _3181_ _2386_ _3195_ _0352_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_0_177_253 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_88_590 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6585__A2 _2934_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7782__A1 _1136_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_49_1099 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_178_798 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_76_752 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_177_286 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5928_ _1819_ _1637_ _2320_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5793__B1 _1615_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_627 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_62_1255 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_61_90 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_118_342 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5859_ _2251_ _1197_ _2252_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__7534__A1 _3581_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_8_562 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_91_766 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_138_2171 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_91_788 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_537 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_161_632 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_173_492 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_44_671 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4899__A2 _1362_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_90_287 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7529_ core_0.execute.sreg_scratch.o_d\[14\] _3646_ _3651_ _3660_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_90_298 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output187_I net187 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_32_855 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_31_343 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_102_732 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_101_220 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_102_776 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_102_798 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_73_1384 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_216_633 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_204_817 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5076__A2 _1522_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6273__B2 net16 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_230_102 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_240_3387 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_98_354 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_240_3398 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_169_754 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_86_527 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_98_387 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5895__I core_0.decode.oc_alu_mode\[2\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7773__A1 _1136_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_129_629 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_183_212 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_39_487 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_627 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_26_115 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_94_593 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_183_267 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_744 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_171_418 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4339__A1 core_0.fetch.prev_request_pc\[14\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_54_457 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_124_301 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_136_161 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_192_790 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_23_791 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_152_632 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5000__A2 _1446_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_229_Left_476 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_151_142 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_22_321 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_112_518 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_152_687 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_105_570 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_50_663 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_685 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5839__A1 _0177_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_387 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_10_527 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_239_769 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4190_ _0754_ _0756_ _0797_ _0808_ _0809_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and4_1
XANTENNA__5854__A4 _1200_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_207_611 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_238_Left_485 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_173_14 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4275__B1 _0844_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4814__A2 core_0.fetch.submitable vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_167_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_EDGE_ROW_167_Right_167 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_82_34 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6900_ _2956_ _3129_ _3134_ _0336_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_7880_ _0071_ clknet_leaf_47_i_clk core_0.decode.i_instr_l\[5\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_4
XFILLER_0_106_30 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_89_387 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6831_ core_0.execute.rf.reg_outputs\[2\]\[6\] _3092_ _3083_ _3095_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_89_398 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_159_242 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_187_562 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_175_702 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_202_371 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7764__A1 _1048_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_159_275 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4578__A1 core_0.ew_data\[3\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_9_326 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6762_ core_0.execute.rf.reg_outputs\[4\]\[9\] _3049_ _3045_ _3055_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_147_437 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_176_2625 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_3974_ core_0.execute.rf.reg_outputs\[1\]\[10\] _0605_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_119_139 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_45_402 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5713_ _2103_ _2110_ _2113_ _2114_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_116_802 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7516__A1 net216 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6693_ core_0.execute.rf.reg_outputs\[6\]\[12\] _3006_ _3004_ _3015_ vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_122_62 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_143_621 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_5_521 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5644_ _2026_ _2034_ _2044_ _2045_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_0_155_481 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_26_660 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_143_632 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_155_492 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_215_3091 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_13_310 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_170_451 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5575_ _1980_ _0742_ _0165_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_14_855 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_5_587 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_143_687 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7314_ _1977_ _3483_ _3488_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__4750__A1 net59 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_13_354 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4526_ _0798_ _1114_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XANTENNA__7819__A2 _1134_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_198_88 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8294_ _0470_ clknet_leaf_45_i_clk core_0.dec_sreg_load vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_229_202 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7245_ _3426_ _3427_ _3428_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_111_551 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_111_562 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4457_ _1051_ _1032_ _1052_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_187_2754 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_217_419 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7176_ _1223_ _1809_ _1810_ _3372_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_4
X_4388_ _0843_ _0947_ _0970_ _0999_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_6127_ _2304_ _2515_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__7047__A3 core_0.execute.alu_mul_div.cbit\[1\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6255__A1 _1061_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6255__B2 _1109_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6058_ net186 _1201_ _2262_ _2447_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_4
XFILLER_0_212_102 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_3_0_0_i_clk clknet_0_i_clk clknet_3_0_0_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XANTENNA__4805__A2 _1307_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5009_ core_0.decode.oc_alu_mode\[11\] _1458_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__inv_4
XPHY_EDGE_ROW_134_Right_134 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__8048__CLK clknet_leaf_119_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6007__A1 net10 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_202_2935 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6007__B2 core_0.execute.sreg_irq_pc.o_d\[3\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_240_488 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_95_324 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_95_335 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_178_562 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6558__A2 _1985_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output102_I net102 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_198_2883 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_165_212 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_198_2894 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_119_640 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_138_459 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_120_1956 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_153_407 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_125_109 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_63_232 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_106_301 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6540__S _2906_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4124__I _0743_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_457 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_174_790 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_619 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_134_632 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_20_750 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_106_356 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_133_142 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_16_181 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6730__A2 _3022_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_161_473 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_161_484 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_663 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_75_1413 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4592__I1 core_0.ew_data\[10\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_242_3416 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6246__A1 _1121_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5049__A2 _1435_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_216_485 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6797__A2 _3064_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_243_282 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_189_838 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_204_647 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_99_652 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_160_2437 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_207_62 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_101_Right_101 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_188_337 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_86_1542 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_188_359 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6942__C _1223_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_86_302 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_28_850 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_87_836 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_59_538 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87_858 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_157_702 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_169_562 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6549__A2 _2716_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_200_831 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_52_37 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_52_48 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_86_368 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_129_437 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_184_532 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_582 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_744 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_144_418 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_171_204 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_109_150 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4034__I net215 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_109_161 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_70_703 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_125_621 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_125_632 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_137_492 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4980__A1 _1419_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_14_107 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_42_438 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_124_142 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_152_451 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_140_602 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7345__I _0722_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_171_2566 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6721__A2 _3027_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_113_838 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_124_164 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_152_473 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_140_624 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_97_1671 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_239_500 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_535 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_97_1682 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_5360_ _1750_ _1807_ _1808_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_140_646 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_11_836 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4311_ _0884_ _0900_ _0922_ _0928_ _0929_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai22_2
XPHY_EDGE_ROW_236_Right_236 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_77_34 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_168_47 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_195 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_858 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5291_ net72 _0810_ _1740_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_168_58 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_120_370 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6485__A1 _1380_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7030_ _1908_ _1637_ _3244_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4242_ _0851_ _0854_ _0857_ _0860_ _0861_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_0_10_379 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_77_89 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_226_238 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4173_ core_0.ew_reg_ie\[4\] core_0.ew_reg_ie\[5\] core_0.ew_reg_ie\[6\] core_0.ew_reg_ie\[7\]
+ _0769_ _0768_ _0792_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux4_4
XFILLER_0_207_441 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6237__A1 _1379_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_235_772 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_124_2001 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_234_271 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_207_485 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_182_2695 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_78_803 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7932_ _0110_ clknet_leaf_24_i_clk core_0.execute.sreg_priv_control.o_d\[4\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_179_337 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7863_ _0055_ clknet_leaf_59_i_clk core_0.fetch.prev_request_pc\[6\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_222_499 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_89_195 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_203_691 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_187_381 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6814_ _2996_ _3065_ _3084_ _0300_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_147_212 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5468__C _1748_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7794_ _0539_ _1134_ _3858_ _1279_ _0506_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__7908__CLK clknet_leaf_83_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_93_839 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_175_543 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_46_1069 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4015__A3 _0548_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_217_3120 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_133_72 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_148_779 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6745_ core_0.execute.rf.reg_outputs\[4\]\[1\] _3043_ _3045_ _3046_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_58_593 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3957_ net91 _0590_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_135_418 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_190_524 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_18_457 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4971__A1 _1419_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_46_788 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_45_265 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6676_ _2998_ _3006_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_46_799 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_33_416 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3888_ _0523_ _0524_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_33_427 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_135_2130 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_6_863 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5627_ _2010_ _2011_ _2013_ _2014_ _2028_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_115_142 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6712__A2 _3021_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_116_698 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_663 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5558_ _0977_ _1956_ _1974_ _0154_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA_input63_I i_req_data[3] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_13_173 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4509_ _1037_ _1074_ _1099_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_8277_ _0453_ clknet_leaf_26_i_clk core_0.execute.pc_high_out\[6\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_2
XPHY_EDGE_ROW_203_Right_203 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
X_5489_ _1367_ _1914_ _1918_ _1921_ _1922_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai22_2
XANTENNA__5279__A2 _0798_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7228_ net82 net81 _3400_ _3413_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and3_1
XTAP_TAPCELL_ROW_57_1198 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_217_216 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_7159_ _1227_ _1364_ _3361_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_70_1354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6228__A1 _2242_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_232_208 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_6_589 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_109_1818 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_225_271 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_146_2270 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_198_613 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_244_16 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_225_282 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_201_617 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_240_263 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_201_628 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_95_110 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_139_702 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_69_858 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_84_839 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5203__A2 _1650_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6400__A1 core_0.execute.alu_mul_div.div_res\[12\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_166_565 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_49_593 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_138_267 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_193_384 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6951__A2 core_0.execute.alu_mul_div.comp vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_81_1483 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_153_226 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_154_749 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4962__A1 _1381_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_153_259 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_427 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_91_382 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_676 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_698 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_134_484 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_279 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6467__A1 _1713_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_208_238 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_217_761 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_217_772 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6953__B _3173_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_232_731 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_189_646 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_232_786 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_59_324 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_176_307 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_87_666 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_185_830 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_59_368 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_129_212 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4860_ _0907_ _1306_ _1343_ _0087_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_75_839 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_129_234 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_170_37 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_184_351 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4791_ core_0.fetch.prev_request_pc\[13\] net225 _0880_ net165 _1300_ vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_0_184_373 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_99_1700 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_117_429 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_144_215 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6530_ _2576_ _2334_ _2905_ _0195_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__4953__B2 _1391_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_574 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_82_360 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_27_276 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_416 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_55_585 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_172_568 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_43_736 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_125_440 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_31_889 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6461_ _1121_ _2085_ _2840_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_103_97 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8200_ _0376_ clknet_leaf_7_i_clk core_0.execute.alu_mul_div.div_res\[9\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_2_310 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5412_ _1853_ _1854_ _0128_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_212_3061 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_2_321 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6392_ core_0.decode.oc_alu_mode\[11\] _2772_ _2773_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xoutput102 net102 dbg_r0[8] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_51_780 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xoutput113 net113 o_instr_long_addr[5] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_101_819 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_112_145 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_140_454 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput124 net124 o_mem_addr[2] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
X_8131_ _0307_ clknet_leaf_112_i_clk core_0.execute.rf.reg_outputs\[2\]\[6\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_2
X_5343_ core_0.execute.alu_mul_div.div_cur\[11\] _1752_ _1791_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__xor2_1
Xoutput135 net135 o_mem_addr_high[3] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
Xoutput146 net146 o_mem_data[1] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_2_387 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xoutput157 net157 o_mem_sel[0] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_239_352 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6458__A1 core_0.ew_data\[13\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput168 net168 o_req_addr[1] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XTAP_TAPCELL_ROW_130_2071 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
Xoutput179 net179 sr_bus_addr[10] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_239_374 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_227_514 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8062_ _0238_ clknet_leaf_109_i_clk core_0.execute.rf.reg_outputs\[6\]\[1\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_11_688 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5274_ _1699_ _1722_ _1723_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_2
XTAP_TAPCELL_ROW_184_2724 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_7013_ core_0.execute.alu_mul_div.mul_res\[5\] _3228_ _3229_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_4225_ net55 core_0.fetch.out_buffer_data_instr\[25\] _0824_ _0844_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_4
XFILLER_0_10_198 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5130__A1 net103 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4367__C _0963_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_128_72 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_4156_ core_0.dec_l_reg_sel\[0\] _0775_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__inv_2
XFILLER_0_223_731 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_207_282 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_3_548 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_4087_ net95 _0521_ _0703_ _0708_ _0709_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai22_4
XTAP_TAPCELL_ROW_223_3190 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_39_978 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6630__A1 _2936_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_93_i_clk_I clknet_4_6__leaf_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7915_ _0006_ clknet_leaf_119_i_clk core_0.decode.oc_alu_mode\[3\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_2
XANTENNA__4383__B _0970_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_195_627 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_194_104 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_194_115 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_148_521 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7846_ _0039_ clknet_leaf_67_i_clk core_0.fetch.out_buffer_data_instr\[23\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_194_137 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3995__A2 _0578_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_53_80 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_66_839 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_104_1759 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7186__A2 _3372_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_176_863 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_195_2853 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_92_135 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_136_727 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7777_ _1136_ _3849_ _0498_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_4989_ _1437_ _1438_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_19_755 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5736__A3 _1696_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_190_310 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_175_384 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6728_ _2986_ _3022_ _3035_ _0263_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_18_265 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_61_500 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4944__B2 _1391_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_151_708 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_18_287 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6146__B1 _2254_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_61_544 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6659_ core_0.execute.rf.reg_outputs\[7\]\[14\] _2935_ _2984_ _2995_ vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__7489__A3 _1206_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_59_1216 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_61_566 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8236__CLK clknet_leaf_36_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6697__A1 _2992_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_103_112 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_5_192 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_103_156 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8329_ _0505_ clknet_leaf_91_i_clk core_0.dec_r_reg_sel\[1\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__dffq_4
XFILLER_0_41_290 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_103_189 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_246_812 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_115_1888 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6449__A1 _2447_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_226_3219 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7110__A2 _3181_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_100_863 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5672__A2 _1491_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6773__B _3057_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_198_410 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6621__A1 _2929_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_198_454 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5424__A2 _1812_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_201_403 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5389__B _1816_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_213_274 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_69_644 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_83_1512 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_68_132 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_96_452 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_154 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_201_469 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_699 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7177__A2 _3372_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_237_3359 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_182_811 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6924__A2 _3130_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_154_524 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_83_168 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_52_511 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_596 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_382 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_142_719 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xinput15 i_core_int_sreg[8] net15 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_25_747 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_4_619 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_155_2369 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
Xinput26 i_mem_data[14] net26 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xinput37 i_mem_exception net37 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
Xinput48 i_req_data[19] net48 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xinput59 i_req_data[29] net59 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__6688__A1 _2983_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_122_432 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_150_741 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_110_605 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_94_1641 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_20_441 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_236_311 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_58_69 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5112__A1 net90 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_209_558 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_179_Left_426 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
X_4010_ core_0.execute.rf.reg_outputs\[1\]\[7\] _0638_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XANTENNA__6860__A1 _2951_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6683__B _3004_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_115_i_clk_I clknet_4_4__leaf_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4982__I _1430_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_0_507 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_0_518 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6612__A1 net24 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_189_476 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5961_ net80 _2268_ _2351_ _2245_ core_0.dec_sreg_irt _2352_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_0_232_594 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_220_745 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_176_115 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_36_948 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_87_452 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7700_ _0766_ _1134_ _3789_ _3799_ _1279_ _0471_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_4912_ _1223_ _1221_ _1377_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_181_47 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_59_165 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3977__A2 _0594_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_90_45 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_176_137 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_48_839 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5892_ _1687_ _1473_ _1470_ _2284_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_181_69 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_47_316 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7168__A2 _1915_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_158_863 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87_496 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7631_ net203 _3733_ _3743_ _3744_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_114_52 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_188_Left_435 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_47_349 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4843_ _1331_ _1333_ _0080_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_157_362 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_43_1028 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_118_727 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6915__A2 _3135_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_185_693 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_23_72 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_184_170 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8259__CLK clknet_leaf_36_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_145_535 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7562_ _3682_ _3683_ _3684_ _3670_ _3685_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__4926__A1 _1381_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4774_ _1290_ _1291_ _0053_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_117_259 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_7_468 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_145_579 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6513_ core_0.execute.alu_mul_div.div_res\[15\] _2891_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__inv_2
XFILLER_0_71_842 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_55_393 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_160_516 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_160_527 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7493_ _3637_ _1208_ _1395_ _3638_ _0425_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_31_706 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_132_2100 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6679__A1 core_0.execute.rf.reg_outputs\[6\]\[5\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_190_2794 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6444_ core_0.execute.alu_mul_div.div_res\[13\] _2332_ _0800_ _2824_ vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA__7340__A2 _3502_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_141_763 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6375_ net74 _2531_ _2756_ _2537_ _2757_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XTAP_TAPCELL_ROW_8_607 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_3_696 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_100_104 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8114_ _0290_ clknet_leaf_107_i_clk core_0.execute.rf.reg_outputs\[3\]\[5\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_228_823 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5326_ core_0.execute.alu_mul_div.div_cur\[3\] _1765_ _1774_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_EDGE_ROW_197_Left_444 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__3901__A2 _0535_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_54_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_54_1157 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_8045_ _0221_ clknet_leaf_93_i_clk core_0.execute.rf.reg_outputs\[7\]\[0\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5257_ _1705_ _1693_ _1525_ _1530_ _1706_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor4_4
XANTENNA__6851__A1 _2996_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_243_837 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_242_314 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4208_ _0723_ net62 _0826_ _0827_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_4
X_5188_ _1632_ _1636_ _1637_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_2
XANTENNA_input26_I i_mem_data[14] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4139_ _0535_ _0536_ _0758_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__6603__A1 _2930_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7201__C _1736_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_223_594 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_167_104 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_167_126 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3968__A2 _0541_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_210_255 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_195_468 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7159__A2 _1364_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4090__A1 _0565_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_327 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_176_660 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5937__B _0799_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_164_811 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7829_ _0022_ clknet_leaf_58_i_clk core_0.fetch.out_buffer_data_instr\[6\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_109_727 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_65_1297 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6906__A2 _3135_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_552 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_749 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_93_488 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_163_343 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_34_522 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_124_719 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4393__A2 _0883_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_61_330 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5590__A1 _1713_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_117_782 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_117_1917 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_163_398 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_61_352 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_151_549 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_output94_I net94 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_104_454 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_131_240 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5342__A1 core_0.execute.alu_mul_div.div_cur\[10\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5893__A2 _2284_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_load_slew216_I _0648_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_246_642 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6059__I _2447_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_234_815 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_4_12__f_i_clk clknet_3_6_0_i_clk clknet_4_12__leaf_i_clk vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_245_196 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_201_Left_448 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_233_347 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_89_717 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_88_205 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_214_594 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_198_262 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_202_745 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_158_104 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_201_233 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6070__A2 _1601_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_202_778 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_186_457 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_33_907 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_57_636 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6950__C _1223_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_60_26 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_60_37 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_606 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4908__A1 _1372_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_210_Left_457 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_154_354 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_13_664 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_71_127 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_231_72 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_53_842 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4384__A2 _0966_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_142_527 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA_clkbuf_leaf_41_i_clk_I clknet_4_11__leaf_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4490_ core_0.decode.i_instr_l\[6\] core_0.decode.i_instr_l\[4\] core_0.decode.i_instr_l\[5\]
+ _1083_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_4
XANTENNA__7322__A2 _2265_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_100_32 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5333__A1 core_0.execute.alu_mul_div.div_cur\[7\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4136__A2 core_0.decode.o_submit vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_110_413 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_100_65 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_21_772 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_100_76 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6160_ _2294_ _2545_ _2546_ _2547_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XTAP_TAPCELL_ROW_168_2527 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_20_260 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_110_457 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_110_468 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_197_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5111_ _1532_ _1555_ _1559_ _1560_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_6091_ core_0.execute.alu_mul_div.div_res\[4\] _2332_ _2479_ _2480_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_85_56 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_176_69 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_236_152 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5097__B1 _1443_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6833__A1 core_0.execute.rf.reg_outputs\[2\]\[7\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
X_5042_ _0576_ _1483_ _1485_ _1490_ _1491_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_0_85_78 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_236_196 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_79_205 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_79_227 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6993_ _3208_ _3210_ _3189_ _3211_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_220_531 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7729__S _1946_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6061__A2 _2254_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_149_137 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5944_ core_0.execute.sreg_data_page _1385_ _2257_ core_0.execute.pc_high_out\[1\]
+ _2336_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_TAPCELL_ROW_179_2656 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_75_422 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87_282 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_192_416 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_146_811 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_101_1729 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_5875_ core_0.dec_sreg_jal_over _1202_ _2268_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or2_2
XFILLER_0_118_524 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_192_2812 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_75_477 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_145_321 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7614_ core_0.dec_sreg_jal_over _0732_ _3730_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_63_628 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4826_ _1320_ _0076_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_90_414 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7561__A2 _3682_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_28_382 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_522 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_138 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_141_72 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_161_814 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_172_151 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7545_ net77 _1742_ _1206_ _3669_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_105_207 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5572__A1 _1980_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_7_276 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4757_ _0726_ _1280_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_43_341 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_298 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_133_549 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_161_858 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_114_741 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_374 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7476_ net210 _2258_ _3627_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
X_4688_ _1236_ _1241_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_160_379 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4127__A2 _0742_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6427_ _1458_ _2806_ _2807_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_113_262 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6358_ _1455_ _2740_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_11_282 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_112_1858 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_228_653 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5309_ core_0.execute.alu_mul_div.div_cur\[8\] _1756_ _1757_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_6289_ _2039_ _2048_ _2629_ _2673_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_0_228_675 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8028_ _0205_ clknet_leaf_56_i_clk net117 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_242_100 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_242_111 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_215_325 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output132_I net132 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_231_829 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_230_317 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_67_1315 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_196_711 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_205_2977 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_168_413 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6052__A2 net203 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_772 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_168_457 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4063__A1 _0567_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_636 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_124 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_149_671 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_183_416 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_109_513 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_123_1987 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_155_118 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_149_682 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_234_3318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_54_606 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_535 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_136_321 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_557 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7552__A2 _1206_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_164_663 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_842 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_191_471 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_81_458 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_124_527 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_136_387 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_10_634 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_50_801 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_152_2339 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_34_363 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_151_346 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_78_1444 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7304__A2 _3391_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6498__B _2286_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_104_240 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_34_396 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_201_86 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_61_193 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5315__A1 core_0.execute.alu_mul_div.div_cur\[4\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_104_251 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_132_571 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_91_1600 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_104_284 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_120_733 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_238_417 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_238_428 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5866__A2 _2257_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7068__A1 core_0.execute.alu_mul_div.mul_res\[9\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_148_Right_148 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_245_3447 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_245_3458 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6815__A1 core_0.ew_reg_ie\[2\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_206_314 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_234_656 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_234_667 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_222_807 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_163_2468 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_89_1584 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_187_722 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_18_723 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_202_531 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_159_424 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7240__A1 net83 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_187_744 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_18_734 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_186_243 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3990_ _0565_ _0524_ _0527_ core_0.execute.rf.reg_outputs\[6\]\[9\] _0620_ vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_0_9_508 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_47 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_57_422 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_282 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_85_731 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7791__A2 _3786_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_202_597 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_146_107 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_71_69 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_242_60 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_84_241 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_242_71 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_466 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_17_308 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_128_855 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_45_628 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5660_ _2055_ _2060_ _2061_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__7543__A2 net19 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_72_447 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4611_ net155 core_0.ew_addr_high\[0\] _1171_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__5554__A1 _0987_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4357__A2 _0942_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5591_ _1990_ _1991_ _1992_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_143_836 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_155_696 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_25_352 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_661 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_143_858 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_174_2597 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_7330_ _1724_ _2328_ _3502_ _3503_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_5_769 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4542_ _1126_ _0002_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_142_357 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7261_ net86 _3398_ _3399_ _3441_ _3442_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__4109__A2 net18 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4473_ _1065_ _1039_ _1066_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_0_111_733 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_40_366 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6212_ _2287_ _1758_ _2420_ _2598_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_111_755 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_229_439 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7192_ _3260_ _3372_ _3381_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_111_766 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_111_788 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_209_3022 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_115_Right_115 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
X_6143_ _2202_ _2529_ _2530_ _0183_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__5609__A2 _1631_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_51_1127 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_237_483 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6074_ _2462_ _2152_ _2148_ _2463_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_2
XANTENNA__4656__B _1214_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_127_2032 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6282__A2 _2294_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5025_ _1472_ _1473_ _1474_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_240_615 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_224_177 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_212_317 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6871__B _3112_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_17_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_136_94 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7231__A1 net82 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_220_350 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_95_539 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_220_361 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6976_ _3175_ _3189_ _3194_ _3195_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__5242__C2 _1690_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_220_383 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_165_416 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5927_ _2300_ _1624_ _2318_ _2319_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_137_129 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_75_263 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_62_1256 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_5858_ net185 _2251_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_180_408 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_75_296 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_180_419 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_17_842 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_161_600 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5545__A1 _1004_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4809_ _0870_ core_0.fetch.submitable _1311_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4348__A2 core_0.decode.i_flush vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_17_Right_17 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_106_527 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_138_2172 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_90_255 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5789_ _2189_ _2190_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_32_801 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_145_184 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_50_119 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7528_ _0580_ _3641_ _3659_ _0439_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_133_368 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_16_396 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7298__A1 _1414_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7207__B _3393_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7459_ _3563_ net76 _3553_ _3612_ _3613_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai211_2
XANTENNA__7298__B2 _1431_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_3_290 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_101_232 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_101_276 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6538__S _2906_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_101_287 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_216_601 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_73_1385 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_26_Right_26 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__6273__A2 _2579_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_216_667 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7470__A1 net37 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_231_604 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5241__I core_0.decode.oc_alu_mode\[6\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4284__A1 core_0.fetch.prev_request_pc\[7\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_231_626 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4284__B2 core_0.fetch.prev_request_pc\[6\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_9_i_clk_I clknet_4_3__leaf_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_240_3388 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7222__A1 _1742_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_219 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_98_399 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_169_777 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_422 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_168_265 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_196_585 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5397__B _1841_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_128_107 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_66_241 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_183_224 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_35_Right_35 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_82_734 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7525__A2 _3646_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_26_127 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6328__A3 _2710_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_109_354 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_217_Right_217 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_81_244 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_125_836 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5536__A1 net81 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6584__I0 core_0.ew_submit vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_124_313 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_136_173 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_23_792 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_125_858 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_81_277 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7289__A1 net74 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_193 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_140_839 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_152_699 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_151_176 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_151_187 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_105_593 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_675 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5839__A2 _2233_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_238_247 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_226_409 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_44_Right_44 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
Xclkbuf_leaf_114_i_clk clknet_4_4__leaf_i_clk clknet_leaf_114_i_clk vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XPHY_EDGE_ROW_152_Left_399 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_237_82 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6264__A2 _2648_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5151__I _1599_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4275__A1 _0892_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_89_311 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_206_177 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_leaf_129_i_clk clknet_4_0__leaf_i_clk clknet_leaf_129_i_clk vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_221_136 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6691__B _3004_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7213__A1 net80 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_159_221 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6830_ _2967_ _3086_ _3094_ _0306_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_77_539 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_106_64 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_75 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_147_405 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_202_383 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4578__A2 net157 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6761_ _2981_ _3042_ _3054_ _0277_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_3973_ _0604_ net196 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XPHY_EDGE_ROW_53_Right_53 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_176_2626 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_18_617 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_174_235 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5712_ _1600_ _2112_ _2113_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_4
XFILLER_0_9_349 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_175_769 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_57_274 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6692_ _2988_ _3000_ _3014_ _0248_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__7516__A2 _3640_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_162_419 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_174_279 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5643_ _2039_ _2043_ _2044_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_128_685 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_73_789 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_31_72 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_14_801 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_5_533 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_94 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_26_683 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_170_441 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5574_ _1980_ _0745_ _0164_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_143_666 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_215_3092 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_198_34 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_41_620 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_5_566 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7313_ _3398_ _3487_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_4525_ core_0.decode.i_instr_l\[3\] core_0.decode.i_instr_l\[2\] _1078_ _1112_ _1113_
+ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_4
XANTENNA__4750__A2 _1241_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_8293_ _0469_ clknet_leaf_12_i_clk core_0.dec_sreg_store vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_142_187 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_664 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7244_ net83 _3413_ net84 _3427_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_4456_ net71 _1051_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_40_185 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_62_Right_62 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_1_772 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_187_2755 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_229_258 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_217_409 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7175_ _3357_ _3371_ _0374_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_4387_ _0959_ _0997_ _0998_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or2_1
X_6126_ _2513_ _2514_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__7452__A1 net37 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_119 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6057_ core_0.execute.sreg_irq_flags.o_d\[4\] _2250_ _2260_ net11 _2446_ vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__4266__A1 core_0.fetch.prev_request_pc\[15\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5008_ core_0.decode.oc_alu_mode\[4\] _1457_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__inv_4
XFILLER_0_96_804 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_197_349 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6007__A2 _2260_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_202_2936 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_95_314 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_71_Right_71 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__7755__A2 _1072_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_221_692 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_93_i_clk clknet_4_6__leaf_i_clk clknet_leaf_93_i_clk vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_95_347 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_178_574 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_198_2884 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6959_ _3154_ _3174_ _3179_ _0350_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_48_241 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_138_449 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_120_1957 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_63_200 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7507__A2 _3640_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_153_419 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_165_279 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_91_553 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_382 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_858 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_146_493 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_20_751 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_63_299 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_642 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_122_839 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_161_496 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_75_1414 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_80_Right_80 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA_clkbuf_leaf_88_i_clk_I clknet_4_12__leaf_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_31_i_clk clknet_4_10__leaf_i_clk clknet_leaf_31_i_clk vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_31_196 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_236_707 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_6_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__7691__A1 _1084_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7691__B2 _1065_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_235_228 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_242_3417 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_235_239 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_4_0__f_i_clk clknet_3_0_0_i_clk clknet_4_0__leaf_i_clk vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
Xclkbuf_leaf_46_i_clk clknet_4_9__leaf_i_clk clknet_leaf_46_i_clk vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__6067__I _2454_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_244_773 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_216_475 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_244_795 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_204_637 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_203_114 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_160_2427 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_160_2438 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_98_141 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_99_664 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_86_1543 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_99_697 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_231_478 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_28_851 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_86_325 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7746__A2 _1062_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_196_371 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_211_180 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_74_509 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_55_712 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_39_274 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_414 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_319 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_82_531 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5509__A1 _1375_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_15_609 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_171_238 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4251__S _0724_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_70_737 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_82_597 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_113_806 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6182__A1 core_0.execute.alu_mul_div.div_res\[6\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_171_2567 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_97_1672 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_4310_ _0898_ _0923_ _0924_ _0927_ _0928_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or4_1
XFILLER_0_168_26 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_2_569 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_10_314 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_168_37 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5290_ core_0.dec_jump_cond_code\[4\] _1738_ core_0.dec_pc_inc _1739_ vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_4
X_4241_ _0824_ net47 _0859_ _0860_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_4
XANTENNA__7682__A1 _1037_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_160_Left_407 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_120_382 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_226_217 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4172_ _0787_ _0788_ _0790_ _0791_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_2
XANTENNA__7434__A1 _3547_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_93_34 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4248__A1 _0865_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_184_69 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_124_2002 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_117_41 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7931_ _0109_ clknet_leaf_14_i_clk core_0.execute.sreg_long_ptr_en vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_2
XTAP_TAPCELL_ROW_182_2696 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_222_445 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4799__A2 _1237_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_117_85 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_89_174 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_222_489 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_188_861 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7862_ _0054_ clknet_leaf_71_i_clk core_0.fetch.prev_request_pc\[5\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__4653__C _0731_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5748__A1 _2018_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6813_ core_0.execute.rf.reg_outputs\[3\]\[15\] _3063_ _3083_ _3084_ vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_187_393 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_92_306 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7793_ core_0.decode.i_instr_l\[15\] _3786_ _3802_ core_0.decode.i_instr_l\[12\]
+ _1133_ _3858_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XTAP_TAPCELL_ROW_46_1059 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_106_1790 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7737__S _1063_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5212__A3 _0778_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_92_317 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_148_769 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_217_3121 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_9_146 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6744_ _1963_ _3045_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
X_3956_ _0585_ _0586_ _0587_ _0588_ _0589_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_0_175_566 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_46_767 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_778 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6675_ _2956_ _2999_ _3005_ _0240_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_3887_ core_0.dec_r_reg_sel\[1\] _0523_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_73_575 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_45_277 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5626_ _2010_ _2011_ _2027_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_135_2131 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6173__A1 _1600_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_115_154 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_171_772 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_60_247 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_839 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_103_316 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_130_102 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_143_485 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5557_ core_0.execute.mem_stage_pc\[12\] _1955_ _1964_ _1974_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__5920__A1 _1482_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_143_496 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4723__A2 _1237_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_170_282 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_450 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_103_349 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_41_472 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4508_ _1040_ core_0.decode.i_instr_l\[2\] _1044_ _1084_ _1098_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_4
X_8276_ _0452_ clknet_leaf_26_i_clk core_0.execute.pc_high_out\[5\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_2
X_5488_ _1230_ _1920_ _1921_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA_input56_I i_req_data[26] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7673__A1 _1034_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7227_ _3406_ _3407_ _3412_ _0385_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_4439_ _1033_ _1034_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_218_729 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_57_1199 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_228_3250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8015__CLK clknet_leaf_53_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4487__A1 _1056_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7158_ core_0.execute.alu_mul_div.div_res\[2\] _3360_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_70_1355 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6109_ _2244_ _2496_ _2497_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_6_579 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7425__A1 core_0.execute.sreg_irq_pc.o_d\[7\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7089_ _1225_ _3248_ _3298_ _1222_ _3299_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_0_225_261 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_198_603 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5720__S _1554_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_109_1819 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_146_2260 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_198_625 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_241_743 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5987__A1 _2300_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8165__CLK clknet_leaf_89_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5987__B2 _1624_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_174_91 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_197_146 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_325 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_25_810 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_84_807 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_96_667 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_138_202 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_369 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5739__A1 _1439_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_139_736 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_166_522 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_712 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6400__A2 _1114_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_193_352 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4411__A1 core_0.fetch.prev_request_pc\[3\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_154_739 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_81_1484 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_153_216 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4962__A2 _0615_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_51_203 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_107_644 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_190 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_52_737 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6164__A1 core_0.decode.oc_alu_mode\[4\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5394__C _1838_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_51_247 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_161_282 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4714__A2 _1237_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_32_472 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_121_146 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_667 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6467__A2 net214 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7664__A1 _3663_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4478__A1 _1038_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_208_228 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7416__A1 _3547_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6219__A2 _2133_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_223_209 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4493__A4 _1085_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_188_102 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5978__A1 _1559_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_3_1_0_i_clk_I clknet_0_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4246__S _0724_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_314 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_87_623 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_188_168 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_169_360 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_200_640 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_185_842 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_74_317 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_86_177 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_27_200 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_129_257 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4790_ _1290_ _1299_ _0061_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_117_408 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_99_1701 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_27_244 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4953__A2 _1394_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_144_238 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_103_76 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_31_879 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_82_383 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6460_ _2078_ _2083_ _2084_ _2839_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_2
XANTENNA__6155__A1 _2403_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_111_i_clk_I clknet_4_4__leaf_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_153_772 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_42_247 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5411_ core_0.execute.alu_mul_div.div_cur\[6\] _1812_ _1841_ _1854_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_212_3051 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_88_34 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_112_102 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_113_636 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_212_3062 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_42_269 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6391_ _2062_ _2066_ _2071_ _2772_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_112_113 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_180_591 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput103 net103 dbg_r0[9] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
X_8130_ _0306_ clknet_leaf_111_i_clk core_0.execute.rf.reg_outputs\[2\]\[5\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xoutput114 net114 o_instr_long_addr[6] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_11_623 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5342_ core_0.execute.alu_mul_div.div_cur\[10\] _1789_ _1790_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__xor2_1
Xoutput125 net125 o_mem_addr[3] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_23_494 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_2_366 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput136 net136 o_mem_addr_high[4] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
Xoutput147 net147 o_mem_data[2] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
Xoutput158 net158 o_mem_sel[1] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA__6458__A2 _2486_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_8061_ _0237_ clknet_leaf_94_i_clk core_0.execute.rf.reg_outputs\[6\]\[0\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_2
XANTENNA__7655__A1 _1078_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput169 net169 o_req_addr[2] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
X_5273_ _1480_ _1700_ _1721_ _1722_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or3_2
XTAP_TAPCELL_ROW_130_2072 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5604__I _1652_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_227_526 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7012_ core_0.execute.alu_mul_div.cbit\[3\] _3227_ _3228_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_10_177 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_184_2725 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_4224_ net54 core_0.fetch.out_buffer_data_instr\[24\] _0824_ _0843_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_4
XFILLER_0_195_57 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5130__A2 _1492_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_227_559 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7407__A1 net204 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_128_51 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4155_ _0773_ _0769_ _0774_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_235_570 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_3_549 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_207_294 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4086_ _0704_ _0705_ _0706_ _0707_ _0708_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_0_97_409 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_223_3191 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_36_i_clk_I clknet_4_11__leaf_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_39_979 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6630__A2 _2972_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7914_ _0005_ clknet_leaf_120_i_clk core_0.decode.oc_alu_mode\[2\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_179_157 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_78_634 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_78_645 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4641__A1 net193 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_66_807 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_78_667 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7845_ _0038_ clknet_leaf_64_i_clk core_0.fetch.out_buffer_data_instr\[22\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_144_94 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_187_190 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_19_723 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_195_2854 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6394__A1 _2300_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_93_648 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_175_352 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_46_520 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7776_ core_0.dec_rf_ie\[2\] _3766_ _3833_ _3848_ _3849_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_46_531 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4988_ _0770_ _0773_ _0769_ _1437_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_0_46_553 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_19_767 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_244 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6727_ core_0.execute.rf.reg_outputs\[5\]\[10\] _3027_ _3031_ _3035_ vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_190_333 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3939_ _0568_ core_0.execute.rf.reg_outputs\[4\]\[13\] _0520_ _0573_ vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA__4944__A2 _1394_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_190_344 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xwire219 _1483_ net219 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_116_430 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_737 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_650 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6658_ _2979_ core_0.ew_data\[14\] _2980_ net26 _2994_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_0_6_683 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_59_1217 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_131_411 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5609_ _1693_ _1631_ _2010_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_4
XFILLER_0_33_269 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6697__A2 _3000_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_131_422 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_143_282 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_5_182 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6589_ _2930_ _2937_ _2938_ _2939_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_2
X_8328_ _0504_ clknet_leaf_89_i_clk core_0.dec_r_reg_sel\[0\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_output162_I net162 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7646__A1 net115 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6449__A2 _2827_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_115_1889 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_8259_ _0435_ clknet_leaf_36_i_clk core_0.execute.sreg_scratch.o_d\[9\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5121__A2 _1435_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6546__S _2906_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_205_209 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4880__A1 core_0.decode.i_imm_pass\[15\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_214_732 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_213_220 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_214_765 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_241_562 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_623 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_201_415 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_68_111 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_158_308 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_83_1513 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_185_138 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_wire211_I _1718_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_167_842 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_56_317 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_68_177 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_56_328 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_204_53 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_194_661 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_127_706 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_83_125 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_49_391 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_154_514 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_37_553 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_83_158 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_204_97 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_64_361 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput16 i_core_int_sreg[9] net16 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_24_214 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_52_523 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6137__A1 core_0.execute.alu_mul_div.div_cur\[5\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput27 i_mem_data[15] net27 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_91_180 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_236 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_135_772 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput38 i_req_data[0] net38 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_24_247 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_80_865 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput49 i_req_data[1] net49 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_12_409 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6688__A2 _2999_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_134_282 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_94_1642 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_32_280 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_122_488 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7637__A1 _3732_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_37 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_20_453 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_236_323 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_229_72 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5112__A2 _1492_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6964__B _1651_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_224_518 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6860__A2 _3107_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_217_570 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_166_2499 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_205_743 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_189_422 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3879__I core_0.dec_r_reg_sel\[2\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_0_508 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_220_702 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_189_444 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5960_ _2347_ _2348_ _2349_ _2350_ _2351_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_0_189_488 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_181_26 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_36_949 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_48_807 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_4911_ _1369_ _1231_ _1223_ _1376_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_176_127 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5891_ _2004_ _2282_ _2283_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_142_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__7168__A3 _1230_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4704__S _1246_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7630_ _0733_ _3729_ _3743_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_59_188 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6376__A1 _1379_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_185_661 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_47_339 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5179__A2 _1436_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4842_ _1280_ net43 _1170_ _1332_ _1333_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_0_28_531 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_43_1029 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_28_553 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7561_ core_0.execute.pc_high_buff_out\[1\] _3682_ _3684_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4773_ core_0.fetch.prev_request_pc\[4\] _1285_ _0881_ net171 _1291_ vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_0_117_238 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_249 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_16_737 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_99_33 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6128__A1 _2300_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_28_597 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6512_ _1088_ _2888_ _2889_ _0799_ _2890_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_0_130_30 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7492_ core_0.execute.sreg_jtr_buff.o_d\[2\] _1208_ _3638_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_132_2101 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6679__A2 _3006_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_153_580 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6443_ _2798_ _2822_ _1114_ _2823_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_113_422 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_125_282 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_190_2795 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_130_74 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_141_742 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6374_ _2754_ _2755_ _2756_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_30_239 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_140_252 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5351__A2 _1702_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_8_608 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_2_174 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7628__A1 core_0.execute.pc_high_buff_out\[2\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_8113_ _0289_ clknet_leaf_111_i_clk core_0.execute.rf.reg_outputs\[3\]\[4\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5325_ _1767_ _1771_ _1772_ _1773_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XANTENNA__3901__A3 _0536_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_228_835 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_475 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4378__C _0963_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6300__A1 _2626_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5256_ _1513_ _1514_ _1515_ _1516_ _1705_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_4
XTAP_TAPCELL_ROW_54_1158 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_139_72 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8044_ _0220_ clknet_leaf_49_i_clk net155 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_47_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_215_507 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4207_ _0824_ _0825_ _0826_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6851__A2 _3087_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5187_ _0776_ _1633_ _1634_ _1635_ _1636_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai211_4
XFILLER_0_208_592 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_242_348 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4138_ core_0.execute.next_ready_delayed _0757_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_143_2230 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_223_551 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_3_72 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_input19_I i_mc_core_int vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_223_562 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_211_702 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6603__A2 core_0.ew_data\[2\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7800__A1 _1039_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4069_ _0532_ _0523_ _0526_ _0692_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_0_211_735 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3968__A3 _0543_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_149_842 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_167_138 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_317 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4090__A2 _0535_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_78_497 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_148_341 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7828_ _0021_ clknet_leaf_53_i_clk core_0.fetch.out_buffer_data_instr\[5\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__6367__A1 _2281_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8203__CLK clknet_leaf_2_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_164_801 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_66_659 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_65_1287 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_65_1298 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_81_607 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_564 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7759_ _1045_ _1071_ _1101_ core_0.decode.i_instr_l\[3\] _3834_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_0_34_512 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_74_681 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_46_383 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_190_152 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6119__A1 _1999_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_163_366 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_117_772 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_123_208 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5590__A2 _1541_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_129_Right_129 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_151_528 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_865 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_104_400 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_117_1918 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_104_411 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5953__B _2190_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_578 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_104_422 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_132_731 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5342__A2 _1789_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_132_797 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_output87_I net87 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7619__A1 net194 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_219_824 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6784__B _3057_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_246_676 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6842__A2 _3092_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_206_529 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4853__A1 _0860_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_242_860 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_201_212 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_97_762 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6070__A3 _1721_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_97_784 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_33_908 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_56_103 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4081__A2 _0594_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_139_330 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_clkbuf_4_4__f_i_clk_I clknet_3_2_0_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_151_18 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_56_125 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_56_136 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_167_683 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_167_694 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_127_536 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4908__A2 _1367_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5030__A1 _1467_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_13_665 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_71_139 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_107_260 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_181_174 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_154_399 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_13_718 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_40_504 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_107_282 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_52_375 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_40_537 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_12_228 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_122_241 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_397 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_548 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_69_69 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5333__A2 _1758_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6530__A1 _2576_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4541__B1 _1064_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_110_447 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_209_301 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5154__I _1596_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_168_2528 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_237_632 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5110_ _1558_ _1559_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XANTENNA__3895__A2 _0530_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_176_37 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6090_ _1433_ _2477_ _2478_ _0799_ _2479_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_0_236_131 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5041_ core_0.execute.rf.reg_outputs\[7\]\[13\] net234 _1435_ core_0.execute.rf.reg_outputs\[6\]\[13\]
+ _1489_ _1490_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_0_85_68 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_29_Left_276 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__6833__A2 _3092_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4844__A1 core_0.decode.i_instr_l\[15\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4695__I1 net65 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_224_359 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_109_86 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_205_562 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5103__B _1460_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6597__A1 _2930_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8226__CLK clknet_leaf_8_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_220_521 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_220_3150 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6992_ _1665_ _3209_ _3210_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_149_105 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5943_ core_0.execute.sreg_irq_pc.o_d\[1\] _2264_ _2265_ core_0.execute.alu_flag_reg.o_d\[1\]
+ _2258_ core_0.execute.trap_flag _2335_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XANTENNA__4072__A2 _0529_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_179_2657 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6713__I _3020_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6349__A1 _2294_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_87_294 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_101_1719 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_158_661 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_136 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5874_ _2255_ _2259_ _2261_ _2266_ _2267_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_0_164_119 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_192_2813 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_7613_ _1209_ _2249_ _3729_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_4
XPHY_EDGE_ROW_38_Left_285 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
X_4825_ _0937_ core_0.decode.i_instr_l\[10\] _1305_ _1320_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_173_642 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_709 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_394 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7544_ _3663_ _3668_ _0446_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__5572__A2 _0743_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4756_ _1051_ _1279_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_172_163 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_865 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6869__B _3112_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_191 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_160_325 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_172_185 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_114_731 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_126_591 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4687_ _0817_ _1237_ _1240_ _0017_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_7475_ core_0.execute.sreg_jtr_buff.o_d\[0\] _1398_ _3626_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_231_3290 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6426_ _2076_ _2805_ _2806_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA_rebuffer11_I net232 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_31_559 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5324__A2 _1600_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6521__A1 _1381_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_250 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6357_ _1137_ _1568_ _1061_ _2739_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_228_621 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_59_91 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_112_1859 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_5308_ _1503_ _1504_ _1756_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_4
XPHY_EDGE_ROW_47_Left_294 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
X_6288_ _2298_ _2666_ _2671_ _2672_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_4
XANTENNA__5088__A1 _0789_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_216_827 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8027_ _0204_ clknet_leaf_53_i_clk net131 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__6824__A2 _3087_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5239_ _1137_ _1451_ _1061_ _1688_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_166_81 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_231_808 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_205_2967 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_67_1316 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
Xclone1 net222 net221 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XANTENNA__6588__A1 net21 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_205_2978 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7785__B1 _3827_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_196_734 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_79_784 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4063__A2 _0524_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_66_401 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5260__A1 core_0.decode.oc_alu_mode\[12\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_103 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_211_598 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_39_648 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_78_294 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_123_1988 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_195_288 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_109_525 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_183_439 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_234_3319 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_191_450 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_53_128 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_93_297 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6760__A1 core_0.execute.rf.reg_outputs\[4\]\[8\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_62_640 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_62_651 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_10_635 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_117_591 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_163_196 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_clkbuf_leaf_5_i_clk_I clknet_4_2__leaf_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_375 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_61_161 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_78_1445 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_22_559 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5315__A2 _1695_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6512__A1 _1088_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_91_1601 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_104_296 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_120_745 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_581 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_219_632 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_120_778 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_219_654 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_245_3448 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5079__A1 _1467_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_219_687 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6815__A2 _2934_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_206_337 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_233_134 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_206_359 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_89_504 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_215_860 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_163_2469 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6579__A1 _2242_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_89_559 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_89_1585 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_214_381 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7776__B1 _3833_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_18_724 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_202_543 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_710 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_97_570 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_37 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_159_469 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_85_743 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_128_801 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_85_754 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_29_158 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_127_322 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_242_83 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5003__A1 _1123_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_489 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_5_704 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_44_139 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4610_ _1170_ core_0.fetch.submitable vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
X_5590_ _1713_ _1541_ _1991_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__7792__C _1279_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5554__A2 _1956_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_26_865 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6689__B _3004_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_142_325 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_154_185 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_759 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4541_ _1124_ _1062_ _1064_ _1125_ _1126_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_TAPCELL_ROW_174_2598 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_108_591 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_4_247 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_312 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_170_667 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_52_172 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_142_369 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7260_ _3439_ _3440_ _3441_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__6503__A1 _2123_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4472_ core_0.decode.i_instr_l\[0\] _1065_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__inv_3
XFILLER_0_229_418 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6211_ _1831_ _2594_ _2596_ _2412_ _2597_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai211_2
X_7191_ _1748_ _3380_ _0381_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_40_389 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_96_45 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_21_570 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_110_244 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_209_3023 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6142_ core_0.ew_data\[5\] _2486_ _2530_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_237_451 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_209_142 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4937__B _1284_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_51_1128 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6073_ _1695_ _1929_ _2462_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6806__A2 _3070_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_224_101 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_94 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5024_ core_0.dec_alu_carry_en core_0.execute.alu_flag_reg.o_d\[1\] _1473_ vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_127_2033 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_213_819 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_240_605 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4293__A2 _0835_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5490__A1 net217 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_178_701 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_177_200 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7231__A2 _3398_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_67_209 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_178_745 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6975_ _2386_ _3192_ _3193_ _3194_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor3_1
XANTENNA__5242__A1 _1686_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5242__B2 _1689_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_88_592 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5926_ _2317_ _2318_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_177_277 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_445 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5793__A2 _1606_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_118_300 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_177_288 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_177_299 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_8_520 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_158_480 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_118_322 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_192_247 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_62_1257 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_75_275 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_91_724 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5857_ net186 _1201_ _1383_ _2250_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and3_2
XFILLER_0_63_426 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_146_664 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4808_ _1045_ core_0.fetch.submitable _1310_ _0068_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__5545__A2 _1956_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_133_314 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_138_2173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_5788_ _1051_ _1953_ _2189_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_0_8_597 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7527_ core_0.execute.sreg_scratch.o_d\[13\] _3646_ _3651_ _3659_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_44_673 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4739_ _0831_ _1238_ _1270_ _0039_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_31_301 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_183 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7458_ net37 _3611_ _3612_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6409_ net75 _2531_ _2789_ _2537_ _2790_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XPHY_EDGE_ROW_55_Left_302 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_101_222 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_4_10__f_i_clk_I clknet_3_5_0_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7389_ _3547_ _3554_ _3555_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_12_592 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_101_299 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_73_1386 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4808__A1 _1045_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5076__A4 _1524_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_243_465 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4284__A2 _0833_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_230_104 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_215_178 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6554__S _2906_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_240_3389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_224_690 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_64_Left_311 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA_clkbuf_leaf_84_i_clk_I clknet_4_12__leaf_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_169_756 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4036__A2 core_0.dec_r_reg_sel\[1\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5233__A1 core_0.decode.oc_alu_mode\[1\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_169_767 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_168_255 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_79_592 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_169_789 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_196_597 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6981__A1 _1226_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_184_737 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_456 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_765 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_184_748 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_489 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_81_212 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_181_Right_181 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__5536__A2 _1953_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6584__I1 net20 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_23_793 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_140_807 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_152_667 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_172 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_312 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4601__I _1165_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_73_Left_320 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_105_583 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_10_507 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_132_391 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_120_597 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_66_37 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_219_484 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4249__S _0724_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_246_292 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_207_668 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7461__A2 _3542_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_237_94 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4275__A2 _0837_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_173_16 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_203_830 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_159_200 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7213__A2 net79 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_209 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_106_32 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_202_340 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_77_529 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_159_233 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3887__I core_0.dec_r_reg_sel\[1\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5224__A1 _0771_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_721 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_187_575 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6760_ core_0.execute.rf.reg_outputs\[4\]\[8\] _3049_ _3045_ _3054_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_57_220 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_147_417 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3972_ _0597_ _0602_ _0603_ _0604_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_4
XTAP_TAPCELL_ROW_176_2627 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_48_1090 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_73_702 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_562 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5711_ _1123_ _2111_ _2112_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_174_247 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_222_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6691_ core_0.execute.rf.reg_outputs\[6\]\[11\] _3006_ _3004_ _3014_ vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_45_437 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_116_804 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_45_448 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_128_675 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5642_ _2042_ _2043_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__6724__A1 _2981_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_73_768 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_183_781 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_115_314 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_115_336 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_170_431 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_31_84 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_545 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5573_ _1980_ _0748_ _0163_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_215_3093 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_7312_ _1395_ _3486_ _0396_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_41_632 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_53_492 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_130_317 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4524_ _1065_ _1039_ _1112_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_8292_ _0468_ clknet_leaf_10_i_clk core_0.dec_sreg_jal_over vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__dffq_4
XFILLER_0_41_676 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7243_ net84 net83 _3413_ _3426_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and3_1
X_4455_ _1037_ _1042_ _1044_ _1049_ _1050_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_229_226 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_40_197 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_187_2756 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5160__B1 _1434_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4386_ _0889_ _0951_ _0997_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_7174_ _3261_ _3355_ core_0.execute.alu_mul_div.div_res\[7\] _3371_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_6125_ _1690_ _2010_ _2511_ _1631_ _2512_ _2513_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_0_147_72 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6056_ core_0.execute.sreg_priv_control.o_d\[4\] _1385_ _2265_ core_0.execute.alu_flag_reg.o_d\[4\]
+ _2445_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_198_807 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4266__A2 _0827_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_212_104 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_106_i_clk_I clknet_4_5__leaf_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5007_ _1131_ _1455_ _1456_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_0_240_435 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_240_457 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_202_2937 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_49_710 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_721 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_163_60 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_138_406 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6958_ core_0.execute.alu_mul_div.mul_res\[0\] _3177_ _3178_ _1451_ _3179_ vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__6963__A1 _1439_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_166_737 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_198_2885 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_49_765 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_178_597 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_193_556 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5909_ _1559_ _1689_ _2301_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_2
XTAP_TAPCELL_ROW_120_1947 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_119_642 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_120_1958 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6889_ _2996_ _3108_ _3127_ _0332_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_64_746 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_134_601 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_826 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_17_640 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6715__A1 _2961_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_63_256 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_106_314 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_119_697 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_134_623 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6566__I1 core_0.ew_reg_ie\[3\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output192_I net192 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_20_752 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_122_807 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_134_667 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__8094__CLK clknet_leaf_109_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_16_183 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_16_194 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_133_166 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_120 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_75_1415 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_31_142 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_114_391 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7140__A1 _1364_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_102_597 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_235_207 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_242_3418 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7443__A2 _3542_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6792__B _3072_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_610 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_231_402 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_203_104 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6284__S _1819_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_632 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_188_317 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_160_2428 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_87_816 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_86_1544 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_86_304 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_28_852 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5206__A1 _0771_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_212_682 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_196_383 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_184_523 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_242 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_702 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_67_562 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_223_63 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_156_247 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_67_584 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_39_286 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_172_729 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_184_589 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_55_757 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_82_543 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6706__A1 _2940_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_42_407 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6182__A2 _1114_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_35_492 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_23_632 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_171_2568 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_2_515 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_112_317 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_22_131 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_97_1673 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_2_537 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_239_502 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_23_687 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3940__A1 _0534_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_239_557 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4240_ core_0.fetch.out_buffer_valid _0858_ _0859_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_227_719 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_120_394 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4171_ core_0.ew_reg_ie\[4\] _0783_ _0789_ _0790_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_184_37 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_172_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_93_57 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_124_2003 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_7930_ _0108_ clknet_leaf_23_i_clk core_0.execute.sreg_data_page vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_234_284 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_182_2697 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_222_435 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5996__A2 _2386_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_89_142 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_222_457 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7861_ _0053_ clknet_leaf_71_i_clk core_0.fetch.prev_request_pc\[4\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_26_95 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_77_326 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_187_361 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6812_ _1963_ _3083_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XANTENNA__5748__A2 _2022_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6945__A1 _1915_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_93_819 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7792_ _0542_ _1134_ _3857_ _1279_ _0505_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_148_737 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_175_523 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_58_551 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_106_1780 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_46_702 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_217_3111 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6743_ _2940_ _3042_ _3044_ _0269_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_217_3122 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_3955_ _0534_ _0535_ _0536_ core_0.execute.rf.reg_outputs\[6\]\[12\] _0588_ vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_0_45_212 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_163_718 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_73_532 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_18_448 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_116_601 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_128_461 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_18_459 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6674_ core_0.execute.rf.reg_outputs\[6\]\[3\] _3000_ _3004_ _3005_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3886_ core_0.execute.rf.reg_outputs\[2\]\[15\] _0522_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_61_716 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5625_ _1999_ _2009_ _2016_ _2025_ _2026_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai211_4
XTAP_TAPCELL_ROW_135_2132 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_6_865 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_104_807 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_115_133 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_116_667 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_60_226 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_54_790 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4184__A1 core_0.decode.o_submit vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_103_306 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_643 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_131_626 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5556_ _0982_ _1956_ _1973_ _0153_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_41_440 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_32_i_clk_I clknet_4_10__leaf_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5920__A2 _1620_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6877__B _3112_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_13_142 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_77_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_41_462 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4507_ _1093_ _1096_ _1097_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_8275_ _0451_ clknet_leaf_26_i_clk core_0.execute.pc_high_out\[4\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_13_175 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5487_ _1226_ _1568_ _1919_ _1920_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_7226_ _3384_ _3411_ _3412_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5133__B1 _1443_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7673__A2 _3773_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4438_ _0721_ _1032_ _1033_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_245_516 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5684__A1 _2078_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input49_I i_req_data[1] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_228_3251 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_7157_ _2331_ _3359_ _3357_ _0368_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_4369_ _0934_ _0942_ _0945_ _0854_ _0983_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_0_226_752 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_70_1356 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6108_ _2455_ _2495_ _2496_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__7425__A2 _3543_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7088_ _1224_ _3297_ _3298_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_146_2261 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7501__B _3516_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6039_ _2425_ _2428_ _2429_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_241_755 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_197_136 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_213_468 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7189__A1 _1748_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_95_101 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_200_107 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5021__B _1451_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output205_I net205 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_25_811 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_95_134 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6936__A1 _1915_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5739__A2 _1448_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_194_832 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_193_320 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_37_702 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_49_562 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_194_865 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_193_331 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_138_247 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_239_3380 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_83_329 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_113_i_clk clknet_4_4__leaf_i_clk clknet_leaf_113_i_clk vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_153_206 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_543 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_81_1485 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_92_863 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_133 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7361__A1 _2565_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_17_492 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4151__I core_0.dec_l_reg_sel\[2\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4175__A1 _0789_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_106_177 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_128_i_clk clknet_4_0__leaf_i_clk clknet_leaf_128_i_clk vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__7113__A1 _1226_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4478__A2 _1039_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5911__S _1482_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6219__A3 _2604_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_217_796 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7411__B _3546_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_244_593 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5978__A2 _1555_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_231_232 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_204_457 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_231_254 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_86_112 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_348 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_3_5_0_i_clk_I clknet_0_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6927__A1 core_0.decode.o_submit vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_28_713 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_184_342 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_157_567 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_212 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_184_364 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_554 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_99_1702 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7727__I0 net192 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7352__A1 core_0.execute.alu_flag_reg.o_d\[3\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_153_762 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_70_535 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_179_26 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5410_ core_0.execute.alu_mul_div.div_cur\[5\] _1814_ _1817_ _1852_ _1853_ vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_113_615 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_42_259 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_568 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_212_3052 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_23_440 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6390_ _2287_ _2067_ _2080_ _1690_ _2770_ _2771_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai221_4
XFILLER_0_23_451 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_113_648 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_334 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_140_434 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput104 net104 o_c_data_page vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
Xoutput115 net115 o_instr_long_addr[7] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
X_5341_ _1508_ _1509_ _1789_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_0_10_101 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput126 net126 o_mem_addr[4] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_100_309 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput137 net137 o_mem_addr_high[5] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_112_169 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput148 net148 o_mem_data[3] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
Xoutput159 net159 o_mem_we vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA__5115__B1 _1443_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_8060_ _0236_ clknet_leaf_98_i_clk core_0.execute.rf.reg_outputs\[7\]\[15\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__7655__A2 _1072_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5272_ _1123_ _1451_ net211 _1720_ _1721_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai211_4
Xclkbuf_leaf_92_i_clk clknet_4_6__leaf_i_clk clknet_leaf_92_i_clk vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_121_692 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_130_2073 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5666__A1 _1803_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_184_2715 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_7011_ _3225_ _3226_ _1366_ _3227_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4223_ _0726_ _0840_ _0841_ _0842_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XPHY_EDGE_ROW_10_Left_257 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_184_2726 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_10_189 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_208_730 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_195_69 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4154_ core_0.dec_l_reg_sel\[1\] _0773_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__inv_4
XANTENNA__7407__A2 _3544_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_208_785 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_207_262 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5418__A1 core_0.execute.alu_mul_div.div_cur\[6\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_37_72 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_83 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4085_ _0567_ _0524_ _0527_ core_0.execute.rf.reg_outputs\[2\]\[1\] _0707_ vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_4
XTAP_TAPCELL_ROW_223_3192 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_7913_ _0004_ clknet_leaf_9_i_clk core_0.decode.oc_alu_mode\[1\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_222_265 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_222_276 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_179_169 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_77_123 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4641__A2 net180 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_210_438 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_148_501 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7844_ _0037_ clknet_leaf_65_i_clk core_0.fetch.out_buffer_data_instr\[21\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xclkbuf_leaf_30_i_clk clknet_4_10__leaf_i_clk clknet_leaf_30_i_clk vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__6918__A1 _2988_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_702 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_93_627 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_176_865 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_195_2855 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_7775_ core_0.decode.i_instr_l\[7\] _3847_ _3848_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__7591__A1 _3682_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_18_212 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_381 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6394__A2 _1560_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4987_ _0770_ _0778_ _1436_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_4
XFILLER_0_148_578 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6726_ _2983_ _3021_ _3034_ _0262_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_18_234 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_74_863 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3938_ core_0.execute.rf.reg_outputs\[7\]\[13\] _0530_ _0572_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_160_61 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_46_587 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_727 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_128_291 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_45_i_clk clknet_4_9__leaf_i_clk clknet_leaf_45_i_clk vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_160_83 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6146__A2 _1385_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_73_384 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6657_ _2941_ _2992_ _2993_ _0234_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_6_662 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_160_94 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_59_1218 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_5608_ _2003_ _2007_ _2008_ _2009_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_4
X_6588_ net21 _1150_ _2938_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_14_451 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_103_136 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_42_782 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_8327_ _0503_ clknet_leaf_80_i_clk core_0.dec_rf_ie\[7\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5539_ _1963_ _1964_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_41_270 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8258_ _0434_ clknet_leaf_36_i_clk core_0.execute.sreg_scratch.o_d\[8\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__7646__A2 _3729_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_112_681 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8132__CLK clknet_leaf_111_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_218_527 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_111_180 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7209_ _2390_ _3391_ _3395_ _3396_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA_output155_I net155 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_100_865 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8189_ _0365_ clknet_leaf_127_i_clk core_0.execute.alu_mul_div.mul_res\[15\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_214_711 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5409__A1 _1233_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_185_80 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6457__I0 _0580_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_226_582 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4880__A2 _1341_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_241_541 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8282__CLK clknet_leaf_29_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6082__A1 _1831_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_241_552 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_101 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_214_799 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_83_1503 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_83_1514 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_213_298 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6562__S _1985_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_201_449 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_96_454 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6909__A1 net101 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_84_605 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_189 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3985__I _0615_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_204_65 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_83_137 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_204_76 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_532 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_193_183 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_126_239 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_92_671 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_64_384 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput17 i_disable net17 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6137__A2 _1432_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput28 i_mem_data[1] net28 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
Xinput39 i_req_data[10] net39 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_80_855 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_107_486 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_40_719 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_162_592 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5896__A1 _2287_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7406__B _3546_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_150_765 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_94_1643 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_110_607 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_60_590 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_150_798 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_20_465 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_237_836 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_237_858 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6964__C core_0.execute.alu_mul_div.cbit\[0\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_74_37 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_74_48 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4871__A2 _1321_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_217_593 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_205_755 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6999__I1 _3215_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6073__A1 _1695_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_0_509 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_245_72 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_205_788 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_245_94 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5820__A1 _2202_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4623__A2 core_0.execute.alu_flag_reg.o_d\[2\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_36_939 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_59_134 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4910_ _1374_ _1375_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_220_769 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_605 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5890_ _1643_ _1476_ _2282_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_87_476 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_74_104 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_90_69 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_158_865 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4841_ _0726_ _1259_ _1332_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_173_802 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_103_1750 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_114_65 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_135_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7573__A1 _3673_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_117_206 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4387__A1 _0959_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_74_148 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_200_493 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7560_ core_0.execute.pc_high_out\[1\] core_0.execute.pc_high_out\[0\] _3683_ vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_56_863 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_184_172 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4772_ _1283_ _1290_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_145_548 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_576 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_727 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6511_ core_0.execute.alu_mul_div.i_mul core_0.execute.alu_mul_div.mul_res\[15\]
+ _2889_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_71_833 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7491_ _0732_ _3637_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__inv_1
XANTENNA__7325__A1 _2711_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_82_170 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_82_181 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_70_332 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_99_67 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4139__A1 _0535_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_31_708 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6442_ _2281_ _2821_ _2822_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_132_2102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_31_719 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_190_2796 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_125_294 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_120 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_70_387 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_131 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6373_ core_0.execute.sreg_scratch.o_d\[11\] _2579_ _2534_ net3 _2755_ vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_113_478 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_8_609 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_101_629 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_2_164 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8112_ _0288_ clknet_leaf_94_i_clk core_0.execute.rf.reg_outputs\[3\]\[3\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__7628__A2 _3731_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5324_ core_0.execute.alu_mul_div.div_cur\[2\] _1600_ _1772_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_2_197 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_100_139 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5639__A1 _1756_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_487 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8043_ _0013_ clknet_leaf_17_i_clk core_0.decode.i_flush vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__dffq_4
XTAP_TAPCELL_ROW_54_1159 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_5255_ _1507_ _1512_ _1517_ _1519_ _1704_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and4_2
XTAP_TAPCELL_ROW_225_3210 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6300__A2 _2672_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_227_346 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4206_ core_0.fetch.out_buffer_data_instr\[31\] _0825_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_48_93 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_227_379 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_243_839 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5186_ core_0.execute.rf.reg_outputs\[6\]\[4\] _1434_ _1437_ core_0.execute.rf.reg_outputs\[2\]\[4\]
+ _1635_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XANTENNA__4862__A2 _1306_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4137_ core_0.decode.i_flush _0755_ _0756_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__4394__C _0963_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_143_2231 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6064__A1 _1378_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7261__B1 _3399_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_155_72 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__7800__A2 _1048_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4068_ _0532_ _0541_ _0543_ _0691_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_0_78_410 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5811__A1 net133 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_168_629 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6382__S _2190_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_307 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4090__A3 _0536_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7827_ _0020_ clknet_leaf_61_i_clk core_0.fetch.out_buffer_data_instr\[4\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__7564__A1 core_0.execute.pc_high_out\[1\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_521 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_532 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6998__S0 core_0.execute.alu_mul_div.cbit\[0\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_65_1288 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4378__A1 _0987_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_236_3350 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_65_159 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_19_554 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_93_468 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7758_ core_0.decode.i_instr_l\[9\] _1132_ _3833_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_191_632 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_163_323 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6709_ core_0.execute.rf.reg_outputs\[5\]\[2\] _3022_ _3016_ _3025_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_34_524 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6119__A2 _2009_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_73_170 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7316__A1 _1400_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_535 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7689_ _3786_ _3788_ _3789_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_62_855 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7316__B2 _1430_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_73_192 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_117_1919 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_154_2360 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5878__A1 core_0.dec_sreg_jal_over vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_30_741 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_774 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_219_836 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_218_313 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_219_858 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_234_817 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_245_154 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4853__A2 _1306_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_233_349 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_1_i_clk_I clknet_4_2__leaf_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_202_703 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_199_765 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_199_776 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_410 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4605__A2 core_0.ew_mem_width vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_198_264 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_69_432 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_198_275 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_33_909 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_29_318 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_201_268 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_96_284 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7555__A1 net194 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_155_824 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4604__I core_0.ew_addr\[0\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_127_526 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_38_863 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_166_172 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4908__A3 _1227_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_166_194 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_502 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5030__A2 net213 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_65_682 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_13_666 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_181_142 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__7307__A1 net76 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_142_507 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_154_378 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_170_827 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_123_710 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_135_570 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_80_663 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_181_186 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_69_26 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_69_37 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_527 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_123_776 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6530__A2 _2334_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_122_275 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_79_i_clk_I clknet_4_13__leaf_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4541__A1 _1124_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4392__I1 _0833_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4541__B2 _1125_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_168_2529 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_209_346 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6294__A1 core_0.decode.oc_alu_mode\[2\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5097__A2 net232 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_209_368 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5040_ _1487_ _1488_ _1489_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_225_839 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_109_54 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4844__A2 _1307_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_205_530 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_189_220 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_79_207 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7094__I0 core_0.execute.alu_mul_div.mul_res\[11\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_192_37 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_79_218 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_195_Right_195 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
X_6991_ _3149_ _1819_ _3209_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_4
XTAP_TAPCELL_ROW_220_3151 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6597__A2 core_0.ew_data\[1\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_88_730 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7794__A1 _0539_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_189_275 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_220_533 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5942_ core_0.execute.alu_mul_div.div_cur\[1\] _2279_ _2330_ _2333_ _2334_ vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai22_4
XFILLER_0_149_139 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_47_104 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_179_2658 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_75_424 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7546__A1 _1209_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5873_ core_0.execute.sreg_irq_pc.o_d\[0\] _2264_ _2265_ core_0.execute.alu_flag_reg.o_d\[0\]
+ _2266_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_0_118_504 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7612_ _3722_ _3673_ _3728_ _1217_ _0454_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_185_470 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_158_684 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_192_2814 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_145_312 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4824_ _1319_ _0075_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_185_492 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_7_212 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_173_632 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_118_548 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_62_107 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5021__A2 _1469_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_62_118 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_524 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7543_ core_0.execute.irq_en net19 _1398_ core_0.execute.sreg_irq_flags.o_d\[4\]
+ _3668_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_4755_ _0825_ _1238_ _1278_ _0047_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_28_384 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_172_153 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_16_535 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_209 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_44_855 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_161_838 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4780__A1 _1290_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_71_663 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7474_ _3581_ _3625_ _0419_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_172_197 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4686_ net49 _1238_ _1240_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_160_348 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_43_376 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_70_162 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_231_3280 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6425_ _2081_ _2774_ _2805_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_70_195 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_141_562 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6521__A2 core_0.execute.sreg_irq_pc.o_d\[15\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4389__C _0877_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_113_275 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4532__A1 _1034_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6356_ _2055_ _2737_ _2738_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_11_262 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5307_ core_0.execute.alu_mul_div.div_cur\[9\] _1754_ _1755_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_227_121 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6287_ _2090_ _2667_ _2670_ _2671_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_2
X_8026_ _0203_ clknet_leaf_56_i_clk net130 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5238_ _1462_ _1469_ _1451_ _1687_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_2
XANTENNA_input31_I i_mem_data[4] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_243_636 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_215_327 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_242_135 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5169_ _0776_ _1614_ _1616_ _1617_ _1618_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__6037__A1 _1137_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_75_91 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_98_527 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xclone2 _0671_ net227 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlyc_4
XTAP_TAPCELL_ROW_205_2968 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_67_1317 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_162_Right_162 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_168_404 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_output118_I net118 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_196_746 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4063__A3 _0527_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_182_92 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_115 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_195_278 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_123_1989 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_66_457 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_136_301 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_176_492 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_93_276 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_94_799 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_148_194 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_164_643 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_559 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_163_131 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_47_682 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_163_142 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_124_518 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6760__A2 _3049_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_191_484 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4771__A1 _1284_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_10_636 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_62_663 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_201_66 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_22_527 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_78_1446 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_104_231 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_105_754 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_34_387 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_34_398 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_201_99 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6512__A2 _2888_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_80_i_clk_I clknet_4_13__leaf_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_91_1602 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_30_593 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_245_3449 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6276__A1 net87 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5079__A2 net182 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6276__B2 _2537_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_219_699 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4287__B1 _0838_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_218_187 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_233_124 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_206_349 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6028__A1 _2412_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_202_500 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_187_702 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_89_1575 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6579__A2 _2202_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_199_562 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_214_371 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_89_1586 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_226_85 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_18_725 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_230_853 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_159_437 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_202_555 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_187_768 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5251__A2 _1600_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_424 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7528__A1 _0580_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_29_126 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_85_766 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_608 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_155_632 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_167_492 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_107 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5003__A2 core_0.decode.oc_alu_mode\[13\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_84_276 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_427 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_154_131 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_154_142 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_182_451 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_26_855 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_25_321 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_727 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_182_473 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4540_ _1066_ _1056_ _1101_ _1041_ _1125_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XTAP_TAPCELL_ROW_174_2599 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_52_140 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_41_836 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_25_387 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_4_259 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_858 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_123_562 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4471_ _1063_ _1064_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA__7700__B2 _3799_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6210_ net223 _2414_ _2595_ _1765_ _2596_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_0_0_410 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4514__A1 _1055_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7190_ _3369_ _3372_ core_0.execute.alu_mul_div.div_res\[14\] _3380_ vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_110_234 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6141_ _2346_ net227 _2528_ _2529_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_209_3024 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7380__I net37 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6267__A1 _2650_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6072_ _2013_ _2460_ _2461_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_29_84 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_51_1129 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5114__B _0779_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5023_ _1470_ _1471_ _1472_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_127_2034 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_213_809 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7216__B1 _3399_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_224_157 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5490__A2 _1650_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_45_72 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_221_842 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_221_853 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_94 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_177_212 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6974_ _1925_ _1927_ core_0.execute.alu_mul_div.cbit\[3\] core_0.execute.alu_mul_div.cbit\[2\]
+ _3193_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XFILLER_0_95_519 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_221_864 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_220_341 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5925_ _1596_ _2313_ _2316_ _2317_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_76_733 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_232 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_118_312 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_479 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5856_ _2248_ _2249_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_158_492 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_62_1258 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_3_Right_3 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
X_4807_ _0869_ core_0.fetch.submitable _1310_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_28_170 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_161_602 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5787_ _2184_ _2187_ _2188_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_2
XANTENNA__6742__A2 _3043_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_138_2163 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_138_2174 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_7526_ _0592_ _3641_ _3658_ _0438_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_4738_ net53 _1253_ _1270_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_44_663 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_160_123 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_102_i_clk_I clknet_4_7__leaf_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_16_387 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_151_2330 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_7457_ core_0.execute.mem_stage_pc\[13\] _3611_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_4669_ _1224_ _1225_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
X_6408_ _2787_ _2788_ _2789_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_EDGE_ROW_2_Left_249 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_101_212 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4505__A1 _1041_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_102_757 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_141_392 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7388_ core_0.execute.mem_stage_pc\[1\] _3554_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_3_292 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_231_Right_231 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
X_6339_ _1379_ _2721_ _2722_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__5803__I _2201_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_216_603 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_73_1387 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_216_625 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4269__B1 _0830_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_243_422 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4808__A2 core_0.fetch.submitable vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_8009_ _0186_ clknet_leaf_55_i_clk core_0.ew_data\[8\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_215_135 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_215_146 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_99_836 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_99_858 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_169_702 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_243_499 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7758__A1 core_0.decode.i_instr_l\[9\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_193_80 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_27_i_clk_I clknet_4_10__leaf_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_168_212 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_86_519 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_98_379 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_169_746 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_211_352 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6430__A1 _2293_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5233__A2 _1124_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_66_221 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_168_278 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_211_396 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6981__A2 _1676_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_156_429 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4154__I core_0.dec_l_reg_sel\[1\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6570__S _2201_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_183_226 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4992__A1 _0770_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_183_237 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_39_479 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_149_492 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_107 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_94_585 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6194__B1 _2579_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6733__A2 _3027_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_164_473 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_23_783 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_137_698 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_191_270 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_652 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_23_794 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_152_635 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_124_337 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_81_279 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_124_348 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_23_836 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_90_780 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_105_540 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_35_696 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_551 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_858 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_105_562 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_120_510 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_699 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_219_430 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_157_18 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_207_603 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_89_302 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5472__A2 _1814_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7749__A1 core_0.decode.i_instr_l\[9\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_199_370 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_203_842 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_159_212 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7213__A3 net72 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_700 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_89_379 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_207_Left_454 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__4027__A3 net231 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_230_683 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_733 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3971_ net90 _0578_ _0603_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_174_215 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5710_ _1596_ _1481_ _2111_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_2
XTAP_TAPCELL_ROW_176_2628 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_48_1091 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6690_ _2986_ _3000_ _3013_ _0247_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_73_714 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_574 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5641_ _2040_ _2041_ _2042_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_127_142 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_215_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6724__A2 _3021_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7375__I _3541_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_5_513 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_652 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_142_101 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_72_268 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5572_ _1980_ _0743_ _0162_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_122_98 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_5_557 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_780 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_215_3094 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_7311_ _3409_ _3481_ _3485_ _3486_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_5_568 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4523_ _1110_ _1111_ _0012_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_8291_ _0467_ clknet_leaf_11_i_clk core_0.dec_sreg_irt vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_4
XPHY_EDGE_ROW_216_Left_463 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_142_189 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7242_ _3420_ _3421_ _3425_ _0387_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_229_205 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_111_532 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4454_ _1046_ _1048_ _1049_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_0_0_240 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_7173_ _3357_ _3370_ _0373_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_4385_ net86 _0996_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XTAP_TAPCELL_ROW_187_2757 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5160__B2 core_0.execute.rf.reg_outputs\[6\]\[6\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_390 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6124_ _1061_ _1693_ _2151_ _1109_ _2512_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_6055_ _2444_ _0181_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5006_ _1452_ _1453_ _1454_ _1455_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_4
XANTENNA__6660__A1 _2941_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XPHY_EDGE_ROW_225_Left_472 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_221_650 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_202_2938 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_96_839 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_163_72 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6957_ _3175_ _1689_ _3178_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_0_220_171 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7883__CLK clknet_leaf_83_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_198_2886 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_48_232 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6963__A2 _1448_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_76_552 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_159_790 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_405 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_714 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5908_ _1641_ _2300_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_119_632 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_120_1948 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4974__A1 _1419_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_91_500 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6888_ core_0.execute.rf.reg_outputs\[1\]\[15\] _3106_ _3124_ _3127_ vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_64_725 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_224 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5839_ _0177_ _2233_ _2234_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_134_613 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6715__A2 _3021_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_107_838 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_384 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_91_566 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_161_410 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4726__A1 net46 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_63_279 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_118_197 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_348 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_20_753 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_234_Left_481 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_161_454 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_44_482 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA_output185_I net185 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7509_ net227 _3648_ _3649_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_75_1416 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6479__A1 core_0.execute.alu_mul_div.div_res\[14\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_114_381 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_31_154 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5961__C core_0.dec_sreg_irt vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_32_699 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_839 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_188_80 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_130_863 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_229_772 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_216_400 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_242_3419 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4149__I _0767_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6100__B1 _2257_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_243_Left_490 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__6651__A1 _2941_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_231_414 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_160_2429 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_203_138 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_86_1545 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_200_801 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_28_853 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6403__A1 _2360_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5206__A2 _0773_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_200_823 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_129_418 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_552 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_156_237 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_109_142 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_223_97 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_235 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_55_769 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6313__B _1457_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6706__A2 _3021_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_124_101 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_137_484 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4612__I _1171_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_192_590 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_588 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_482 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_152_465 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_2_505 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5390__A1 _1747_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_140_616 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_171_2569 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_2_527 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_62_290 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_97_1674 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_50_452 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3940__A2 _0535_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_23_699 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5142__A1 net102 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_10_349 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_120_384 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5693__A2 _2092_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_207_400 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4170_ _0782_ _0789_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XANTENNA__6983__B core_0.execute.alu_mul_div.cbit\[1\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_219_282 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_234_241 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_207_477 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_93_47 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_124_2004 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6642__B2 net36 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_93_69 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_179_307 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3898__I _0533_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4653__B1 _1211_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_182_2698 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_117_65 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_165_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_7860_ _0052_ clknet_leaf_62_i_clk core_0.fetch.prev_request_pc\[3\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_78_839 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6811_ _2994_ _3065_ _3082_ _0299_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_148_716 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7791_ core_0.decode.i_instr_l\[14\] _3786_ _3802_ core_0.decode.i_instr_l\[11\]
+ _1133_ _3857_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_0_147_204 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6945__A2 _1702_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_106_1781 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6742_ core_0.execute.rf.reg_outputs\[4\]\[0\] _3043_ _3031_ _3044_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_217_3112 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4956__B2 _1391_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_46_714 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_137 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_500 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_3954_ _0539_ core_0.execute.rf.reg_outputs\[4\]\[12\] _0520_ _0587_ vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_18_416 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__7319__B _3384_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6673_ _1963_ _3004_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_46_769 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3885_ _0517_ _0520_ _0521_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_4
XANTENNA__6223__B _2279_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_61_706 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_257 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_155_270 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_33_408 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5624_ _2021_ _2024_ _2025_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_183_590 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_45_279 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_6_855 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_73_599 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_135_2133 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_5_343 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_238 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_115_156 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_170_251 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5555_ core_0.execute.mem_stage_pc\[11\] _1955_ _1964_ _1973_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__4184__A2 core_0.execute.alu_mul_div.i_mul vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5381__A1 _1233_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_130_104 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4506_ _1043_ _1094_ _1095_ _1083_ _1096_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_2
X_8274_ _0450_ clknet_leaf_23_i_clk core_0.execute.pc_high_out\[3\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_2
X_5486_ _1226_ _1501_ _1919_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_130_159 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_112_863 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7225_ net81 _3408_ _3410_ _3411_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4437_ _0812_ _1031_ _1032_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_0_111_384 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_228_3252 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_7156_ _1369_ _1227_ _1364_ _3358_ _3359_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_4368_ net74 _0982_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XPHY_EDGE_ROW_92_Left_339 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__6893__B _3124_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_238_591 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_226_731 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6107_ _2494_ _2495_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__inv_1
XTAP_TAPCELL_ROW_70_1357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6385__S _2113_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7087_ _1229_ _3275_ _3296_ _3297_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4299_ core_0.fetch.prev_request_pc\[0\] _0851_ _0914_ core_0.fetch.prev_request_pc\[1\]
+ core_0.fetch.prev_request_pc\[2\] _0860_ _0917_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai222_4
XFILLER_0_226_786 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6633__A1 _2929_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_146_2262 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6038_ _1997_ _2426_ _2427_ _1831_ _1686_ _2428_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_0_197_104 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_240_244 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_68_305 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_197_148 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_69_839 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_83_91 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_200_119 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_194_811 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_96_658 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4247__I0 net65 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_25_812 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6936__A2 _1559_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7989_ _0166_ clknet_leaf_20_i_clk core_0.execute.sreg_irq_flags.i_d\[2\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_166_524 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output100_I net100 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_138_226 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_166_535 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_178_395 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8061__CLK clknet_leaf_94_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_239_3381 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4947__B2 _1391_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_193_354 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_64_522 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_76_382 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_166_579 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7229__B net82 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6133__B _2520_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_81_1486 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5528__I _1955_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_64_555 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_153_229 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4432__I _0748_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_257 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_9_693 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_91_352 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_119_484 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_24_419 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_181 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_162_741 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_157_2391 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_45_780 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_107_668 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7361__A2 _2606_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_134_465 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5372__A1 core_0.execute.alu_mul_div.div_cur\[0\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3922__A2 _0528_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7113__A2 _1491_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_636 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5124__A1 _0782_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_130_671 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_102_384 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_47_18 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6872__A1 _2977_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_102_395 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_217_742 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_216_241 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6624__A1 _2936_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_5_570 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_188_104 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_232_745 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_231_244 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3989__A2 _0594_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_231_277 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6027__C _1831_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_327 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_86_124 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_231_299 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_197_682 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6927__A2 _1088_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_234_85 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_196_170 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_86_168 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_200_664 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_55_500 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_157_557 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_200_675 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_45_1050 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_55_533 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_842 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_6_107 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_55_544 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_99_1703 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_103_34 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_172_527 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_184_387 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_55_566 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_27_268 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_15_419 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_125_432 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7352__A2 _3510_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5363__A1 _1374_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_152_251 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4166__A2 core_0.execute.sreg_long_ptr_en vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_23_430 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_302 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_212_3053 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_35_290 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_836 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_3_858 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_51_772 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5340_ _1755_ _1757_ _1786_ _1787_ _1788_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai211_4
Xoutput105 net105 o_c_instr_long vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_88_69 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_EDGE_ROW_149_Left_396 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
Xoutput116 net116 o_mem_addr[0] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
Xoutput127 net127 o_mem_addr[5] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_50_271 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput138 net138 o_mem_addr_high[6] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_140_479 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_10_124 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput149 net149 o_mem_data[4] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
X_5271_ core_0.decode.oc_alu_mode\[12\] _1719_ _1720_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_4
XTAP_TAPCELL_ROW_130_2074 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_239_377 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7010_ _2001_ _1665_ _1929_ _1631_ _1226_ _1228_ _3226_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux4_2
X_4222_ _0726_ net46 _0841_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_10_168 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6863__A1 _2956_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5666__A2 _1500_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_184_2716 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_56_1190 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7602__B _3672_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_208_753 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_207_230 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4153_ _0768_ _0769_ _0771_ _0772_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_235_550 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_128_64 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6615__A1 _2930_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5418__A2 _1838_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_223_723 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_222_200 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4084_ _0517_ core_0.execute.rf.reg_outputs\[4\]\[1\] net229 _0706_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_2
XTAP_TAPCELL_ROW_108_1810 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_179_104 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6091__A2 _2332_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4517__I core_0.decode.oc_alu_mode\[4\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_223_767 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_223_3193 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_222_244 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7912_ _0103_ clknet_leaf_81_i_clk core_0.decode.i_jmp_pred_pass vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__8084__CLK clknet_leaf_109_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_78_614 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_194_107 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_188_660 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4641__A3 net179 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7843_ _0036_ clknet_leaf_65_i_clk core_0.fetch.out_buffer_data_instr\[20\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_78_658 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_203_480 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_194_129 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_72 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6918__A2 _3130_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_187_170 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_148_535 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4929__A1 _1392_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_176_855 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_77_179 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4986_ _1434_ _1435_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_148_557 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7774_ _1317_ _3842_ _3847_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_175_343 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_195_2856 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_46_511 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_18_202 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6394__A3 _2642_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6725_ core_0.execute.rf.reg_outputs\[5\]\[9\] _3027_ _3031_ _3034_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3937_ _0568_ _0542_ _0544_ core_0.execute.rf.reg_outputs\[1\]\[13\] _0571_ vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_0_191_836 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_19_769 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_191_858 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_73_352 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_18_268 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_6_630 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_514 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6656_ core_0.execute.rf.reg_outputs\[7\]\[13\] _2962_ _2984_ _2993_ vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__6888__B _3124_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5607_ _1676_ _1600_ _2008_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_30_870 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6587_ net35 _1148_ _2937_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_59_1219 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_42_750 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_8326_ _0502_ clknet_leaf_81_i_clk core_0.dec_rf_ie\[6\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5538_ _0722_ _1963_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XANTENNA_input61_I i_req_data[30] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_8257_ _0433_ clknet_leaf_32_i_clk core_0.execute.sreg_scratch.o_d\[7\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_112_671 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5469_ core_0.execute.alu_mul_div.div_cur\[15\] _1711_ _1807_ _1903_ vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_7208_ _3392_ _3394_ _3395_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_100_855 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4704__I1 net69 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_8188_ _0364_ clknet_leaf_127_i_clk core_0.execute.alu_mul_div.mul_res\[14\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_245_336 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7139_ _1915_ net214 _3344_ _1364_ _3345_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XANTENNA_output148_I net148 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_226_561 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6606__A1 net23 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7803__B1 _3866_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_226_594 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_214_734 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_214_745 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_241_531 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_2_540 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_241_564 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_198_457 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4093__A1 _0568_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_113 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_83_1504 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_38_970 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5459__S _1373_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6909__A2 _3135_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7031__A1 _1908_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_157 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_166_310 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_159_2420 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_139_557 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_182_803 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_77_691 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_127_719 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_65_842 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_166_365 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4396__A2 _0950_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_154_527 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_166_387 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4162__I core_0.dec_l_reg_sel\[2\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_182_858 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_37_588 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_363 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput18 i_irq net18 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__6798__B _3072_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_91_171 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_135_763 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput29 i_mem_data[2] net29 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__5345__A1 core_0.execute.alu_mul_div.div_cur\[11\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_709 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_772 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5896__A2 _1603_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_94_1644 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_150_777 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_103_660 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_103_671 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_236_303 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6845__A1 _2990_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_477 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_176_Right_176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_244_380 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7270__A1 net87 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_205_767 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6073__A2 _1929_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4084__A1 _0517_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_260 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_232_575 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87_422 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_99_282 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_232_597 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_220_737 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_176_107 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_clkbuf_leaf_75_i_clk_I clknet_4_13__leaf_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_157_310 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_47_319 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4840_ core_0.decode.i_instr_l\[14\] _1307_ _1331_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_87_488 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_511 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_157_343 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_28_522 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_103_1751 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_28_533 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_145_516 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4771_ _1284_ _1289_ _0052_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_7_416 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_145_527 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_184_162 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_609 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_128_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_184_184 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_352 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6510_ _2886_ _2887_ _2888_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_0_173_858 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_672 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_15_205 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_83_683 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7490_ _3635_ _3636_ _1284_ _0424_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_70_311 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_172_357 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7325__A2 _2734_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_130_32 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_172_379 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6441_ _2802_ _2804_ _2807_ _2820_ _2821_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XANTENNA__4139__A2 _0536_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_157_Left_404 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_43_558 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_113_413 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_190_2797 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_30_208 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_141_755 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6372_ core_0.execute.sreg_priv_control.o_d\[11\] _1386_ _2577_ core_0.execute.sreg_irq_pc.o_d\[11\]
+ _2754_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_140_232 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_130_98 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_23_271 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_140_254 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7089__A1 _1225_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_23_282 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_8111_ _0287_ clknet_leaf_109_i_clk core_0.execute.rf.reg_outputs\[3\]\[2\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5323_ _1768_ _1769_ _1770_ _1771_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_4
XFILLER_0_100_107 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_228_804 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_140_298 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6836__A1 _2981_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_8042_ _0219_ clknet_leaf_47_i_clk core_0.ew_mem_width vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_2
X_5254_ _1701_ _1702_ _1703_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_TAPCELL_ROW_114_1880 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_239_196 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_143_Right_143 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_225_3211 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_4205_ core_0.fetch.out_buffer_valid _0824_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
Xclkbuf_leaf_112_i_clk clknet_4_4__leaf_i_clk clknet_leaf_112_i_clk vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_5185_ core_0.execute.rf.reg_outputs\[1\]\[4\] _1615_ _1436_ core_0.execute.rf.reg_outputs\[4\]\[4\]
+ net219 _1634_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi221_4
X_4136_ core_0.execute.hold_valid core_0.decode.o_submit _0755_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XPHY_EDGE_ROW_166_Left_413 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_208_594 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7261__A1 net86 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6064__A2 core_0.execute.sreg_irq_pc.o_d\[4\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_143_2232 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5111__I1 _1555_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4067_ net96 _0690_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__inv_2
XFILLER_0_3_96 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7800__A3 _1069_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_127_i_clk clknet_4_1__leaf_i_clk clknet_leaf_127_i_clk vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_64_93 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5811__A2 _2209_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_210_247 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7013__A1 core_0.execute.alu_mul_div.mul_res\[5\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
X_7826_ _0019_ clknet_leaf_58_i_clk core_0.fetch.out_buffer_data_instr\[3\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_19_511 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7564__A2 _3672_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_93_436 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_47_831 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_47_842 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_65_1289 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_171_72 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_175_151 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_236_3340 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5575__A1 _1980_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4378__A2 _0966_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_148_376 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_609 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_108_218 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7757_ _3831_ _3832_ _1284_ _0495_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_136_527 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_148_387 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4969_ _1381_ _0592_ _1422_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_108_229 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6708_ _2946_ _3021_ _3024_ _0254_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XPHY_EDGE_ROW_175_Left_422 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_74_694 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7688_ _1098_ _1099_ _3787_ _3788_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_4
XANTENNA__7316__A2 core_0.execute.sreg_irq_pc.o_d\[15\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_116_251 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_144_571 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6639_ _2979_ core_0.ew_data\[8\] _2980_ net35 _2981_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XTAP_TAPCELL_ROW_154_2361 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_144_593 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_772 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5878__A2 _2270_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_104_457 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6130__C _1831_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_104_468 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_591 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8309_ _0485_ clknet_leaf_75_i_clk net179 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_4
XANTENNA__6827__A1 core_0.execute.rf.reg_outputs\[2\]\[4\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_100_630 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_100_663 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_110_Right_110 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_234_807 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6637__I _2929_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_184_Left_431 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_233_339 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_165_2490 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7252__A1 _1414_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7252__B2 _1431_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_198_254 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_69_422 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_214_597 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_202_737 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5697__B net211 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_202_748 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_69_444 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_158_107 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7004__A1 _1637_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_96_252 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5015__B1 _0692_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_60_18 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_leaf_91_i_clk clknet_4_6__leaf_i_clk clknet_leaf_91_i_clk vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__7555__A2 _3675_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_56_138 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_84_447 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4369__A2 _0942_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_193_Left_440 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__5566__A1 _1977_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_182_611 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_154_313 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_42_1020 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5917__S _1603_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_53_801 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4908__A4 _1230_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_155_858 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_182_644 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_71_119 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_300 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7307__A2 _3467_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_13_667 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_65_694 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_154_368 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_245_Right_245 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_25_536 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_142_519 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_108_774 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7417__B _3553_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5318__A1 core_0.execute.alu_mul_div.div_cur\[3\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_135_593 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_181_198 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5869__A2 _1382_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_49 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_0_614 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_100_57 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4541__A2 _1062_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_241 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_85_26 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6294__A2 _1585_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_85_48 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_236_155 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_224_317 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7243__A1 net84 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4067__I net96 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6990_ _3198_ _3206_ _3207_ _3208_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__7794__A2 _1134_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_232_372 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_220_3152 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_5941_ _2331_ _2332_ _2279_ _2333_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA__7378__I _3541_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_245_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_220_567 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_88_786 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5872_ net186 _1198_ _1201_ _2265_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and3_4
XTAP_TAPCELL_ROW_179_2659 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_59_i_clk clknet_4_14__leaf_i_clk clknet_leaf_59_i_clk vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__7546__A2 _2257_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7611_ _3675_ _3726_ _3727_ _3673_ _3728_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_29_842 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_118_516 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4823_ _0936_ core_0.decode.i_instr_l\[9\] _1305_ _1319_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_192_2815 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8122__CLK clknet_4_7__leaf_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_28_341 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_145_346 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4754_ net62 _1241_ _1278_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_56_683 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7542_ _3663_ _3667_ _0445_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_50_51 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_90_439 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_173_688 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_212_Right_212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_43_333 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5309__A1 core_0.execute.alu_mul_div.div_cur\[8\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_173_699 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_160_327 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7473_ core_0.execute.sreg_irq_pc.o_d\[15\] _3542_ _3624_ _3625_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4685_ _0814_ _1237_ _1239_ _0016_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_160_338 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8272__CLK clknet_leaf_26_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_114_755 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_174 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6424_ _1457_ _2803_ _2804_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_2
XTAP_TAPCELL_ROW_231_3281 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_12_720 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_731 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_113_265 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_114_799 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_12_753 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6355_ _2698_ _2060_ _2064_ _2737_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__4532__A2 _1116_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_3_496 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_113_298 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5306_ _1753_ _1754_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XANTENNA__6809__A1 _2992_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6286_ _2294_ _2669_ _2670_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_52_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_228_667 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_227_133 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_216_807 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_8025_ _0202_ clknet_leaf_38_i_clk net129 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5237_ core_0.decode.oc_alu_mode\[9\] _1686_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__inv_3
XFILLER_0_216_829 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4296__A1 _0824_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_215_317 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5168_ core_0.execute.rf.reg_outputs\[4\]\[7\] _1436_ _1437_ core_0.execute.rf.reg_outputs\[2\]\[7\]
+ _1617_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_224_840 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_input24_I i_mem_data[12] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_208_391 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__7234__A1 _3409_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6037__A2 _1931_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4119_ core_0.execute.pc_high_out\[0\] net105 _0739_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_5099_ _1544_ _1545_ _1546_ _1547_ _1548_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and4_2
XTAP_TAPCELL_ROW_67_1318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_205_2969 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7785__A2 _1133_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_223_383 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_79_753 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5796__A1 _2187_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_78_285 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_94_734 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_149_663 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_505 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_19_330 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_94_767 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7809_ _1038_ _1094_ _3870_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_93_255 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_136_313 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_137_836 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_94_789 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_136_335 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_137_858 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_191_430 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_417 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_160 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4220__A1 _0835_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_47_694 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_163_176 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_10_637 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_105_722 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_61_152 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_78_1447 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_105_766 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output92_I net92 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_201_89 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_clkbuf_leaf_23_i_clk_I clknet_4_8__leaf_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_104_276 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_120_725 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_238_409 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_91_1603 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6568__S _2201_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_219_612 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_218_111 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_218_133 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6276__A2 _2531_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7473__A1 core_0.execute.sreg_irq_pc.o_d\[15\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_219_678 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_234_626 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_206_317 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_218_177 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7225__A1 net81 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_89_1576 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_202_512 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7776__A2 _3766_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_187_725 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_18_726 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_186_213 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_202_545 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_186_224 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6316__B _1121_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_97_550 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7198__I _1209_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_230_865 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_97_572 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_85_723 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7528__A2 _3641_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_174_419 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_138 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_233 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_195_780 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_458 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_100_1710 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_38_661 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_84_288 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_127_346 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8295__CLK clknet_leaf_88_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_37_160 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4211__A1 _0723_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7147__B _3189_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_25_344 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_111_34 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_170_647 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_80_461 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_174 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_697 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4470_ _1033_ _1063_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_4
XANTENNA__7700__A2 _1134_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_150_360 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5711__A1 _1123_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_111_747 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7661__I _1132_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6140_ _2497_ _2527_ core_0.dec_mem_access _2528_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_0_444 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_209_3025 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_195_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7464__A1 net37 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6071_ _2425_ _2423_ _1997_ _2460_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XTAP_TAPCELL_ROW_51_1119 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_111_1850 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_5022_ _1462_ _1469_ _1450_ _1471_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or3_2
XTAP_TAPCELL_ROW_127_2035 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7216__A1 net80 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_224_169 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_221_832 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_45_84 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5778__A1 _1713_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6973_ _3154_ _3190_ _3191_ _3192_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_178_747 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4825__I0 _0937_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_88_572 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5924_ _1559_ _2315_ _2316_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__7519__A2 _3646_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_76_745 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_177_279 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_119_836 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5855_ net186 _1383_ _2247_ _2248_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_0_61_72 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_91_715 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_62_1259 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_63_417 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_119_858 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_173_430 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_233_3310 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6740__I _3041_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_61_94 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4806_ _0944_ _1306_ _1309_ _0067_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_16_311 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5786_ _2185_ _2186_ _2187_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_2
XTAP_TAPCELL_ROW_138_2164 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7057__B _3175_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_134_839 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7525_ core_0.execute.sreg_scratch.o_d\[12\] _3646_ _3651_ _3658_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_160_102 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4737_ _1269_ _0038_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4753__A2 _1238_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5950__A1 _1378_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_133_349 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_31_303 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_151_2320 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_7456_ _3581_ _3610_ _0416_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_4668_ core_0.execute.alu_mul_div.cbit\[2\] _1224_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_31_347 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6407_ core_0.execute.sreg_scratch.o_d\[12\] _2579_ _2534_ net4 _2788_ vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_4599_ _1164_ net143 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_3_282 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7387_ _3540_ _3553_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XANTENNA__8018__CLK clknet_leaf_24_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_12_561 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6338_ net73 _2531_ _2720_ _2537_ _2721_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_12_594 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_101_268 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6258__A2 _2642_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_177_82 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6269_ _2346_ _2653_ _2654_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_73_1388 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4269__A1 core_0.fetch.prev_request_pc\[12\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4269__B2 core_0.fetch.prev_request_pc\[13\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_216_637 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_8008_ _0185_ clknet_leaf_55_i_clk core_0.ew_data\[7\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_2
XANTENNA__7207__A1 _1195_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_243_467 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_243_489 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_162_2460 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7758__A2 _1132_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_224_692 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_193_92 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_98_358 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_212_865 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4435__I core_0.decode.i_flush vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_169_769 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_39_414 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_168_268 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_183_205 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_149_460 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_184_739 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4992__A2 _0767_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_81_203 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_346 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5694__C _2092_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_82_737 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_94_597 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_82_748 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_19_171 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_236 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_212_66 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_23_784 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_136_165 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_151_102 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_164_485 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5941__A1 _2331_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50_601 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_163 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4170__I _0782_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_117_390 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_22_314 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_34_174 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_151_179 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_105_574 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_667 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7694__A1 _1055_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_112_Left_359 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_132_371 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_120_522 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_120_577 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7446__A1 _3547_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6097__I _2201_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6249__A2 _2633_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_101_780 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_207_615 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_206_103 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7430__B _3545_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_13_Right_13 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_234_489 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7749__A2 _1032_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4680__A1 _0721_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_121_Left_368 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_230_651 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4345__I _0877_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5224__A3 _0779_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_187_566 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3970_ _0598_ _0599_ _0600_ _0601_ _0602_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_0_175_706 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_202_375 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_230_695 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_159_279 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_176_2629 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_168_791 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_48_1092 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_127_132 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6185__A1 _2360_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_45_439 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5640_ _1758_ _1619_ _2041_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_31_42 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_72_236 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_247 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_116_839 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_122_66 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_183_783 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_170_411 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5571_ _1980_ _0733_ _0161_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XPHY_EDGE_ROW_22_Right_22 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__5932__A1 _2322_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_26_664 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5176__I _1482_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_110_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_182_282 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_675 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_143_658 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_208_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_41_612 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7310_ _0964_ _3482_ _3484_ _3485_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_4522_ _1042_ _1095_ _1078_ _1064_ _1111_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai211_2
XPHY_EDGE_ROW_130_Left_377 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_215_3095 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_198_37 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_25_185 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8290_ _0466_ clknet_leaf_10_i_clk core_0.dec_sys vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_40_122 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_142_168 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_80_291 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7241_ _3384_ _3424_ _3425_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4453_ core_0.decode.i_instr_l\[6\] _1047_ core_0.decode.i_instr_l\[5\] _1048_ vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or3_4
XFILLER_0_40_155 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4499__A1 _1038_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_111_555 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7172_ _3358_ _3369_ core_0.execute.alu_mul_div.div_res\[6\] _3370_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_111_566 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4384_ _0991_ _0966_ _0994_ _0995_ _0877_ net176 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_0_40_199 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5160__A2 _1608_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_187_2758 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6123_ _1137_ _1693_ _1456_ _2511_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_0_274 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6054_ core_0.ew_data\[3\] _2443_ _2190_ _2444_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XPHY_EDGE_ROW_31_Right_31 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__5999__A1 _2388_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5005_ core_0.decode.oc_alu_mode\[1\] core_0.decode.oc_alu_mode\[6\] core_0.decode.oc_alu_mode\[7\]
+ core_0.decode.oc_alu_mode\[4\] _1454_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_0_56_83 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6660__A2 _2994_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_212_139 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_96_807 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_15_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_202_2939 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_49_712 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7070__C1 _3178_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_221_673 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6956_ _3176_ _3177_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_3
XFILLER_0_72_71 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_88_380 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_198_2887 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_49_767 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_165_216 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5907_ _2296_ _2298_ _2299_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_48_255 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_76_564 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_9_842 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_120_1949 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6887_ _2994_ _3108_ _3126_ _0331_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_48_277 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_76_597 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_40_Right_40 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_36_439 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5838_ _2227_ _2231_ _2230_ _2233_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_0_119_699 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_174_794 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4726__A2 _1253_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5923__A1 _1554_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_161_422 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_173_282 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5769_ _1510_ _1511_ _2170_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_TAPCELL_ROW_20_754 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_7508_ _3639_ _3648_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_121_319 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_161_488 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7515__B _3651_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_32_667 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_20_807 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_75_1417 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6479__A2 _1114_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7676__A1 _3663_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output178_I net178 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7439_ core_0.execute.mem_stage_pc\[10\] _3596_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_114_393 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7428__A1 _3547_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_235_209 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6100__B2 core_0.execute.pc_high_out\[5\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7250__B _1395_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_612 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6651__A2 _2988_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_216_489 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_204_629 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4662__A1 _1209_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_243_286 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_207_66 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_98_133 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_99_667 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_197_842 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_86_1546 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_28_843 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_86_317 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7600__A1 _3682_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6403__A2 _2783_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_28_854 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_196_352 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4414__A1 _0883_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_200_835 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_211_172 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_184_536 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_715 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_94_361 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_184_569 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_94_383 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_137_441 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_748 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_165_761 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4178__B1 _0765_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_180_720 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_42_409 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5914__A1 _1554_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_125_636 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4717__A2 _1237_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_23_623 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_63_792 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_171_2559 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_180_775 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_124_168 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_140_628 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_442 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_97_1675 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7667__A1 _3663_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_168_18 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3940__A3 _0536_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_121_842 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_10_317 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_239_559 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_22_199 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5142__A2 _1492_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6890__A2 _2934_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_219_261 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_207_445 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_234_231 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6642__A2 core_0.ew_data\[9\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_207_489 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_124_2005 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_179_319 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_182_2699 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4653__B2 _1172_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_78_807 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_222_459 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_158_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_77_328 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6810_ core_0.execute.rf.reg_outputs\[3\]\[14\] _3063_ _3072_ _3082_ vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_187_352 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_89_199 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_202_161 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4405__A1 _1008_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7790_ _0536_ _1134_ _3856_ _1950_ _0504_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XTAP_TAPCELL_ROW_106_1782 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6741_ _3041_ _3043_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA__4956__A2 _1394_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3953_ core_0.execute.rf.reg_outputs\[7\]\[12\] _0530_ _0586_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_217_3113 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6504__B _2090_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_46_737 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_58_597 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_133_76 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_190_506 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_128_452 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6672_ _2951_ _2999_ _3003_ _0239_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_6_801 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3884_ net228 _0520_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_42_96 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_73_556 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5623_ _2022_ _2023_ _2024_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_143_422 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_155_282 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_333 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_206 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_155_293 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_135_2134 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_5554_ _0987_ _1956_ _1972_ _0152_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_103_319 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_14_667 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_13_133 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7658__A1 _1043_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7335__B _3507_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_130_127 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4505_ _1041_ _1071_ _1095_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_5485_ _1364_ _1917_ _1367_ _1918_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_8273_ _0449_ clknet_leaf_22_i_clk core_0.execute.pc_high_out\[2\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_13_166 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_123_190 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7224_ net81 _3408_ _3409_ _3410_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_4436_ core_0.decode.input_valid core_0.decode.i_submit _1030_ _1031_ vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_4
XANTENNA__5133__A2 net232 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6330__A1 _1088_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_111_352 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_228_3253 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_4367_ _0977_ _0966_ _0981_ _0963_ net164 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_4
X_7155_ _1372_ _1809_ _1810_ _3358_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_4
XANTENNA__6881__A2 _3114_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4892__A1 _1280_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6106_ _1378_ _2492_ _2493_ _2494_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_70_1347 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_7086_ _1229_ _3295_ _3296_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_70_1358 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_4298_ core_0.fetch.prev_request_pc\[3\] _0857_ _0860_ core_0.fetch.prev_request_pc\[2\]
+ _0916_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_225_242 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_241_702 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7850__CLK clknet_leaf_68_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_213_404 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6037_ _1137_ _1931_ _1061_ _2427_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_146_2263 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_225_275 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_198_617 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_241_735 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_197_116 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_179_842 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_68_317 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_96_626 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_68_328 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8206__CLK clknet_leaf_129_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7988_ _0165_ clknet_leaf_31_i_clk core_0.execute.prev_pc_high\[7\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_25_813 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_221_492 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4947__A2 _1394_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6939_ _1227_ _1683_ _3160_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_49_575 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_239_3382 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_190_71 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_650 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_147_772 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_193_388 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_247 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_81_1487 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_91_331 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_92_865 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_8_171 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_409 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_162_731 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_206 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_52_729 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_157_2392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_162_753 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_91_386 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_106_157 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_157_Right_157 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__5372__A2 _1819_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_161_263 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_134_488 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_162_797 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7649__A1 _1217_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_32_453 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_103_842 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_60_795 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6872__A2 _3107_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4883__A1 core_0.decode.i_flush vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_217_765 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_217_776 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6624__A2 _2967_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_5_571 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_4_15__f_i_clk clknet_3_7_0_i_clk clknet_4_15__leaf_i_clk vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__4635__A1 core_0.de_jmp_pred vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_231_212 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_188_116 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_99_486 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_169_352 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_200_632 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_129_238 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5060__A1 _1460_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_45_1051 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_184_355 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7139__C _1364_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_82_331 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_99_1704 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_144_219 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_578 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_125_422 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_137_282 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_103_68 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_206 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_125_444 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6155__A4 _2541_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5363__A2 _1809_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_124_Right_124 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_113_628 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_125_488 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_212_3054 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_2_314 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_88_37 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_140_436 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput106 net106 o_c_instr_page vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_11_615 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xoutput117 net117 o_mem_addr[10] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
Xoutput128 net128 o_mem_addr[6] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_2_369 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_clkbuf_leaf_71_i_clk_I clknet_4_13__leaf_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput139 net139 o_mem_data[0] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
X_5270_ _1543_ _1548_ _1719_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or2_4
XANTENNA__5115__A2 net232 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6312__A1 _2633_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4221_ core_0.fetch.out_buffer_data_instr\[17\] _0840_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_120_171 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_130_2075 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_227_518 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6863__A2 _3107_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_227_529 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_184_2717 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_56_1180 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_4152_ _0770_ _0771_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_235_562 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_223_702 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6615__A2 core_0.ew_data\[4\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_37_74 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4083_ core_0.execute.rf.reg_outputs\[7\]\[1\] _0529_ _0705_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_222_212 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_108_1811 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_7911_ _0102_ clknet_leaf_26_i_clk net156 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_223_3183 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_223_3194 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_195_609 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7025__C1 _3209_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4734__S _1246_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_222_289 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7842_ _0035_ clknet_leaf_67_i_clk core_0.fetch.out_buffer_data_instr\[19\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__6379__A1 _2244_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4641__A4 net182 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_203_470 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_203_492 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_77_158 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_350 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7773_ _1136_ _3846_ _0497_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__4929__A2 _1390_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4985_ _0781_ _0773_ core_0.dec_l_reg_sel\[0\] _1434_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_4
XANTENNA__5051__A1 net91 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_195_2857 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6724_ _2981_ _3021_ _3033_ _0261_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_3936_ _0564_ _0528_ _0566_ _0569_ _0570_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai211_4
XFILLER_0_129_772 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_135_208 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_545 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_190_314 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_18_247 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_865 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_128_271 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_144_731 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6655_ _2979_ core_0.ew_data\[13\] _2980_ net25 _2992_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_0_61_504 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5606_ _1643_ _1476_ _2004_ _2006_ _2007_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai31_4
XTAP_TAPCELL_ROW_30_871 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_119_1940 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_61_559 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_82_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6586_ _2935_ _2936_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_5_174 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_116_499 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_171_594 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8325_ _0501_ clknet_leaf_79_i_clk core_0.dec_rf_ie\[5\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5537_ _1961_ _1172_ _1962_ _1950_ _0145_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__5364__I _1811_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_131_458 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_100_801 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8256_ _0432_ clknet_leaf_32_i_clk core_0.execute.sreg_scratch.o_d\[6\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_41_294 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6303__A1 _1114_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_112_661 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_169_72 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5468_ _1898_ _1817_ _1902_ _1748_ _0136_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XANTENNA_input54_I i_req_data[24] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7207_ _1195_ core_0.execute.sreg_irq_pc.o_d\[2\] _3393_ _3394_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4419_ _0883_ _1022_ _1023_ _0963_ net169 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XFILLER_0_246_849 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8187_ _0363_ clknet_leaf_125_i_clk core_0.execute.alu_mul_div.mul_res\[13\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5399_ core_0.execute.alu_mul_div.div_cur\[5\] _1811_ _1843_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_7138_ _1915_ _1549_ _3344_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__7803__A1 core_0.decode.i_instr_l\[13\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7803__B2 core_0.decode.i_instr_l\[10\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_198_403 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7069_ _3273_ _3280_ _3281_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_2_541 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_69_615 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_output210_I net210 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5290__A1 core_0.dec_jump_cond_code\[4\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_241_587 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_213_278 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_83_1505 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_38_971 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_185_119 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_136 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_EDGE_ROW_226_Right_226 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__7031__A2 _1631_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_169 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_159_2421 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_204_34 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_77_670 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5042__A1 _0576_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5539__I _1963_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_194_653 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4443__I core_0.decode.i_instr_l\[0\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_383 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_534 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_49_394 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_139 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_204_78 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6790__A1 _2961_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_181_314 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_353 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_80_802 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_147_580 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_107_422 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_119_282 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_52_515 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xinput19 i_mc_core_int net19 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_64_397 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5345__A2 _1752_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_162_594 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_20_401 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_94_1645 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_32_283 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_818 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_102_171 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6845__A2 _3087_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_236_326 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_217_562 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_205_702 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_217_573 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_204_201 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4608__A1 _0726_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_232_521 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6038__C _1686_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5281__A1 _1430_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_181_18 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_clkbuf_leaf_18_i_clk_I clknet_4_8__leaf_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_220_749 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87_467 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_90_49 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_157_322 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_75_629 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_114_34 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4353__I _0965_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_74_128 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_103_1752 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_157_366 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4770_ core_0.fetch.prev_request_pc\[3\] _1285_ _0881_ net170 _1289_ vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_0_28_545 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6781__A1 _2940_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_172_303 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_185_697 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6989__B _3175_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_83_640 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_865 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_145_539 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_138_591 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_126_753 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_55_397 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6440_ _2812_ _2813_ _2819_ _2820_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_99_69 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_130_55 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_190_2787 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_141_734 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_190_2798 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_2_111 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_125_296 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_180_391 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6371_ _2663_ _2723_ _2753_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_51_581 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8110_ _0286_ clknet_leaf_102_i_clk core_0.execute.rf.reg_outputs\[3\]\[1\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_2
X_5322_ core_0.execute.alu_mul_div.div_cur\[1\] _1556_ _1557_ _1770_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_0_2_177 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_8041_ _0218_ clknet_leaf_55_i_clk core_0.ew_mem_access vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__6836__A2 _3086_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_139_42 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5253_ _1528_ _1529_ _1702_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_0_227_326 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_489 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_114_1881 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4698__I1 net66 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_225_3212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_4204_ _0723_ net58 _0822_ _0823_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_4
X_5184_ core_0.execute.rf.reg_outputs\[5\]\[4\] _1604_ _1605_ core_0.execute.rf.reg_outputs\[7\]\[4\]
+ _1606_ core_0.execute.rf.reg_outputs\[3\]\[4\] _1633_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_0_208_562 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4135_ _0731_ _0753_ _0754_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_2
XTAP_TAPCELL_ROW_143_2233 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7261__A2 _3398_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4066_ net212 net203 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_3
XANTENNA__5272__A1 _1123_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_78_412 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_211_727 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_78_423 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_204_790 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_176_620 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7825_ _0018_ clknet_leaf_60_i_clk core_0.fetch.out_buffer_data_instr\[2\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_35_930 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_148_333 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_59_670 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4263__I _0881_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_523 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_176_664 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_65_139 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_236_3341 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_7756_ core_0.dec_jump_cond_code\[4\] _3766_ _3832_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_136_517 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_163_303 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5575__A2 _0742_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4968_ _1419_ _1421_ _0117_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_58_191 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6772__A1 _2992_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_74_651 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6899__B _3124_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_62_802 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6707_ core_0.execute.rf.reg_outputs\[5\]\[1\] _3022_ _3016_ _3024_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3919_ core_0.execute.rf.reg_outputs\[2\]\[14\] _0554_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_163_347 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7687_ _1038_ _1102_ _3787_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_190_144 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4899_ _1231_ _1362_ _1363_ _1365_ _0104_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai31_1
X_6638_ _2979_ core_0.ew_mem_width _2980_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_4
XTAP_TAPCELL_ROW_154_2362 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_21_209 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_132_745 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_171_380 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6569_ _2925_ _0214_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_131_244 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8308_ _0484_ clknet_leaf_74_i_clk net193 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_4
XTAP_TAPCELL_ROW_7_600 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7523__B _3651_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_246_624 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8239_ _0415_ clknet_leaf_39_i_clk core_0.execute.sreg_irq_pc.o_d\[11\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__6827__A2 _3092_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_30_798 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_245_112 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4838__A1 _1280_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4689__I1 net60 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_165_2491 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_242_852 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7252__A2 core_0.execute.sreg_irq_pc.o_d\[7\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_199_745 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5978__B _2300_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4882__B _0881_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_97_765 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_215_66 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7004__A2 _3178_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_139_322 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_69_478 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_215_88 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_96_275 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_215_99 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_210_760 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_69_Right_69 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_37_320 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6763__A1 _2983_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5566__A2 _1957_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_865 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_127_539 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_42_1021 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_65_662 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_673 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_731 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_108_742 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_13_668 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_154_358 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_170_807 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_41_999 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_107_252 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5318__A2 _1765_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6515__A1 core_0.execute.alu_mul_div.div_cur\[15\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_122_211 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5869__A3 _1197_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_122_233 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_150_597 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_EDGE_ROW_78_Right_78 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_110_439 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_648 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6818__A2 _3087_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4829__A1 _1280_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_236_123 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_20_297 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_236_134 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_53_1150 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7779__B1 _3833_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7911__CLK clknet_leaf_26_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7243__A2 net83 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5254__A1 _1701_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_220_3153 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_125_22 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87_220 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5940_ _0799_ _2332_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_177_417 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_87_Right_87 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_125_66 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_618 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_125_77 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87_275 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_140_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5871_ _2263_ _2264_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA__5006__A1 _1452_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_238_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_87_286 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6054__I0 core_0.ew_data\[3\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7610_ net216 _3675_ _3727_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_32_900 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_87_297 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_4822_ _1317_ core_0.fetch.submitable _1318_ _0074_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__5557__A2 _1955_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_192_2816 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_157_174 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_8_737 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_44_802 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_146_859 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_90_418 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7541_ core_0.execute.sreg_irq_flags.o_d\[3\] _1398_ _1357_ _3667_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_4753_ _0845_ _1238_ _1277_ _0046_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_173_656 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_161_818 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_71_632 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_83_492 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5309__A2 _1756_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7472_ _0553_ _3546_ _3541_ _3623_ _3624_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_172_177 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4684_ net38 _1238_ _1239_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_126_583 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6423_ _2074_ _2801_ _2803_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_113_222 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_114_745 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_116_1910 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_31_529 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_231_3282 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_12_710 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_96_Right_96 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_24_592 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6354_ _2052_ _2735_ _2736_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_59_72 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_228_613 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_11_253 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5305_ _1505_ _1506_ _1753_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__6809__A2 _3065_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_227_101 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_264 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6285_ _2668_ _2602_ _2102_ _2669_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_8024_ _0201_ clknet_leaf_37_i_clk net128 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5236_ _1480_ _1602_ _1681_ _1684_ _1685_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_0_45_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4296__A2 net46 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5493__A1 core_0.execute.alu_mul_div.cbit\[0\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_242_104 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5167_ core_0.execute.rf.reg_outputs\[1\]\[7\] _1615_ _1434_ core_0.execute.rf.reg_outputs\[6\]\[7\]
+ _1616_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_242_137 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5798__B _2183_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4118_ _0734_ _0737_ _0738_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__7234__A2 _3418_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_16_Left_263 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_98_518 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5098_ core_0.execute.rf.reg_outputs\[1\]\[15\] _1484_ _1486_ core_0.execute.rf.reg_outputs\[5\]\[15\]
+ core_0.execute.rf.reg_outputs\[6\]\[15\] _1435_ _1547_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi222_2
XANTENNA__5245__A1 _1466_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input17_I i_disable vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_223_373 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_67_1319 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_211_524 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4049_ _0516_ _0523_ _0526_ core_0.execute.rf.reg_outputs\[2\]\[4\] _0674_ vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_1
XANTENNA__5796__A2 _2194_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_765 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_182_72 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_195_258 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_117 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_93_212 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_66_437 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7808_ _0789_ _1134_ _3869_ _1279_ _0509_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_176_461 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_66_459 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_109_517 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5548__A2 _1172_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_176_472 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_109_539 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_176_483 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_148_185 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7739_ net183 core_0.decode.i_imm_pass\[14\] _1063_ _3821_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_164_667 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4220__A2 _0836_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_46_172 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_481 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_46_183 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XPHY_EDGE_ROW_25_Left_272 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__7237__C _1736_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_10_627 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_10_638 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_117_583 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_367 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_61_142 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7170__A1 _3357_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_78_1448 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_104_244 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_91_1604 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output85_I net85 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_104_288 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_120_737 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_219_624 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_246_410 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_167_2520 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7934__CLK clknet_leaf_32_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7473__A2 _3542_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4287__A2 _0836_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5484__A1 _1915_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_218_189 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6584__S _2929_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_34_Left_281 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
Xclkbuf_4_3__f_i_clk clknet_3_1_0_i_clk clknet_4_3__leaf_i_clk vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__7700__C _1279_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_230_811 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5236__A1 _1480_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_89_1577 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_214_384 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_202_524 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_186_203 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6984__A1 core_0.execute.alu_mul_div.cbit\[1\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_18_727 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5787__A2 _2187_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_85_702 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_97_562 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_186_247 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_69_275 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_139_130 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_85_746 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_139_152 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6736__A1 _2994_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_210_590 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_100_1711 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_155_623 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4598__I0 core_0.ew_data\[5\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_26_802 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_43_Left_290 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_25_301 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6332__B _1117_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4211__A2 net59 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_111_i_clk clknet_4_4__leaf_i_clk clknet_leaf_111_i_clk vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_65_481 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_25_323 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_632 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_492 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_142_317 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_25_356 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_170_637 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_80_473 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_337 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_126_i_clk clknet_4_1__leaf_i_clk clknet_leaf_126_i_clk vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_96_26 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_96_37 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_562 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_96_48 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_209_3015 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_209_3026 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_0_478 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_111_1840 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7464__A2 _3616_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6070_ _2111_ _1601_ _1721_ _2113_ _2110_ _2459_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai32_4
XFILLER_0_29_64 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input9_I i_core_int_sreg[2] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_225_627 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_188_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_237_487 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5021_ _1462_ _1469_ _1451_ _1470_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_4
XTAP_TAPCELL_ROW_127_2036 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7216__A2 _3398_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_206_863 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5411__B _1841_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_221_844 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6972_ core_0.execute.alu_mul_div.cbit\[3\] _3180_ _3185_ _3191_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_1
XANTENNA__6975__A1 _2386_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5778__A2 net214 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_178_737 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_221_855 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4825__I1 core_0.decode.i_instr_l\[10\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_220_343 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_220_354 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5923_ _1554_ _1631_ _2314_ _2315_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_76_713 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_75_212 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_177_269 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_220_387 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_48_437 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4742__S _1246_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_192_217 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5854_ _2246_ net192 _1199_ _1200_ _2247_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_0_118_314 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_61_62 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_122_1980 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_29_662 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_63_407 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_267 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_158_494 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4805_ _1039_ _1307_ _1309_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_233_3311 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_5785_ core_0.execute.rf.reg_outputs\[3\]\[0\] _1606_ _1615_ core_0.execute.rf.reg_outputs\[1\]\[0\]
+ _2186_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_134_807 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_146_667 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_28_172 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7524_ _0604_ _3641_ _3657_ _0437_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_138_2165 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_4736_ core_0.fetch.out_buffer_data_instr\[22\] net52 _1246_ _1269_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_90_259 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_440 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5950__A2 core_0.execute.sreg_irq_pc.o_d\[1\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_160_125 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_126_391 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_160_136 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7455_ core_0.execute.sreg_irq_pc.o_d\[12\] _3542_ _3609_ _3610_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_151_2321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_43_175 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4667_ _1222_ _1223_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XANTENNA__7152__A1 _1375_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_160_158 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6406_ core_0.execute.sreg_priv_control.o_d\[12\] _1386_ _2577_ core_0.execute.sreg_irq_pc.o_d\[12\]
+ _2787_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_101_203 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_114_586 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7386_ _1980_ _3552_ _0404_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_4598_ core_0.ew_data\[5\] core_0.ew_data\[13\] _1150_ _1164_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_101_236 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6337_ _2718_ _2719_ _2720_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_clkbuf_4_3__f_i_clk_I clknet_3_1_0_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7455__A2 _3542_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6268_ _2623_ _2625_ _2652_ _2356_ _2653_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
Xclkbuf_leaf_90_i_clk clknet_4_6__leaf_i_clk clknet_leaf_90_i_clk vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_TAPCELL_ROW_73_1389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_177_94 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_244_3440 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4269__A2 _0823_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5466__A1 _1233_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_8007_ _0184_ clknet_leaf_54_i_clk core_0.ew_data\[6\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_243_424 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5219_ _0771_ _0768_ core_0.execute.rf.reg_outputs\[7\]\[2\] _1668_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_2
X_6199_ _1379_ core_0.execute.sreg_irq_pc.o_d\[7\] _2584_ _2585_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_243_457 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_230_107 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_224_671 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5321__B core_0.execute.alu_mul_div.div_cur\[0\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_162_2461 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_169_726 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_211_321 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_196_523 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6966__A1 _1223_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_551 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_79_562 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_169_759 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_168_247 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_724 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_94_510 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_211_376 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6931__I core_0.execute.alu_mul_div.mul_res\[0\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6718__A1 core_0.execute.rf.reg_outputs\[5\]\[6\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_137_623 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6194__A2 _1386_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_212_34 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7391__A1 _0709_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_35_632 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_492 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_23_785 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_124_317 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_191_272 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5941__A2 _2332_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_151_114 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_191_294 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3952__A1 _0539_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_304 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_leaf_43_i_clk clknet_4_9__leaf_i_clk clknet_leaf_43_i_clk vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__7143__A1 core_0.execute.alu_mul_div.mul_res\[15\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_173_2590 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_50_646 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_132_361 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_leaf_58_i_clk clknet_4_14__leaf_i_clk clknet_leaf_58_i_clk vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_120_589 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_246_240 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_207_605 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8112__CLK clknet_leaf_94_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_234_457 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_237_86 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_215_671 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6406__B1 _2577_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4680__A2 _0727_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6957__A1 _3175_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_159_214 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_159_225 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_202_343 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_230_663 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_187_556 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_202_365 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_85_510 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_57_212 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_79 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_202_387 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_176_2619 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_48_1093 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_85_576 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_116_807 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_122_34 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6185__A2 _2571_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_122_45 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_128_667 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7382__A1 _3547_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4196__A1 _0724_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5570_ _1283_ _1980_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_25_131 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_5_537 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_25_142 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_170_445 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3943__A1 core_0.dec_r_reg_sel\[2\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_31_98 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_559 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4521_ _1109_ _1062_ _1110_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_108_391 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_215_3096 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7134__A1 _3189_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_101 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_103_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_130_309 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7240_ net83 _3422_ _3423_ _1735_ _3424_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_40_145 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7685__A2 _1095_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4452_ core_0.decode.i_instr_l\[4\] _1047_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__inv_1
XANTENNA__5696__A1 _1124_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4499__A2 _1039_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_189 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7171_ _1369_ _1227_ _1364_ _3369_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_2
X_4383_ _0844_ _0947_ _0970_ _0995_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XTAP_TAPCELL_ROW_187_2759 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6122_ _2506_ _2508_ _2509_ _2510_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA__7437__A2 _3543_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6053_ _2346_ _2441_ _2442_ _2443_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_56_51 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_56_62 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_73 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5004_ core_0.decode.oc_alu_mode\[9\] core_0.decode.oc_alu_mode\[11\] core_0.decode.oc_alu_mode\[3\]
+ core_0.decode.oc_alu_mode\[2\] _1453_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_0_212_107 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_206_682 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6948__A1 _1225_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_178_523 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7070__B1 _3173_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_702 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7070__C2 _1585_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6955_ _3175_ _3172_ _3176_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA_clkbuf_leaf_66_i_clk_I clknet_4_15__leaf_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_48_201 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4423__A2 _0947_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5620__A1 _2018_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_48_212 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6751__I _3041_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5906_ _2102_ _2297_ _2298_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or2_4
XFILLER_0_48_234 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_49_757 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_138_Right_138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_198_2888 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6886_ core_0.execute.rf.reg_outputs\[1\]\[14\] _3106_ _3124_ _3126_ vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_159_792 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_91_502 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_119_645 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_204 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_146_431 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5837_ _2227_ _2230_ _2231_ _2232_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_29_470 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7373__A1 _1209_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_29_492 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_17_632 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_119_689 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4187__A1 core_0.ew_mem_access vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_63_248 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_91_557 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5923__A2 _1631_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5768_ _2051_ _2058_ _2169_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_146_497 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_44_451 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7507_ _1403_ _3640_ _3647_ _0430_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_32_613 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_20_755 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_4719_ net43 _1253_ _1260_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__7125__A1 _1994_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6700__B _3016_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_133_158 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_16_186 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5699_ core_0.decode.oc_alu_mode\[12\] _1553_ _2100_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_75_1407 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_7438_ _3581_ _3595_ _0413_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_31_134 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_75_1418 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5687__A1 _1124_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8135__CLK clknet_leaf_104_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_130_865 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7369_ _3535_ _3536_ _3537_ _0402_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_228_251 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7531__B _3651_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_216_424 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8285__CLK clknet_leaf_29_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6100__A2 _1385_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_216_457 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_99_602 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4111__A1 core_0.execute.prev_sys vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_243_265 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_207_34 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_98_101 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6939__A1 _1227_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_98_145 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_86_1547 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_28_844 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_196_331 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_211_151 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4890__B _1284_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_212 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5611__A1 _2010_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_196_375 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_105_Right_105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__7739__I0 net183 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_278 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_418 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_535 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_137_464 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_192_570 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4178__A1 core_0.ew_submit vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4178__B2 _0796_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_164_272 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_35_451 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5914__A2 _1568_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_180_732 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3925__A1 _0539_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7116__A1 _1364_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6610__B _1978_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_152_489 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_97_1676 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_50_454 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_22_167 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_31_690 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4350__A1 core_0.fetch.prev_request_pc\[14\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7419__A2 _3543_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_219_251 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7441__B _3553_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_207_457 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_93_38 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_124_2006 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_117_45 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4356__I net76 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_117_67 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_222_449 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_188_832 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_117_89 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_188_865 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4405__A2 _0966_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_543 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6740_ _3041_ _3042_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_86_863 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3952_ _0539_ _0542_ _0544_ core_0.execute.rf.reg_outputs\[1\]\[12\] _0585_ vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_4
XTAP_TAPCELL_ROW_106_1783 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_217_3114 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_9_139 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_133_66 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_220_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6671_ core_0.execute.rf.reg_outputs\[6\]\[2\] _3000_ _2984_ _3003_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3883_ _0518_ core_0.dec_r_reg_sel\[1\] _0519_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_0_128_464 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4169__A1 core_0.ew_reg_ie\[5\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5622_ _1715_ _1934_ _2023_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_143_412 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_771 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_135_2135 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8158__CLK clknet_leaf_88_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_143_445 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_345 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5553_ core_0.execute.mem_stage_pc\[10\] _1955_ _1964_ _1972_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_143_489 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4504_ _1046_ _1068_ _1094_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_8272_ _0448_ clknet_leaf_26_i_clk core_0.execute.pc_high_out\[1\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_41_454 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_170_286 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5484_ _1915_ _1491_ _1916_ _1917_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__5669__A1 _1752_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7223_ _3397_ _3409_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_13_178 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_112_865 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4435_ core_0.decode.i_flush _1030_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_1_562 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6330__A2 _2711_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_228_3243 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_7154_ _1727_ _3356_ _3357_ _0367_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_111_386 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4366_ _0965_ _0978_ _0980_ _0981_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_0_10_863 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_50 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_228_3254 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_67_72 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6105_ _1378_ core_0.execute.sreg_irq_pc.o_d\[5\] _2493_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_70_1348 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_7085_ _1909_ _1568_ _3294_ _3295_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_241_3410 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_207_Right_207 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
X_4297_ core_0.fetch.prev_request_pc\[1\] _0914_ _0915_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_225_232 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6094__A1 _2360_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6036_ _1121_ _2009_ _2146_ _1107_ _1059_ _2426_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_0_225_265 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_198_607 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_146_2264 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5841__A1 _2232_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_241_747 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_83_93 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7987_ _0164_ clknet_leaf_30_i_clk core_0.execute.prev_pc_high\[6\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_221_460 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7594__A1 _3675_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_194_802 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_95_126 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_194_813 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_25_814 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_138_206 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_554 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6938_ _1231_ _1831_ _1601_ _1926_ _1225_ _3159_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_0_178_397 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_92_800 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_239_3383 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_64_524 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_190_94 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6869_ core_0.execute.rf.reg_outputs\[1\]\[6\] _3114_ _3112_ _3117_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_76_384 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7346__A1 core_0.execute.alu_flag_reg.o_d\[2\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_147_762 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_81_1488 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_92_855 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_106_103 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_626 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_174_581 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_107_648 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_462 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_125 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_157_2393 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output190_I net190 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_161_242 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_162_765 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_44_270 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4580__A1 core_0.ew_data\[4\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_161_286 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_32_465 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_121_139 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_20_627 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6321__A2 _2642_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_236_508 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_130_695 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_217_722 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_8_Left_255 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_244_541 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6085__A1 _1690_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6085__B2 _1929_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7821__A2 _3767_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_5_572 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5832__A1 _2226_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_169_320 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_197_640 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87_627 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_231_279 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7585__A1 core_0.execute.pc_high_buff_out\[4\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_240_791 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4399__A1 _1004_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_184_312 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_200_644 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_863 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_157_537 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_28_705 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5060__A2 net179 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_184_334 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_727 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_822 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_45_1052 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_94_170 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_55_535 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_137_250 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_27_248 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_99_1705 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_12_34 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_125_412 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_82_354 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_103_58 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_70_527 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5899__A1 _1059_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_153_754 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7436__B _3545_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5899__B2 _1107_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_82_387 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_793 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_179_18 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_35_292 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_212_3055 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_50_240 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput107 net107 o_icache_flush vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA_clkbuf_leaf_14_i_clk_I clknet_4_8__leaf_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput118 net118 o_mem_addr[11] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_11_627 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput129 net129 o_mem_addr[7] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_23_487 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_191 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_121_640 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_239_346 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_121_684 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_239_368 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4220_ _0835_ _0836_ _0837_ _0838_ _0839_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor4_4
XANTENNA__4174__I1 core_0.ew_reg_ie\[1\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_130_2076 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_184_2718 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_208_711 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_56_1181 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4874__A2 _1341_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4151_ core_0.dec_l_reg_sel\[2\] _0770_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_235_530 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_207_221 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6076__A1 _1999_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_207_243 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5403__C _1822_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4082_ _0533_ _0524_ _0527_ core_0.execute.rf.reg_outputs\[6\]\[1\] _0704_ vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_4
XANTENNA__4087__B1 _0703_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_170_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_108_1812 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_222_224 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7910_ _0101_ clknet_leaf_52_i_clk core_0.fetch.pc_reset_override vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_223_769 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_223_3184 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_7841_ _0034_ clknet_leaf_67_i_clk core_0.fetch.out_buffer_data_instr\[18\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__7025__C2 _1613_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_188_662 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7576__A1 _3682_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5036__C1 net218 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_176_802 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_52 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7772_ core_0.dec_rf_ie\[1\] _3766_ _3833_ _3845_ _3846_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_4984_ core_0.execute.alu_mul_div.i_mul _1433_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_144_98 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_92_107 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_195_2847 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5051__A2 _1492_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_148_559 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_195_2858 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6723_ core_0.execute.rf.reg_outputs\[5\]\[8\] _3027_ _3031_ _3033_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_46_524 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3935_ _0568_ core_0.execute.rf.reg_outputs\[3\]\[13\] _0549_ _0569_ vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_0_46_535 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_855 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6654_ _2941_ _2990_ _2991_ _0233_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_160_53 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_34_719 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_190_348 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_116_434 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_160_75 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6000__A1 _2360_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5605_ _1558_ _2005_ _2006_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__7346__B _3516_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_73_398 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_142 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6585_ core_0.ew_reg_ie\[7\] _2934_ _2935_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_2
XTAP_TAPCELL_ROW_119_1941 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_171_562 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_30_872 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_6_687 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8324_ _0500_ clknet_leaf_86_i_clk core_0.dec_rf_ie\[4\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_131_426 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5536_ net81 _1953_ _1962_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_41_240 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_103_128 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_75_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_8255_ _0431_ clknet_leaf_25_i_clk core_0.execute.sreg_scratch.o_d\[5\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5467_ core_0.execute.alu_mul_div.div_cur\[13\] _1838_ _1816_ _1901_ _1902_ vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XANTENNA__6303__A2 _2686_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7500__A1 _0709_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_112_684 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7206_ _3386_ _1195_ _3393_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_4418_ net80 _0883_ _1023_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_246_828 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8186_ _0362_ clknet_leaf_125_i_clk core_0.execute.alu_mul_div.mul_res\[12\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5398_ _1840_ _1842_ _0126_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA_input47_I i_req_data[18] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7137_ core_0.execute.alu_mul_div.mul_res\[14\] _1941_ _3343_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__and2_1
X_4349_ _0965_ _0966_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_226_563 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7068_ core_0.execute.alu_mul_div.mul_res\[9\] _3279_ _3280_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__7803__A2 _3788_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5814__A1 _2205_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6019_ _2306_ _2303_ _1559_ _2409_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_2_531 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_241_544 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4173__S0 _0769_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_2_542 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_213_257 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_68_104 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_69_627 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_179_640 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_201_419 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_190_Right_190 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__7567__A1 core_0.execute.pc_high_out\[1\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_83_1506 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8323__CLK clknet_leaf_83_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_222_780 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_38_972 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_167_813 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_output203_I net203 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_178_161 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_49_340 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_159_2422 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_193_120 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5042__A2 _1483_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_139_559 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_204_57 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_193_142 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_524 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7319__A1 net78 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_64_321 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6790__A2 _3064_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_37_557 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_401 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_119_261 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_135_710 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_9_481 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_9_492 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_52_527 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_64_387 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_91_173 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_134_242 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_220_34 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_91_184 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_135_776 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_60_560 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_150_757 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_32_262 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_94_1635 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_60_582 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_94_1646 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4305__A1 core_0.fetch.prev_request_pc\[7\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_457 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_103_695 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_102_183 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_236_338 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_229_390 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6058__A1 net186 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_205_725 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_244_382 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5805__A1 _2183_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4608__A2 _0727_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_245_42 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5281__A2 net194 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7558__A1 _3637_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_87_446 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_169_150 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_197_470 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_197_492 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6230__A1 _2576_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_74_107 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_103_1753 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_184_142 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_524 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_200_485 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_23_66 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_55_332 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_56_855 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6781__A2 _3064_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_28_557 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_16_699 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4792__A1 _1290_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_365 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_126_732 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_218 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_82_162 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_99_59 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_858 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_141_702 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_153_584 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_190_2788 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_153_595 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_180_370 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6370_ _2749_ _2750_ _2751_ _2752_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_4
XFILLER_0_130_78 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_774 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_58_1210 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_2_123 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_140_234 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_11_402 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5321_ _1551_ _1552_ core_0.execute.alu_mul_div.div_cur\[0\] _1769_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XANTENNA__6297__A1 _2311_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_8040_ _0217_ clknet_leaf_81_i_clk core_0.ew_reg_ie\[7\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__dffq_2
X_5252_ _1526_ _1527_ _1701_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_0_11_479 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_121_492 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_114_1882 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_139_54 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4847__A2 _1336_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4203_ _0723_ _0821_ _0822_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_225_3213 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_5183_ net98 _1446_ _1632_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__6049__A1 core_0.execute.alu_mul_div.div_cur\[3\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7246__B1 _3399_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4134_ _0738_ _0741_ _0752_ _0753_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_0_235_360 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_235_382 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_223_533 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_143_2223 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_4065_ _0680_ _0683_ _0688_ _0521_ net97 _0689_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai32_4
XTAP_TAPCELL_ROW_143_2234 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_211_706 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5272__A2 _1451_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_64_73 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_78_435 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7824_ _0017_ clknet_leaf_61_i_clk core_0.fetch.out_buffer_data_instr\[1\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_35_931 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_93_416 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6221__A1 _2281_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5024__A2 core_0.execute.alu_flag_reg.o_d\[1\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_148_345 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4967_ core_0.execute.sreg_priv_control.o_d\[11\] _1393_ _1420_ _1391_ _1421_ vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_58_170 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7755_ _3769_ _1072_ _1032_ _1084_ _3831_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai211_2
XTAP_TAPCELL_ROW_236_3342 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6772__A2 _3043_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_557 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_129_570 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_164_849 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4783__A1 core_0.fetch.prev_request_pc\[9\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3918_ _0553_ net200 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_6706_ _2940_ _3021_ _3023_ _0253_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__4783__B2 net176 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_190_123 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7686_ _3777_ _3783_ _3784_ _3785_ _3786_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_4
X_4898_ _1364_ _1221_ _1365_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_73_162 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_387 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_34_527 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6637_ _2929_ _2979_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_8
XFILLER_0_190_156 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_6_451 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_61_346 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_154_2363 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_116_275 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_61_368 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_426 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_131_212 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_EDGE_ROW_89_Left_336 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
X_6568_ core_0.dec_rf_ie\[4\] core_0.ew_reg_ie\[4\] _2201_ _2925_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_131_256 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_8307_ _0483_ clknet_leaf_76_i_clk net192 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_4
X_5519_ core_0.execute.sreg_data_page _0807_ _1949_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_6499_ _1109_ _1989_ _2876_ _1987_ _2741_ _2877_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_0_131_278 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_219_828 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8238_ _0414_ clknet_leaf_40_i_clk core_0.execute.sreg_irq_pc.o_d\[10\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_7_601 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_100_621 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_218_305 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4299__B1 _0914_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4299__C2 _0860_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4838__A2 net42 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8338__D _0514_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_218_349 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_8169_ _0345_ clknet_leaf_85_i_clk net91 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_4
XFILLER_0_245_168 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7788__A1 _1136_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_165_2492 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_98_Left_345 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_241_352 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_69_402 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6460__A1 _2078_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5263__A2 _1524_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_201_205 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_214_599 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_201_216 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_198_267 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_186_418 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_96_254 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_167_632 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_179_492 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6212__A1 _2287_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_56_107 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5015__A2 _0661_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_210_772 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_127_507 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_210_794 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_855 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6763__A2 _3042_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_42_1011 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_182_624 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_42_1022 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4774__A1 _1290_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_107_220 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_13_669 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_52_313 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_398 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_538 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_231_88 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_858 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_123_702 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_135_562 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6515__A2 _1117_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7712__A1 _1382_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_107_264 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_108_798 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_135_573 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_357 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_275 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_69_18 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_100_26 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_100_37 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7714__B _3808_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_766 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_110_429 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6110__S _1625_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_265 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_236_102 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_53_1151 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_233_842 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_189_223 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_205_566 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6451__A1 _1380_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5254__A2 _1702_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_88_722 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_232_374 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_220_3154 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_149_109 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_48_608 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5870_ _1196_ _1201_ _2262_ _2263_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_0_158_643 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_427 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_201_772 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_157_142 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_4821_ _0938_ _1170_ _1318_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_32_901 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_28_310 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_133_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6754__A2 _3049_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_145_304 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_192_2817 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_28_343 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_64_1280 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_7540_ _3663_ _3666_ _0444_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_4752_ net61 _1241_ _1277_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4765__A1 _1284_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_145_337 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_83_460 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_611 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6512__C _0799_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_16_527 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_141_66 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_43_324 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_398 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_154_860 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7471_ _3547_ net78 _3540_ _3622_ _3623_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_172_167 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4683_ _1236_ _1238_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_55_195 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7703__A1 _3773_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6422_ _2074_ _2801_ _2802_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_113_212 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_116_1900 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_43_379 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_699 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_231_3283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_24_582 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_3_454 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7624__B _1216_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5190__A1 _1625_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6353_ _2058_ _2695_ _2056_ _2735_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_3_498 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5304_ _1510_ _1511_ _1752_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_4
X_6284_ _2120_ _2094_ _1819_ _2668_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_59_84 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_59_95 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8023_ _0200_ clknet_leaf_36_i_clk net127 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__4539__I _1123_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5235_ _1682_ _1683_ _1684_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or2_2
XANTENNA__6690__A1 _2986_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_243_628 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5166_ _1608_ _1615_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_38_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_236_691 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_72 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_166_85 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4117_ core_0.execute.prev_pc_high\[2\] _0735_ _0736_ core_0.execute.prev_pc_high\[1\]
+ _0737_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_224_864 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5097_ core_0.execute.rf.reg_outputs\[7\]\[15\] net232 _1443_ core_0.execute.rf.reg_outputs\[3\]\[15\]
+ _1546_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_223_352 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4048__A3 _0518_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6442__A1 _2281_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5245__A2 net188 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4048_ _0516_ _0540_ _0518_ core_0.execute.rf.reg_outputs\[1\]\[4\] _0673_ vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_1
XANTENNA__7886__CLK clknet_leaf_81_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_66_405 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_79_788 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_149_632 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_182_84 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_107 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_94_747 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7807_ core_0.decode.i_instr_l\[15\] _3788_ _3866_ core_0.decode.i_instr_l\[12\]
+ _1132_ _3869_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_0_176_451 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6745__A2 _3043_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_94_769 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5999_ _2388_ _2389_ _2390_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_0_149_698 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_419 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_136_337 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7738_ _3820_ _0488_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_163_123 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_191_454 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_302 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4220__A3 _0837_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_35_836 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_62_633 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_858 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_105_702 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_562 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_10_628 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_7669_ _0514_ _1084_ _1072_ _3772_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_62_655 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_144_370 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_154 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_132_521 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_34_379 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_839 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_62_699 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_78_1449 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_132_543 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_160_863 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5181__A1 net99 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_91_1605 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_120_749 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_output78_I net78 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_30_585 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_246_422 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_167_2521 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_100_451 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_246_444 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6681__A1 core_0.execute.rf.reg_outputs\[6\]\[6\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5484__A2 _1491_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_227_680 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_233_138 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_215_842 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_89_508 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_215_864 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_214_330 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6433__A1 _2090_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4039__A3 _0518_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_89_1578 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_18_728 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_159_418 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_241_182 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_230_845 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_69_232 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4995__A1 _0770_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_85_714 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_416 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_84_213 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_298 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_449 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_178_2650 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_195_782 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6736__A2 _3022_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_84_257 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_100_1712 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_154_101 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_242_87 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4598__I1 core_0.ew_data\[13\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_154_123 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5944__B1 _2257_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_53_611 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_182_454 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_52_121 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_218 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_132 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_142_329 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_452 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_154_189 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_34 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_111_58 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_111_69 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_80_496 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5172__A1 _1553_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_390 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_150_384 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_21_574 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_209_3016 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_111_1841 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_209_146 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6672__A1 _2951_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5020_ _1464_ _1465_ _1467_ _1468_ _1469_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XTAP_TAPCELL_ROW_127_2037 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_119_Right_119 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_205_352 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_221_812 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5227__A2 net219 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6424__A1 _1457_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_232_171 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_220_311 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6971_ core_0.execute.alu_mul_div.cbit\[3\] _3185_ _3180_ _3190_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_177_204 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_88_541 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_204_2960 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_232_193 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_220_333 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5922_ _1553_ _2019_ _2314_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_88_574 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_88_585 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_220_377 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_48_427 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5853_ net187 _2246_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__inv_1
XANTENNA__6727__A2 _3027_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_145_101 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4738__A1 net53 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_8_524 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_91_717 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_118_326 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_122_1981 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_4804_ _0816_ _1306_ _1308_ _0066_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_233_3312 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_63_419 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_75_279 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5784_ _1442_ _2185_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_28_162 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_17_836 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4735_ _1268_ _0037_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7523_ core_0.execute.sreg_scratch.o_d\[11\] _3646_ _3651_ _3657_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_138_2166 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_17_858 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_133_318 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_161_627 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_160_104 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_133_329 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7454_ _0592_ _3546_ _3545_ _3608_ _3609_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_4666_ core_0.execute.alu_mul_div.cbit\[3\] _1222_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XTAP_TAPCELL_ROW_151_2322 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_32_839 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_142_863 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6405_ _2785_ _2759_ _2786_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_43_187 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5163__A1 net100 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_102_716 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_31_349 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7385_ core_0.execute.sreg_irq_pc.o_d\[0\] _3543_ _3551_ _3552_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4597_ _1163_ net142 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_12_541 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_141_384 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_clkbuf_leaf_62_i_clk_I clknet_4_14__leaf_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6336_ core_0.execute.sreg_scratch.o_d\[10\] _2579_ _2534_ net2 _2719_ vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__7073__C _1372_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_177_51 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6267_ _2650_ _2651_ _2652_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_4
XTAP_TAPCELL_ROW_244_3441 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_243_403 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_216_617 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6663__A1 _2941_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_8006_ _0183_ clknet_leaf_54_i_clk core_0.ew_data\[5\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_2
X_5218_ core_0.execute.rf.reg_outputs\[3\]\[2\] _1667_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_215_105 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6198_ _1378_ _2583_ _2584_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_149_2295 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_5149_ _1467_ _1196_ _1598_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_212_801 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6415__A1 core_0.ew_data\[12\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_162_2451 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_193_72 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_162_2462 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_79_530 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_169_738 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output116_I net116 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8064__CLK clknet_leaf_94_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4977__A1 _1419_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_596 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7529__B _3651_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_438 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6718__A2 _3027_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6433__B _2626_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_67_769 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_183_229 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_82_728 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_780 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7391__A2 _3544_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_75_791 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_23_786 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_117_381 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_133_830 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_151_126 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_688 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3952__A2 _0542_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_165 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_173_2591 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_62_485 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_62_496 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_576 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_160_671 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5563__I net78 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_120_524 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_132_384 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_219_422 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_207_617 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6654__A1 _2941_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_246_274 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_219_488 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_50_1110 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6406__A1 core_0.execute.sreg_priv_control.o_d\[12\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6327__C _2626_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_89_327 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_203_834 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_199_362 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_214_171 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_202_311 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6957__A2 _1689_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4968__A1 _1419_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_15_34 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_159_237 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_187_568 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_85_522 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6709__A2 _3022_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_769 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_48_1083 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_48_1094 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_73_706 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_85_566 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_408 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_128_679 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_61_1250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_182_251 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_38_493 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_170_413 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_441 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_549 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4520_ core_0.decode.oc_alu_mode\[9\] _1109_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_108_381 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3943__A2 core_0.dec_r_reg_sel\[1\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_81_772 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_14_839 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_142_148 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_170_457 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_215_3097 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_26_699 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_53_485 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_53_496 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_124_863 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_338 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7174__B core_0.execute.alu_mul_div.div_res\[7\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5145__A1 _1482_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4451_ core_0.decode.i_instr_l\[3\] _1045_ _1046_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_0_151_682 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_123_384 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5696__A2 _2019_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4499__A3 _1069_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6893__A1 net88 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7170_ _3357_ _3368_ _0372_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_4382_ _0959_ _0993_ _0994_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_1_766 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_111_568 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6121_ _2506_ _2508_ _1458_ _2509_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_238_786 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6645__A1 _2936_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6052_ core_0.dec_mem_access net203 _2442_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_EDGE_ROW_7_Right_7 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
X_5003_ _1123_ core_0.decode.oc_alu_mode\[13\] _1452_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_4
XANTENNA__4817__I core_0.decode.i_instr_l\[7\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4120__A2 _0739_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_221_642 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7070__A1 core_0.execute.alu_mul_div.mul_res\[9\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4959__A1 _1414_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6954_ _0803_ _3175_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_88_360 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_166_719 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5905_ _1721_ _2108_ _1625_ _2297_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__7349__B _3495_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_220_185 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_198_2889 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_76_544 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6885_ _2992_ _3108_ _3125_ _0330_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_64_717 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5836_ _0649_ _1444_ _1607_ _2231_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_4
XFILLER_0_17_600 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_173_240 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7373__A2 _2577_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_134_605 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4187__A2 core_0.ew_submit vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5384__A1 core_0.execute.alu_mul_div.div_cur\[3\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_17_644 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5767_ _2161_ _2162_ _2167_ _2168_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_134_627 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_387 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5584__S _1985_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_118_189 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7506_ core_0.execute.sreg_scratch.o_d\[4\] _3646_ _3516_ _3647_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_20_756 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_17_688 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4718_ core_0.fetch.out_buffer_data_instr\[14\] _1259_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_5698_ _2097_ _2098_ _1554_ _2099_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__7125__A2 _3209_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_130_800 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7437_ core_0.execute.sreg_irq_pc.o_d\[9\] _3543_ _3594_ _3595_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_75_1408 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_102_502 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6333__B1 _2713_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4649_ _1206_ _1208_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_31_146 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_102_524 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_188_72 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_130_855 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_141_192 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7368_ core_0.execute.alu_flag_reg.o_d\[4\] _3510_ _3516_ _3537_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XPHY_EDGE_ROW_203_Left_450 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_40_691 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_12_382 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_228_230 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6319_ _1109_ _2057_ _2701_ _2702_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_7299_ _1742_ _3467_ _3475_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6636__A1 _2936_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_110_i_clk clknet_4_5__leaf_i_clk clknet_leaf_110_i_clk vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_231_406 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_99_636 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4662__A3 _0810_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6939__A2 _1683_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_86_1548 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_28_845 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_67_500 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_212_686 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_211_163 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_125_i_clk clknet_4_1__leaf_i_clk clknet_leaf_125_i_clk vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__7259__B net86 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_95_842 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_39_246 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_211_196 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7739__I1 core_0.decode.i_imm_pass\[14\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_149_270 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_223_67 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_109_112 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_149_292 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7364__A2 _2434_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5375__A1 _1375_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_35_430 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_750 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_124_126 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_63_772 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_35_474 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_152_457 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_62_271 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_863 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5127__A1 net89 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_180_799 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_22_135 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_97_1677 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_120_310 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_132_170 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6875__A1 core_0.execute.rf.reg_outputs\[1\]\[9\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_120_354 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_120_387 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_120_398 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6627__A1 _2929_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4637__I net186 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_234_288 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5850__A2 core_0.dec_sreg_jal_over vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7052__A1 _3261_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_10_i_clk_I clknet_4_3__leaf_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_203_664 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_230_461 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_203_675 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_201_2930 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_187_365 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_202_174 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3951_ _0581_ _0528_ _0582_ _0583_ _0584_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai211_4
XFILLER_0_187_387 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_58_555 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_106_1784 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_46_706 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_9_129 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_352 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_217_3115 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_168_590 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6670_ _2946_ _2999_ _3002_ _0238_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_3882_ core_0.dec_r_reg_sel\[0\] _0518_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_42_76 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7355__A2 _2777_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_128_454 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_155_240 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5621_ _1761_ _1613_ _2022_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_2
XANTENNA__4169__A2 _0779_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_115_104 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_213_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_143_424 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_155_284 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5552_ _0991_ _1956_ _1971_ _0151_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_5_335 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_115_137 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_135_2136 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_143_457 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_171_766 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_5_357 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_115_159 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_170_243 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4503_ _1084_ _1092_ _1093_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5118__A1 _1561_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5417__B _1822_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_130_107 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8271_ _0447_ clknet_leaf_22_i_clk core_0.execute.pc_high_out\[0\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_41_444 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5483_ _1909_ net214 _1916_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_130_129 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6866__A1 _2961_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5669__A2 _1568_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4434_ _0742_ net115 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_2
X_7222_ _1742_ _3400_ _3408_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_112_855 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_41_488 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7632__B _1216_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7153_ _1747_ _3357_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
X_4365_ _0946_ _0955_ _0979_ _0980_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_1
XTAP_TAPCELL_ROW_228_3244 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6104_ net83 _2268_ _2491_ _2245_ _2492_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__6618__A1 _2936_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_171_Right_171 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
X_7084_ _1909_ _1576_ _3294_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_67_84 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7351__C _3510_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4296_ _0824_ net46 _0913_ _0914_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_4
XTAP_TAPCELL_ROW_70_1349 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_241_3400 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_226_756 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6094__A2 _2482_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6035_ _1765_ _1665_ _2425_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_2
XTAP_TAPCELL_ROW_146_2265 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_20_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XPHY_EDGE_ROW_61_Left_308 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
Xrebuffer10 _0784_ net232 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlya_2
XFILLER_0_241_759 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_240_236 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_leaf_42_i_clk clknet_4_9__leaf_i_clk clknet_leaf_42_i_clk vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_240_247 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7043__A1 _2587_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_83_72 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_83_83 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_95_105 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7986_ _0163_ clknet_leaf_28_i_clk core_0.execute.prev_pc_high\[5\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_89_680 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_25_815 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_95_138 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_77_842 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6937_ _3157_ _3158_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_166_527 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_178_387 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_193_324 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_49_566 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_193_335 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_239_3384 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_57_i_clk clknet_4_14__leaf_i_clk clknet_leaf_57_i_clk vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_6868_ _2967_ _3107_ _3116_ _0322_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__7346__A2 _3510_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8102__CLK clknet_leaf_107_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_81_1489 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_119_476 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_162_711 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_685 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5819_ net134 _2209_ _2217_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6711__B _3016_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6799_ _2981_ _3064_ _3076_ _0293_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_106_115 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_174_593 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_146_295 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_45_772 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_157_2394 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_70_Left_317 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_134_457 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_159 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_17_496 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_output183_I net183 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_170_2550 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4580__A2 net157 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_102_387 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6609__A1 _2930_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_217_734 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_218_34 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_217_745 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_218_45 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7282__A1 _2752_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6085__A2 _2013_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4096__A1 _0568_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_5_573 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_99_422 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_232_737 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_244_597 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_232_748 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_181_2690 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_231_258 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_231_269 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5045__B1 _1443_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7585__A2 _3682_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_197_674 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_157_505 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4399__A2 _0966_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_196_162 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5596__A1 _1765_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_185_858 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_67_352 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4192__I _0810_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_200_667 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_196_195 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_138_741 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_45_1053 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_55_525 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_138_752 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7337__A2 _3495_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_184_368 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_99_1706 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_109_Left_356 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_55_558 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5348__A1 core_0.execute.alu_mul_div.div_cur\[11\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_153_722 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_137_284 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_23_400 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_35_271 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_23_411 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_35_282 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_23_422 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_212_3056 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_152_287 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_23_455 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_51_764 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput108 net108 o_instr_long_addr[0] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_50_263 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xoutput119 net119 o_mem_addr[12] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_195_18 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4174__I2 core_0.ew_reg_ie\[2\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_121_696 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_130_2077 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_184_2719 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_56_1182 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_120_195 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4150_ core_0.dec_l_reg_sel\[0\] _0769_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XPHY_EDGE_ROW_118_Left_365 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_208_734 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput90 net90 dbg_r0[11] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_128_34 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_128_45 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6076__A2 _2009_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4081_ _0700_ _0594_ _0701_ _0702_ _0703_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai211_4
XANTENNA__4087__A1 net95 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_207_266 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4087__B2 _0708_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5823__A2 _2215_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_108_1813 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_223_3185 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_163_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_222_247 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7025__A1 _2567_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7840_ _0033_ clknet_leaf_70_i_clk core_0.fetch.out_buffer_data_instr\[17\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_188_652 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5036__B1 _1443_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_842 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_53_64 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5587__A1 _1987_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_175_302 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_230_280 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7771_ core_0.decode.i_instr_l\[8\] _1315_ _3842_ _3845_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__nor3_2
X_4983_ core_0.execute.alu_mul_div.i_mod _1432_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_19_706 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_74_801 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_175_335 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_195_2848 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6722_ _2977_ _3021_ _3032_ _0260_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XPHY_EDGE_ROW_127_Left_374 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_58_374 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3934_ _0567_ _0568_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_86_683 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_216 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7328__A2 _2434_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_129_763 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_18_249 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_116_402 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5339__A1 core_0.execute.alu_mul_div.div_cur\[9\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_73_344 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6653_ core_0.execute.rf.reg_outputs\[7\]\[12\] _2962_ _2984_ _2991_ vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_160_65 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_156_593 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_772 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6000__A2 _2390_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8275__CLK clknet_leaf_26_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5604_ _1652_ _2005_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_73_388 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_160_87 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4011__A1 core_0.execute.rf.reg_outputs\[7\]\[7\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_116_457 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_160_98 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_240_Right_240 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
X_6584_ core_0.ew_submit net20 _2929_ _2934_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_4
XFILLER_0_42_731 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_30_873 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_119_1942 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_54_591 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8323_ _0499_ clknet_leaf_83_i_clk core_0.dec_rf_ie\[3\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5535_ core_0.execute.mem_stage_pc\[3\] _1961_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__6839__A1 _2983_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_8254_ _0430_ clknet_leaf_24_i_clk core_0.execute.sreg_scratch.o_d\[4\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5466_ _1233_ _1894_ _1900_ _1809_ _1901_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XANTENNA__7500__A2 _3640_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_4417_ _1021_ _0860_ _0946_ _1022_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XPHY_EDGE_ROW_136_Left_383 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
X_7205_ _1381_ net202 _3392_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__5511__A1 core_0.execute.alu_mul_div.div_cur\[0\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
X_8185_ _0361_ clknet_leaf_123_i_clk core_0.execute.alu_mul_div.mul_res\[11\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_2
X_5397_ core_0.execute.alu_mul_div.div_cur\[4\] _1812_ _1841_ _1842_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_10_661 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4348_ core_0.fetch.pc_flush_override core_0.decode.i_flush _0965_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__or2_2
X_7136_ core_0.execute.alu_mul_div.mul_res\[15\] _3342_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_226_531 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_226_553 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7067_ _1372_ _3185_ _3278_ _3279_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4279_ _0888_ _0896_ _0897_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_214_715 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_185_84 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_185_95 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_214_737 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6018_ _1644_ _2300_ _1624_ _1549_ _2408_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_1
XTAP_TAPCELL_ROW_2_532 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4173__S1 _0768_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_241_556 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_83_1507 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7567__A2 core_0.execute.pc_high_out\[0\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_38_973 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_139_516 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_145_Left_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_166_302 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_330 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_609 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7969_ _0146_ clknet_leaf_45_i_clk core_0.execute.mem_stage_pc\[4\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_166_313 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_194_633 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_352 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_159_2423 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_167_858 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_77_672 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_64_311 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_204_69 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_119_240 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7537__B core_0.execute.prev_sys vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_80_804 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_190_861 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4002__A1 _0565_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_64_399 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_17_271 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_17_282 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5057__B _1460_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5750__A1 _1715_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_94_1636 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_150_769 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_594 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4305__A2 _0833_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5502__A1 _1908_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6550__I0 net117 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_469 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_236_317 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_229_66 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7255__A1 net85 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_217_575 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_205_715 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_189_416 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_204_247 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7007__A1 core_0.execute.alu_mul_div.mul_res\[4\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_252 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4915__I _1378_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_87_414 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_245_98 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7558__A2 _1953_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5569__A1 _1419_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_650 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_56_801 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_68_661 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_514 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_74_119 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_103_1743 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8298__CLK clknet_leaf_48_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_103_1754 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4241__A1 _0824_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_28_536 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_114_69 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_145_519 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_200_497 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_185_699 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7447__B _3553_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_83_664 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_172_349 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_71_837 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_174 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_153_552 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_731 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_113_405 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_126_799 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_180_360 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xrebuffer1 _0548_ net226 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_125_276 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_190_2789 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_70_369 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_140_213 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_180_382 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_58_1211 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_5320_ _1556_ _1557_ core_0.execute.alu_mul_div.div_cur\[1\] _1768_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_140_257 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_594 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_239_122 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_436 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_228_807 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6577__I _2929_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7494__A1 _1430_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5251_ _1644_ _1600_ _1700_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__6297__A2 _2642_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4202_ core_0.fetch.out_buffer_data_instr\[28\] _0821_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_114_1883 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_139_66 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5182_ _1446_ _1629_ _1630_ _1631_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XTAP_TAPCELL_ROW_225_3214 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_208_531 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7246__A1 net84 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6049__A2 _2279_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4133_ _0747_ _0751_ _0752_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_223_501 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7797__A2 _3778_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_208_597 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4064_ _0684_ _0685_ _0686_ _0687_ _0688_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_4
XTAP_TAPCELL_ROW_143_2224 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_64_41 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_223_545 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_3_66 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_3_88 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_69_1340 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_207_2991 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_64_85 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_195_408 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_210_217 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_64_96 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7823_ _0016_ clknet_leaf_60_i_clk core_0.fetch.out_buffer_data_instr\[0\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_148_313 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_149_836 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_35_932 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_149_858 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6221__A2 _2606_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_176_644 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7754_ _3829_ _3830_ _0494_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4232__A1 _0824_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4966_ _1400_ _0604_ _1420_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_236_3343 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_19_536 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_631 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_191_614 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_190_102 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6705_ core_0.execute.rf.reg_outputs\[5\]\[0\] _3022_ _3016_ _3023_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3917_ net94 _0521_ _0538_ _0552_ _0553_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai22_4
XANTENNA__5980__A1 _1601_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_62_804 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7685_ _1090_ _1095_ _1084_ _3785_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_191_658 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4897_ core_0.execute.alu_mul_div.cbit\[1\] _1364_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
X_6636_ _2936_ _2977_ _2978_ _0228_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_73_174 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_766 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_144_563 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_154_2364 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_131_202 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5732__A1 _1765_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6567_ _2924_ _0213_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_42_561 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_263 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8306_ _0482_ clknet_leaf_76_i_clk net191 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_4
XFILLER_0_14_274 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7804__C _1279_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5518_ net104 _1948_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_6498_ _2287_ _1719_ _2286_ _2876_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__7485__A1 _1392_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_246_604 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8237_ _0413_ clknet_leaf_34_i_clk core_0.execute.sreg_irq_pc.o_d\[9\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_7_602 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_5449_ _1796_ _1801_ _1886_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__4299__A1 core_0.fetch.prev_request_pc\[0\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3904__I core_0.dec_r_reg_sel\[1\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_218_317 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_246_648 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8168_ _0344_ clknet_leaf_84_i_clk net90 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_4
XANTENNA__7237__A1 _1414_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7237__B2 _1431_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7119_ _1222_ _3227_ _3327_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_8099_ _0275_ clknet_leaf_113_i_clk core_0.execute.rf.reg_outputs\[4\]\[6\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_199_725 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_165_2493 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_153_Left_400 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_199_769 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_198_279 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_97_767 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_167_622 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_57_i_clk_I clknet_4_14__leaf_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_179_482 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6212__A2 _1758_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_139_346 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_96_288 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4223__A1 _0726_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_182_603 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_127_519 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_154_305 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_42_1012 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_231_34 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_64_141 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_65_664 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5971__A1 _1458_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_92_450 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_37_366 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5971__B2 _1457_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_166_198 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_182_647 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_231_67 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_686 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_147_390 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_837 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_174 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_135_541 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7712__A2 _0514_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5723__A1 _1124_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5184__C1 _1606_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_80_667 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_135_596 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_162_382 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_123_769 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_33_594 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_122_257 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_122_279 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7476__A1 net210 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_255 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6523__I0 _2893_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_237_626 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_85_18 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7228__A1 net82 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_53_1152 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_18_34 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_109_58 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_245_670 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7779__A2 _3766_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_189_202 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_88_734 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_220_3155 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4462__A1 _1038_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_189_279 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_177_419 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_87_233 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_198_780 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_197_290 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_47_108 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7400__A1 _3547_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4820_ core_0.decode.i_instr_l\[8\] _1317_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__4214__A1 _0724_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_32_902 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_118_508 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_200_272 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_158_688 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_192_2818 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_7_205 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_145_316 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_173_625 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4751_ _0828_ _1238_ _1276_ _0045_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_44_804 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_64_1281 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5962__A1 _1195_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_16_506 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5476__I _1908_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_56_675 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_126_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_71_623 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4682_ _1236_ _1237_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA__5409__C _1822_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7470_ net37 _3621_ _3622_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_114_703 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_71_667 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6421_ _2069_ _2799_ _2800_ _2801_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_40_990 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5714__A1 _1714_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_116_1901 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_70_166 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_231_3284 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6352_ _2626_ _2733_ _2734_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__5190__A2 _1631_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_594 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_70_199 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_113_279 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5303_ core_0.execute.alu_mul_div.div_cur\[14\] _1713_ _1751_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_6283_ _2113_ _2499_ _2667_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_12_789 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_8022_ _0199_ clknet_leaf_35_i_clk net126 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5234_ net188 net204 _1460_ _1683_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_4
XFILLER_0_227_136 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_209_851 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7640__B _1216_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5165_ core_0.execute.rf.reg_outputs\[5\]\[7\] _1604_ _1605_ core_0.execute.rf.reg_outputs\[7\]\[7\]
+ _1606_ core_0.execute.rf.reg_outputs\[3\]\[7\] _1614_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XANTENNA__6690__A2 _3000_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_166_53 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_208_383 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4116_ core_0.execute.pc_high_out\[1\] _0732_ _0736_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_0_223_320 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5096_ _0789_ core_0.execute.rf.reg_outputs\[4\]\[15\] _0779_ _1545_ vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_75_95 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4555__I core_0.decode.oc_alu_mode\[2\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4047_ core_0.execute.rf.reg_outputs\[6\]\[4\] _0661_ _0662_ core_0.execute.rf.reg_outputs\[5\]\[4\]
+ core_0.execute.rf.reg_outputs\[4\]\[4\] _0663_ _0672_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi222_2
XFILLER_0_78_200 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_223_375 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4453__A1 core_0.decode.i_instr_l\[6\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_168_408 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_78_244 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_91_72 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_78_277 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_176_430 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_182_96 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7806_ _0773_ _1134_ _3868_ _1279_ _0508_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_149_655 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_148_143 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_93_236 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5998_ core_0.execute.alu_mul_div.div_cur\[2\] _0800_ _2389_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_191_400 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_46_130 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7737_ net182 core_0.decode.i_imm_pass\[13\] _1063_ _3820_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__5953__A1 _2242_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4949_ _1381_ net215 _1408_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_74_450 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_164_647 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_62_601 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_461 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_686 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_163_135 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4220__A4 _0838_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_117_541 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_174 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_34_325 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7668_ core_0.dec_sreg_jal_over _1062_ _3771_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_7_772 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_191_488 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_10_629 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_132_500 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_807 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_62_667 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6619_ net25 _1148_ _2964_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4508__A2 core_0.decode.i_instr_l\[2\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7599_ core_0.execute.pc_high_buff_out\[6\] _3681_ _3717_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_104_235 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5181__A2 net219 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_15_594 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7458__A1 net37 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_91_1606 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_167_2511 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_30_597 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_167_2522 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6130__A1 _1601_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_246_478 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_218_169 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6681__A2 _3006_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_199_500 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_226_34 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_215_854 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_214_342 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4465__I core_0.decode.oc_alu_mode\[6\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7630__A1 _0733_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_199_555 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6433__A2 _2501_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_89_1579 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_226_89 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_214_397 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_18_729 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_202_559 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4995__A2 _0767_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_167_430 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_85_737 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6197__A1 net85 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6197__B2 _2537_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_195_772 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5244__I0 net189 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7980__CLK clknet_leaf_43_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_178_2651 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_84_247 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_38_642 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_100_1713 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_128_839 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_194_271 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_653 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_167_496 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4747__A2 _1238_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_26_804 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_127_338 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5944__B2 core_0.execute.pc_high_out\[1\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_65_461 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_154_146 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5229__C _1559_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_53_634 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_37_196 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_182_477 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7697__A1 _1038_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_151_831 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_40_306 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_151_842 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_40_317 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_177 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5172__A2 _1620_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_339 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_111_717 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_96_28 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_104_780 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_110_238 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_209_103 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_209_3017 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_189_2780 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_111_1842 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4132__B1 _0745_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7460__B _3541_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6672__A2 _2999_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_237_489 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_225_629 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_218_681 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_127_2038 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_136_34 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_206_865 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_136_45 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7621__A1 _3732_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6970_ _3176_ _3189_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_136_78 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_220_323 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6975__A3 _3193_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_66_1310 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_204_2961 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_5921_ _1625_ _1592_ _2312_ _2313_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_88_564 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_243_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6804__B _3072_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_76_737 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6188__A1 core_0.ew_data\[6\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5852_ core_0.dec_sreg_jal_over _2245_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_3
XFILLER_0_76_748 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_236 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_185_260 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_29_642 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_122_1971 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_4803_ _1038_ _1307_ _1308_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4738__A2 _1253_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_28_130 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5935__A1 _1480_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_122_1982 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_173_422 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_61_86 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5783_ _1711_ _2183_ _2184_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_146_647 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_233_3313 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_8_558 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7522_ _0615_ _3640_ _3656_ _0436_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_4734_ core_0.fetch.out_buffer_data_instr\[21\] net51 _1246_ _1268_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_138_2167 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_145_168 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_173_488 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_667 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_32_807 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__7688__A1 _1098_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7453_ _3563_ net75 _3553_ _3607_ _3608_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_4665_ core_0.execute.alu_mul_div.comp _0804_ _1220_ _0754_ _1221_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__oai211_4
XTAP_TAPCELL_ROW_151_2323 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6404_ _2753_ _2785_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_31_339 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_141_352 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5163__A2 net219 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_380 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_12_520 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6360__A1 _1568_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7384_ _0720_ _3544_ _3545_ _3550_ _3551_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_4596_ core_0.ew_data\[4\] core_0.ew_data\[12\] _1150_ _1163_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_114_588 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6335_ core_0.execute.sreg_priv_control.o_d\[10\] _1386_ _2577_ core_0.execute.sreg_irq_pc.o_d\[10\]
+ _2718_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_177_30 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6266_ core_0.execute.alu_mul_div.div_cur\[8\] _0800_ _2651_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_8005_ _0182_ clknet_leaf_54_i_clk core_0.ew_data\[4\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_2
XTAP_TAPCELL_ROW_244_3442 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_5217_ _0771_ _0773_ core_0.execute.rf.reg_outputs\[5\]\[2\] _1666_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__and3_1
XANTENNA__6663__A2 _2996_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_216_629 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6197_ net85 _2531_ _2582_ _2537_ _2583_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_215_117 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_149_2296 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_215_139 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5148_ _1578_ _1594_ _1596_ _1597_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA_input22_I i_mem_data[10] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_98_306 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6415__A2 _2486_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_162_2452 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_5079_ _1467_ net182 _1528_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_4
XANTENNA__4426__A1 net72 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_224_695 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_212_857 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_168_216 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_211_345 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6714__B _3016_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_94_512 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_94_523 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6179__A1 _2281_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_149_452 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_225 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_177_772 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_247 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_192_720 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_136_102 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_176_271 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4729__A2 _1238_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_149_496 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_94_589 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_163 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_23_787 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_152_628 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_35_656 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_117_360 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7545__B _1206_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_152_639 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_453 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_155 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_151_138 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3952__A3 _0544_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_133_842 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_EDGE_ROW_185_Right_185 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_34_177 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_22_317 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_173_2592 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_105_555 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_output90_I net90 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_120_514 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5065__B _1459_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_30_372 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_30_383 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_246_220 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_101_772 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6654__A2 _2990_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_50_1111 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4665__A1 core_0.execute.alu_mul_div.comp vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5862__B1 _2250_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_237_66 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5862__C2 _2254_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4409__B _0970_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_89_306 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_199_330 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7603__A1 core_0.execute.pc_high_out\[6\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6406__A2 _1386_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_199_352 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_199_374 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_106_26 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_199_385 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_704 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_737 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_230_687 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_48_1084 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_174_219 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_73_718 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_155_422 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_26_601 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_61_1240 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_183_764 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_31_34 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_122_47 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_122_58 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_143_617 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6590__A1 _2930_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_5_517 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_170_403 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_807 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_215_3087 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3943__A3 _0518_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_13_306 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_215_3098 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_80_272 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_152_Right_152 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_151_650 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6342__A1 _2244_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5145__A2 _1585_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_123_352 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_4450_ core_0.decode.i_instr_l\[2\] _1045_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_4
XFILLER_0_229_209 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7876__CLK clknet_leaf_83_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4381_ core_0.fetch.prev_request_pc\[9\] _0992_ _0993_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__6893__A2 _3130_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6120_ _2014_ _2507_ _2013_ _2508_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_21_394 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_193_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7190__B core_0.execute.alu_mul_div.div_res\[14\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5703__B net211 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6645__A2 _2983_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6051_ _2403_ _2407_ _2440_ _2360_ _2441_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_225_426 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_72_1380 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4656__A1 core_0.dec_jump_cond_code\[4\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5002_ _1450_ _1451_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_147_66 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5422__C _1838_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_206_651 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4408__A1 _0959_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_221_621 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_233_492 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__7070__A2 _3177_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_221_654 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4959__A2 _0626_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6953_ core_0.execute.alu_mul_div.mul_res\[0\] _3155_ _3173_ _3174_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_49_715 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_221_665 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_178_558 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_72_63 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5904_ _2294_ _2295_ _2296_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_6884_ core_0.execute.rf.reg_outputs\[1\]\[13\] _3114_ _3124_ _3125_ vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_48_247 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_76_556 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_8_311 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_64_707 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_118_102 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_409 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5835_ _2203_ _2226_ _2230_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_118_113 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_729 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_17_612 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_17_623 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_63_228 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_366 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5766_ _2166_ _2167_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_91_559 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5384__A2 _1811_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_44_431 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7505_ _3639_ _3646_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA__7365__B _3495_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4717_ _1257_ _1237_ _1258_ _0029_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_16_155 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_115_842 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_32_615 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5697_ _1123_ _1934_ net211 _1720_ _2098_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai211_2
XTAP_TAPCELL_ROW_20_757 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_161_458 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_177 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7436_ _0626_ _3544_ _3545_ _3593_ _3594_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_32_659 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5136__A2 _1584_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_75_1409 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6333__A1 core_0.execute.alu_mul_div.div_cur\[10\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
X_4648_ core_0.execute.sreg_jtr_buff.o_d\[0\] _0731_ _1206_ _1207_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_0_4_583 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_142_683 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_31_169 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_4_594 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6884__A2 _3114_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7367_ net204 _3495_ _3496_ _3536_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_4579_ _1154_ net148 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_188_84 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4895__A1 core_0.execute.alu_mul_div.cbit\[0\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6318_ _2286_ _1789_ _1576_ _1455_ _2638_ _2701_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_0_229_765 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7298_ _1414_ core_0.execute.sreg_irq_pc.o_d\[13\] _1424_ _1431_ _1736_ _3474_ vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XANTENNA__6709__B _3016_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_229_776 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6636__A2 _2977_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6249_ _2040_ _2633_ _2634_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4647__A1 _1172_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_243_212 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_99_615 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_99_648 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_207_58 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_224_481 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_212_621 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_98_147 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_196_311 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_86_1549 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_28_846 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_211_142 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5072__A1 _1467_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_196_344 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_95_832 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_67_556 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_269 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_578 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_137_422 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_175_2610 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_94_375 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_48_781 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_94_397 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_125_617 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_137_488 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_192_594 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_180_734 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_23_615 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_570 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3925__A3 _0549_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_103 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_330 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_152_469 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_648 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6324__A1 _2123_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5127__A2 _1492_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_97_1678 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6875__A2 _3114_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_120_322 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_132_193 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_219_242 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_235_702 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_219_253 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_186_2750 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_207_404 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4918__I net178 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_207_415 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4638__A1 net189 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_207_437 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_188_801 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_26_34 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_89_136 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_187_300 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_215_492 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_203_632 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_187_311 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7052__A2 _1451_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5063__A1 _1508_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_201_2920 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_58_523 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_221_Right_221 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
X_3950_ _0568_ core_0.execute.rf.reg_outputs\[3\]\[12\] _0549_ _0583_ vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_0_147_208 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_86_865 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_106_1785 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_128_411 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_175_539 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_46_718 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_217_3116 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_156_731 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_45_206 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3881_ _0516_ _0517_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_58_589 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_128_444 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_155_230 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5620_ _2018_ _2020_ _2021_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_73_548 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_155_252 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_26_431 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_109_680 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_170_211 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5551_ core_0.execute.mem_stage_pc\[9\] _1957_ _1964_ _1971_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_26_475 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_135_2137 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_206_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_53_272 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4502_ _1071_ _1073_ _1092_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_0_13_125 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5118__A2 _1566_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6315__A1 _2045_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_170_266 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8270_ _0446_ clknet_leaf_22_i_clk core_0.execute.sreg_irq_flags.o_d\[4\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_14_659 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5482_ _1909_ _1915_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_13_158 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7221_ _1414_ core_0.execute.sreg_irq_pc.o_d\[3\] _1401_ _1431_ _1736_ _3407_ vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi221_4
X_4433_ _0745_ net114 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__6866__A2 _3107_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4877__A1 _0830_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8054__CLK clknet_leaf_103_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7152_ _1375_ _3355_ _3356_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4364_ core_0.fetch.prev_request_pc\[12\] _0954_ _0979_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_228_3245 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_10_865 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6103_ _2488_ _2489_ _2490_ _2491_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__6618__A2 _2961_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4295_ core_0.fetch.out_buffer_valid _0840_ _0913_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7083_ _3177_ _3292_ _3293_ _0360_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_225_212 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4629__A1 core_0.execute.alu_flag_reg.o_d\[4\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_158_98 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_241_3401 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7291__A2 _3467_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6034_ _1121_ _2421_ _2423_ _1107_ _2424_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XTAP_TAPCELL_ROW_146_2266 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_197_108 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xrebuffer11 net232 net233 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlya_2
XFILLER_0_174_75 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7043__A2 _3181_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7985_ _0162_ clknet_leaf_29_i_clk core_0.execute.prev_pc_high\[4\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_13_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6264__B _0798_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_178_333 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_221_451 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5054__A1 _1466_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_194_804 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_221_473 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_89_692 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_25_816 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6936_ _1915_ _1559_ _3156_ _3157_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_193_303 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_119_411 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_190_63 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_119_422 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_239_3385 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_193_347 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_190_74 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6867_ core_0.execute.rf.reg_outputs\[1\]\[5\] _3114_ _3112_ _3116_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_49_589 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_147_742 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_9_653 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_81_1479 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_5818_ _2213_ _2215_ _2216_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__7807__C _1132_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6798_ core_0.execute.rf.reg_outputs\[3\]\[8\] _3070_ _3072_ _3076_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_8_163 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_119_488 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_162_723 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_174 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_697 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_762 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_91_378 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_157_2395 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_5749_ _2010_ _2013_ _2149_ _2150_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_2
XANTENNA__3907__I _0518_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_106_149 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_161_244 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_60_732 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_115_650 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_44_283 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5109__A2 _1557_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_170_2551 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_32_445 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7419_ core_0.execute.sreg_irq_pc.o_d\[6\] _3543_ _3579_ _3580_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__6857__A2 _3108_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output176_I net176 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_629 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_4_391 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_217_702 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_102_399 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6609__A2 core_0.ew_data\[3\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7806__A1 _0773_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7282__A2 _3391_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4096__A2 _0535_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5293__A1 _1172_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_5_574 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5997__C _1432_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_181_2680 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_234_34 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_212_440 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_197_642 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_87_629 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_127_i_clk_I clknet_4_1__leaf_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6242__B1 _2133_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_86_128 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_234_89 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5596__A2 _1665_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6793__A1 _2967_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_196_174 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_68_865 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_184_314 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_55_504 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6902__B _3124_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_45_1054 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_137_241 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5348__A2 _1752_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_137_274 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_192_380 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_125_436 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_192_391 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_152_255 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_2_306 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_212_3057 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_2_317 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_180_597 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_51_776 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput109 net109 o_instr_long_addr[1] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_133_480 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_489 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_11_629 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_50_275 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4859__A1 core_0.decode.i_imm_pass\[5\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_10_128 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_130_2067 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4174__I3 core_0.ew_reg_ie\[3\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_130_2078 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_56_1183 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
Xoutput80 net80 dbg_pc[2] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
Xoutput91 net91 dbg_r0[12] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_235_521 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_207_212 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4080_ _0567_ core_0.execute.rf.reg_outputs\[3\]\[1\] net226 _0702_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_0_235_554 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_128_68 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_222_Left_469 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_37_66 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4087__A2 _0521_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5284__A1 core_0.dec_jump_cond_code\[4\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6481__B1 _2534_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_223_727 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_222_204 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_108_1803 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_179_108 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_108_1814 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_223_3186 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_188_620 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7025__A2 _3181_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_53_10 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_144_34 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6233__B1 _2577_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_156_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_176_804 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_59_832 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_203_484 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_77_139 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7770_ _1136_ _3844_ _0496_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_148_517 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_58_331 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5587__A2 _1549_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4982_ _1430_ _1431_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_187_174 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_148_539 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6721_ core_0.execute.rf.reg_outputs\[5\]\[7\] _3027_ _3031_ _3032_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_86_662 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_195_2849 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_3933_ _0516_ _0567_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_175_347 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_312 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6652_ _2979_ core_0.ew_data\[12\] _2980_ net24 _2990_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_0_190_317 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5339__A2 _1754_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_128_263 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_144_723 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_231_Left_478 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_6_634 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5603_ _1558_ _1652_ _2004_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_0_171_520 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6583_ _0785_ _2190_ _2933_ _0220_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__4011__A2 _0529_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_54_570 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_171_553 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_119_1943 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_30_874 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_8322_ _0498_ clknet_leaf_83_i_clk core_0.dec_rf_ie\[2\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5534_ _1959_ _1956_ _1960_ _0144_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_103_108 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_131_417 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_188 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6839__A2 _3086_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_8253_ _0429_ clknet_leaf_15_i_clk core_0.execute.sreg_scratch.o_d\[3\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_42_798 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5465_ _1232_ _1899_ _1900_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_7204_ _3390_ _3391_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_246_808 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4416_ core_0.fetch.prev_request_pc\[2\] _1020_ _1021_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
Xclkbuf_leaf_124_i_clk clknet_4_1__leaf_i_clk clknet_leaf_124_i_clk vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_8184_ _0360_ clknet_leaf_123_i_clk core_0.execute.alu_mul_div.mul_res\[10\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_2
XANTENNA__5511__A2 _1812_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5396_ _0802_ _1841_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_111_174 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7135_ _2855_ _3181_ _3341_ _0364_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4347_ net77 _0964_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_3
XFILLER_0_238_381 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_240_Left_487 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
X_7066_ _1224_ _3276_ _3277_ _1371_ _3278_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_4278_ _0891_ _0893_ _0895_ _0896_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__5275__A1 _1451_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_241_502 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6017_ _2356_ _2406_ _2407_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_2_533 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_241_579 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_69_629 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_38_963 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_83_1508 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_38_974 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_68_128 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_194_601 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7968_ _0145_ clknet_leaf_11_i_clk core_0.execute.mem_stage_pc\[3\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5578__A2 _0177_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_77_640 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_167_837 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_179_697 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_77_662 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_159_2424 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_178_185 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_204_37 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6919_ net91 _3135_ _3139_ _3145_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_194_667 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_193_144 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_76_161 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7899_ _0090_ clknet_leaf_73_i_clk core_0.decode.i_imm_pass\[8\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_182_807 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_166_369 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_37_537 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_64_323 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_64_334 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_37_559 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_147_572 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6527__A1 core_0.ew_addr\[0\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_193_199 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_91_142 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_64_378 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_119_296 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4002__A2 _0524_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_134_244 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_135_767 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5750__A2 _1631_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_32_231 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_150_737 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_94_1637 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5852__I core_0.dec_sreg_jal_over vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_53_i_clk_I clknet_4_14__leaf_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5502__A2 _1934_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6550__I1 _2752_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6169__B _1686_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4468__I core_0.decode.oc_alu_mode\[7\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_2_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4069__A2 _0523_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_220 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_204_237 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_99_264 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7558__A3 _1205_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_158_815 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87_459 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5569__A2 _0735_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_157_325 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_158_859 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4777__B1 _0881_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_114_37 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_67_150 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_157_347 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_200_465 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_684 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_103_1744 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4241__A2 net47 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_83_621 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_632 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_95_492 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_184_166 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6518__A1 _2447_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_172_317 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_55_356 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_138_583 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_184_188 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_83_676 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_126_734 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_43_518 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_15_209 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_165_391 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_389 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7191__A1 _1748_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_181_851 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_36_592 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_197 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xrebuffer2 _0699_ net222 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_113_417 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_626 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_58_1212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_41_i_clk clknet_4_11__leaf_i_clk clknet_leaf_41_i_clk vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_24_798 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_140_269 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_239_134 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7494__A2 _0810_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5250_ _1693_ _1698_ _1452_ _1699_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or3_2
XFILLER_0_121_483 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_139_34 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4201_ _0816_ _0819_ _0820_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_114_1884 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_5181_ net99 net219 _1630_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_TAPCELL_ROW_225_3215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_56_i_clk clknet_4_11__leaf_i_clk clknet_leaf_56_i_clk vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__7246__A2 _3398_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4132_ core_0.execute.prev_pc_high\[5\] _0748_ _0745_ core_0.execute.prev_pc_high\[6\]
+ _0750_ _0751_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_0_236_863 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5257__A1 _1705_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4063_ _0567_ _0524_ _0527_ core_0.execute.rf.reg_outputs\[2\]\[3\] _0687_ vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_2
XTAP_TAPCELL_ROW_143_2225 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_155_66 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5430__C _1822_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_69_1341 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_207_2992 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_78_415 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_188_450 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4480__A2 _1045_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_204_782 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7822_ _0015_ clknet_leaf_18_i_clk core_0.execute.alu_mul_div.comp vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_4
XANTENNA__6757__A1 _2972_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8242__CLK clknet_leaf_43_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_176_612 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_35_933 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4768__B1 _0881_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_80_30 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7753_ core_0.decode.i_instr_l\[10\] _0514_ _1070_ _3830_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_46_301 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4965_ _1283_ _1419_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_164_807 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4232__A2 net45 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_176_667 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_58_172 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_171_76 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_175_155 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_236_3344 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_58_183 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6704_ _3020_ _3022_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_19_548 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6509__A1 _1719_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_3916_ _0545_ _0546_ _0550_ _0551_ _0552_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_0_19_559 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7684_ _1044_ _1112_ _1094_ _3784_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_4896_ _0804_ _1221_ _1363_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_73_142 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_15_690 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3991__A1 _0517_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6635_ core_0.execute.rf.reg_outputs\[7\]\[7\] _2962_ _1978_ _2978_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_74_698 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_116_233 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_186 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_154_2365 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_80_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6566_ core_0.dec_rf_ie\[3\] core_0.ew_reg_ie\[3\] _2201_ _2924_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_132_737 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_144_597 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_242 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_89_72 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_8305_ _0481_ clknet_leaf_74_i_clk net190 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_4
XFILLER_0_131_236 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5517_ _1947_ _0140_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6497_ _2872_ _1991_ _2874_ _2875_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_112_450 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8236_ _0412_ clknet_leaf_36_i_clk core_0.execute.sreg_irq_pc.o_d\[8\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xclkbuf_3_7_0_i_clk clknet_0_i_clk clknet_3_7_0_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_100_601 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_112_461 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5448_ _1884_ _1885_ _0133_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__7485__A2 _1206_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input52_I i_req_data[22] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6532__I1 _2390_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_112_483 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4299__A2 _0851_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4288__I _0835_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_246_638 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8167_ _0343_ clknet_leaf_87_i_clk net89 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_4
XFILLER_0_245_126 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_470 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5379_ _1767_ _1771_ _1826_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_196_95 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7118_ _1372_ _3324_ _3325_ _3326_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_100_689 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7820__C _1216_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_8098_ _0274_ clknet_leaf_113_i_clk core_0.execute.rf.reg_outputs\[4\]\[5\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5248__A1 _1124_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6445__B1 _2823_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_242_822 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_199_715 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_226_384 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7049_ _1911_ _1936_ core_0.execute.alu_mul_div.cbit\[1\] _3262_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_226_395 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_29_Right_29 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_241_321 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_198_214 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_165_2494 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_97_702 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_198_247 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_97_724 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_201_218 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6748__A1 _2951_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_139_314 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5956__C1 _2258_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_194_453 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_210_796 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_77_492 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_194 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_42_1013 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_154_317 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_166_177 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_805 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_108_734 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_147_380 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_182_659 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_181_136 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_38_Right_38 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__7173__A1 _3357_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5184__B1 _1605_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_162_372 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5723__A2 _1491_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6920__A1 _2990_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_150_523 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_702 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_122_247 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7476__A2 _2258_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_209_307 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8115__CLK clknet_leaf_111_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5487__A1 _1226_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_236_104 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_53_1153 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_236_159 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7228__A2 net81 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_218_863 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_47_Right_47 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__5239__A1 _1137_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_233_833 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_205_524 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_232_321 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_220_3156 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_87_212 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4462__A2 _1043_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_177_409 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_220_527 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_34_34 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6739__A1 core_0.ew_reg_ie\[4\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_201_730 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_198_792 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_199_Right_199 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_146_807 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_158_667 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4214__A2 net53 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_28_312 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_56_621 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5411__A1 core_0.execute.alu_mul_div.div_cur\[6\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4661__I _1218_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4750_ net59 _1241_ _1276_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_192_2819 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_185_486 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_157_177 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XPHY_EDGE_ROW_56_Right_56 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_64_1282 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_55_142 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_687 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_172_147 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4681_ _0813_ _1235_ _1236_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_0_43_326 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_126_553 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_12_660 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6420_ _1803_ _1501_ _2800_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_40_991 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5714__A2 _1501_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_114_737 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6911__A1 net102 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_116_1902 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_12_702 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7193__B _3357_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_114_759 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_231_3285 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5706__B net211 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6351_ _2432_ _2666_ _2732_ _2733_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_12_724 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_113_258 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_11_212 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5302_ core_0.execute.alu_mul_div.div_cur\[15\] _1711_ _1750_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_12_757 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__7467__A2 _3542_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6282_ _2133_ _2294_ _2666_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__5478__A1 _1909_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_8021_ _0198_ clknet_leaf_31_i_clk net125 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_59_97 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5233_ core_0.decode.oc_alu_mode\[1\] _1124_ _1682_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_209_830 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_65_Right_65 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
X_5164_ _1446_ _1611_ _1612_ _1613_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_0_236_660 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_75_41 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_242_107 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_52 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_166_65 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4115_ core_0.execute.pc_high_out\[2\] _0732_ _0735_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_4
X_5095_ core_0.execute.rf.reg_outputs\[2\]\[15\] _1438_ _1544_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_79_702 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_223_354 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4046_ _0671_ net205 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_223_365 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5650__A1 _1752_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_757 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7368__B _3516_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7805_ core_0.decode.i_instr_l\[14\] _3788_ _3866_ core_0.decode.i_instr_l\[11\]
+ _1132_ _3868_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_0_78_289 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5997_ core_0.execute.alu_mul_div.div_res\[2\] _0798_ _2385_ _2387_ _1432_ _2388_
+ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XPHY_EDGE_ROW_74_Right_74 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__5402__A1 _1374_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_149_667 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_166_Right_166 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_115_80 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_59_492 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7736_ _3819_ _0487_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_136_317 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4948_ _1301_ _1407_ _0111_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_148_177 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5953__A2 net201 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_191_434 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_46_142 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_46_153 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_19_367 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_304 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3964__A1 _0533_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_191_456 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_47_698 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7155__A1 _1372_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7667_ _3663_ _3770_ _0467_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_4879_ _0886_ _1321_ _1353_ _0096_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_191_467 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_635 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_117_553 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_61_112 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_564 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_117_575 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6618_ _2936_ _2961_ _2963_ _0225_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_7598_ core_0.execute.pc_high_out\[6\] _3715_ _3716_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__6902__A1 net98 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_144_383 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4508__A3 _1044_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_15_562 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_132_545 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6549_ _2576_ _2716_ _2915_ _0204_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_104_247 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_160_865 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_30_521 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_120_729 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_91_1607 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_219_616 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_83_Right_83 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__5469__A1 core_0.execute.alu_mul_div.div_cur\[15\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
X_8219_ _0395_ clknet_leaf_42_i_clk net76 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_4
XTAP_TAPCELL_ROW_167_2512 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_218_115 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6130__A2 _2309_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_218_137 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__8288__CLK clknet_leaf_48_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4141__A1 _0542_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_215_811 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_226_181 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_226_192 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_230_803 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7630__A2 _3729_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_201 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_241_151 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_202_516 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_69_212 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_214_387 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_202_527 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_187_729 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6961__I _3176_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_186_217 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_97_554 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_92_Right_92 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_85_716 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_242_34 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6197__A2 _2531_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_128_807 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__7394__A1 _1357_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_242_45 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_178_2652 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_242_56 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5244__I1 net205 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_133_Right_133 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_155_615 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_100_1714 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_182_412 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_139_188 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5944__A2 _1385_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4414__C _0963_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_37_142 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_93_760 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_37_164 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_65_473 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3955__A1 _0534_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_182_445 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7146__A1 _3175_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_170_629 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7697__A2 _1101_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_80_454 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_108_597 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_465 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5526__B _1284_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_123_556 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_150_353 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_150_364 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_96_18 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7449__A2 _3542_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_209_3018 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_189_2781 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_29_56 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_111_1843 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7460__C _3613_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_225_619 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6357__B _1061_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_224_107 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_218_671 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5880__A1 core_0.dec_sreg_jal_over vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_127_2039 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_205_321 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_206_855 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_205_376 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_45_66 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_233_696 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_66_1300 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_5920_ _1482_ _1620_ _2312_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_204_2962 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_220_346 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7188__B core_0.execute.alu_mul_div.div_res\[13\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_75_204 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_88_587 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5851_ _2243_ _2244_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XANTENNA__6188__A2 _2486_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_152_34 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_236_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_192_209 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_152_45 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_29_632 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4199__A1 _0724_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_100_Right_100 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
X_4802_ _1305_ _1307_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XTAP_TAPCELL_ROW_122_1972 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_172_Left_419 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
X_5782_ _1121_ _2087_ _2136_ _2139_ _2182_ _2183_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XTAP_TAPCELL_ROW_233_3303 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_56_451 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5935__A2 _2311_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_61_76 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_233_3314 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_7521_ core_0.execute.sreg_scratch.o_d\[10\] _3646_ _3651_ _3656_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_145_136 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4733_ _1267_ _0036_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_29_698 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6820__B _3083_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_138_2168 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_71_432 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_161_629 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7452_ net37 _3606_ _3607_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_4_710 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4664_ core_0.decode.i_flush _1051_ _1220_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__5699__A1 core_0.decode.oc_alu_mode\[12\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_9_66 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_151_2324 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6403_ _2360_ _2783_ _2784_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5436__B _1838_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_142_865 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7383_ _1357_ net72 _3546_ _3549_ _3550_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_4595_ _1162_ net141 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_52_690 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_77_1440 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_3_264 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6334_ _2360_ _2716_ _2717_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_40_863 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_286 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_565 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_101_228 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6265_ core_0.execute.alu_mul_div.div_res\[8\] _0798_ _2647_ _2649_ _1432_ _2650_
+ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XPHY_EDGE_ROW_181_Left_428 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_228_435 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_228_446 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_228_457 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8004_ _0181_ clknet_leaf_48_i_clk core_0.ew_data\[3\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_2
X_5216_ net97 _1492_ _1664_ _1665_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_4
XFILLER_0_86_73 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_177_86 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_110_795 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_177_97 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_244_3443 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6196_ _2578_ _2580_ _2581_ _2582_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_43_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_EDGE_ROW_235_Right_235 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_215_129 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_149_2297 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_5147_ _1595_ _1596_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XANTENNA__7612__A2 _3673_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_162_2453 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_224_674 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_223_151 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_193_74 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5078_ _0584_ _0589_ _1461_ _0591_ _1527_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai211_4
XANTENNA_input15_I i_core_int_sreg[8] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_169_718 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5623__A1 _2022_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_196_515 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4029_ _0516_ _0523_ _0526_ core_0.execute.rf.reg_outputs\[2\]\[6\] _0656_ vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_0_39_418 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_190_Left_437 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__6179__A2 _2565_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_177_762 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_149_464 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_183_209 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_137_615 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_192_732 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_164_423 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_19_142 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_207 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_191_220 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3937__A1 _0568_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_101 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_19_175 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__7128__A1 _2797_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7719_ net188 core_0.decode.i_imm_pass\[4\] _1946_ _3811_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_191_253 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_74_270 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_124_309 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_136_169 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_192_798 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_23_788 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_90_741 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_151_106 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_164_489 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5139__B1 _1443_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_62_443 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_570 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_605 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_62_465 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_173_2593 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_90_796 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_15_392 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output83_I net83 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6956__I _3176_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7300__A1 net76 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_30_395 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_101_784 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_219_468 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_50_1112 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4665__A2 _0804_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5862__A1 core_0.execute.pc_high_buff_out\[0\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5862__B2 core_0.execute.sreg_irq_flags.o_d\[0\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_202_Right_202 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_237_78 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_215_652 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7603__A2 _3673_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5614__A1 _2013_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_203_858 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_98_863 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_230_655 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_502 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_97_373 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_524 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_230_699 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7367__A1 net204 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8303__CLK clknet_leaf_76_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_174_209 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_48_1085 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_195_592 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_613 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_122_37 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3928__A1 net93 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_61_1241 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6640__B _1978_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_66_793 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6590__A2 core_0.ew_data\[0\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_31_46 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_155_489 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_5_529 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_182_286 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_26_679 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_142_139 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_215_3088 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_41_616 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_189 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_124_865 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_40_115 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1_702 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_80_295 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_137 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4380_ core_0.fetch.prev_request_pc\[8\] _0951_ _0992_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_22_863 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_111_559 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7471__B _3540_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5153__I0 _1560_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6050_ _2438_ _2439_ _2440_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_0_237_276 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input7_I i_core_int_sreg[15] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_186_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_72_1381 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_5001_ _1439_ _1448_ _1449_ _1450_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_56_54 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_206_630 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_87 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_206_663 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5605__A1 _1558_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_206_696 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_178_515 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6952_ core_0.decode.o_submit _3172_ _3173_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__5081__A2 _1527_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_48_204 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_53 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5903_ _1699_ _2133_ _2295_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_0_88_384 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6883_ _0722_ _3124_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_76_535 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_88_395 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_48_237 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_76_568 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5834_ _2202_ _2228_ _2229_ _0174_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_119_626 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_8_334 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_173_220 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5765_ _2163_ _2165_ _2166_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_17_646 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_118_169 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_134_629 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_146_489 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6042__S _2102_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7504_ net212 _3640_ _3645_ _0429_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_4716_ net42 _1253_ _1258_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_20_747 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_5696_ _1124_ _2019_ _2091_ _2092_ _2097_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_0_127_692 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_20_758 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_16_167 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7435_ _3563_ net87 _3553_ _3592_ _3593_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_126_191 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_4_551 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4647_ _1172_ _1205_ _1206_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_4
XANTENNA__7530__A1 _0563_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_71_295 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6333__A2 _1117_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_142_662 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_141_150 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4344__A1 net78 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_141_161 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7366_ _3528_ _3533_ _3534_ _3535_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4578_ core_0.ew_data\[3\] net157 _1154_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_97_61 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4895__A2 core_0.execute.alu_mul_div.cbit\[1\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_97_72 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_102_559 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6317_ _2698_ _2060_ _2699_ _2700_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_12_384 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7297_ _2825_ _3391_ _3473_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_228_243 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_244_703 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6248_ _2460_ _2632_ _2154_ _2149_ _2159_ _2633_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai221_4
XFILLER_0_216_416 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4647__A2 _1205_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6179_ _2281_ _2565_ _2566_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_99_627 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_197_802 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7597__A1 core_0.execute.pc_high_out\[5\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6725__B _3031_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8326__CLK clknet_leaf_81_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output121_I net121 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6217__S _2102_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_86_1539 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_28_847 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_67_502 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5072__A2 net184 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_196_356 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4280__B1 _0886_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_211_176 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_196_367 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7349__A1 _1458_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_0_494 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_137_401 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_94_365 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_175_2611 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_109_136 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_137_445 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_527 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_94_387 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7556__B _1216_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_164_242 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_35_432 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_125_629 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_106_843 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_23_627 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_796 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_22_115 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_865 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_97_1679 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4335__A1 _0892_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_123_i_clk_I clknet_4_1__leaf_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50_457 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_133_695 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_31_682 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_219_221 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_120_378 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_186_2740 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6088__A1 _2295_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_101_592 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4638__A2 net188 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_219_298 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_117_26 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_117_37 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_222_419 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6635__B _1978_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5063__A2 _1509_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_201_2921 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_203_699 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_97_181 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_48_i_clk_I clknet_4_12__leaf_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_86_855 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_97_192 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4810__A2 core_0.fetch.submitable vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_42_34 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_4_2__f_i_clk_I clknet_3_1_0_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_106_1786 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_85_354 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_217_3117 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_42_45 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3880_ _0515_ _0516_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_8
XTAP_TAPCELL_ROW_197_2880 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6012__A1 _1378_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7466__B _3541_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_171_702 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_183_562 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_38_281 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_741 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4574__A1 core_0.ew_data\[1\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5550_ _0996_ _1956_ _1970_ _0150_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_54_763 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_135_2127 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_115_139 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_135_2138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_5_348 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4501_ _1089_ _1091_ _0011_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5481_ _1911_ _1913_ _1229_ _1914_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_101_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_112_802 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_170_278 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_137 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7220_ _2440_ _3391_ _3406_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4326__A1 _0725_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4432_ _0748_ net113 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_151_481 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4877__A2 _1321_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_111_345 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_6_34 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7151_ _1838_ _1810_ _3355_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_4363_ _0934_ _0942_ _0945_ _0823_ _0978_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_0_10_855 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6079__A1 net223 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_228_3246 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6102_ core_0.execute.sreg_scratch.o_d\[5\] _2254_ _2249_ core_0.execute.pc_high_buff_out\[5\]
+ _2490_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_67_53 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7082_ core_0.execute.alu_mul_div.mul_res\[10\] _3177_ _3293_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__7815__A2 _1094_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_158_77 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4294_ core_0.fetch.prev_request_pc\[2\] _0860_ _0912_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__5826__A1 _2219_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_241_3402 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6033_ _2422_ _2366_ _2000_ _2423_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_4
XTAP_TAPCELL_ROW_146_2267 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_225_279 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_174_43 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__7579__A1 net203 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xrebuffer12 net232 net234 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlya_2
XFILLER_0_233_290 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7984_ _0161_ clknet_leaf_28_i_clk core_0.execute.prev_pc_high\[3\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__6251__A1 _1107_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5054__A2 net192 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_89_671 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_95_107 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_194_816 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6935_ _1915_ _1689_ _1230_ _3156_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_76_310 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_25_817 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_76_321 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_190_53 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_239_3375 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_239_3386 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6866_ _2961_ _3107_ _3115_ _0321_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_9_632 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_49_579 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6003__A1 core_0.ew_data\[2\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_64_527 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_76_387 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5817_ _0681_ _1444_ _2214_ _2215_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_6797_ _2977_ _3064_ _3075_ _0292_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_91_335 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_741 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7751__A1 _3663_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_161_201 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4565__A1 _0727_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5748_ _2018_ _2022_ _2149_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_91_368 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_161_212 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_44_251 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_157_2396 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_162_757 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_262 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_72_582 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5679_ _2069_ _2080_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__inv_2
XFILLER_0_161_267 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_161_278 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_170_2552 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_199_95 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_103_824 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_32_457 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7418_ net215 _3544_ _3545_ _3578_ _3579_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_0_4_381 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_660 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_799 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7349_ _1458_ _1990_ _3495_ _3519_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA_output169_I net169 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_490 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_130_687 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_229_552 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7806__A2 _1134_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_217_769 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4096__A3 _0536_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5293__A2 _1739_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6490__A1 _2360_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_5_575 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_181_2681 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_197_632 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_87_619 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6174__C _1479_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_86_107 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6242__A1 _1831_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5045__A2 net232 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_169_345 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_169_356 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_200_636 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6793__A2 _3064_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_855 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_185_838 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_354 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_28_719 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_138_732 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_45_1055 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_184_359 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_95_696 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_83_858 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_153_702 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_138_787 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_36_741 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_37 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_82_346 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4556__A1 _1078_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_125_448 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_140_407 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_212_3058 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_35_295 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_105_150 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_121_632 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_133_492 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4859__A2 _1341_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_130_2068 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_208_703 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_56_1184 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
Xoutput81 net81 dbg_pc[3] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA__5808__A1 _2205_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput92 net92 dbg_r0[13] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA__4865__S _1305_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_223_706 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6481__B2 net6 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_222_216 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_108_1804 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_223_3187 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_188_632 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5036__A2 _1438_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_231_772 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_187_142 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4981_ _1209_ _1430_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_203_496 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6784__A2 _3065_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_149_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_175_315 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4795__A1 _1301_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_354 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3932_ _0565_ _0541_ _0543_ core_0.execute.rf.reg_outputs\[5\]\[13\] _0566_ vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_4
X_6720_ _1963_ _3031_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_46_505 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5992__B1 _2295_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_719 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_527 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_173 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6651_ _2941_ _2988_ _2989_ _0232_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_46_549 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_160_34 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_rebuffer5_I _0879_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_4_Left_251 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
X_5602_ _2000_ _2002_ _2003_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_128_275 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_116_426 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_143_212 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_160_67 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6582_ net155 _2190_ _2933_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_42_722 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_119_1944 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_8321_ _0497_ clknet_leaf_80_i_clk core_0.dec_rf_ie\[1\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5533_ core_0.execute.mem_stage_pc\[2\] _1957_ _1217_ _1960_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_30_875 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_14_457 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_171_598 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8252_ _0428_ clknet_leaf_15_i_clk core_0.execute.sreg_scratch.o_d\[2\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5464_ _1751_ _1805_ _1899_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_41_276 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7203_ _1430_ _1381_ _3390_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_4415_ core_0.fetch.prev_request_pc\[1\] core_0.fetch.prev_request_pc\[0\] _1020_
+ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_2_863 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_169_76 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_8183_ _0359_ clknet_leaf_124_i_clk core_0.execute.alu_mul_div.mul_res\[9\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_111_142 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5395_ core_0.execute.alu_mul_div.div_cur\[3\] _1814_ _1817_ _1839_ _1840_ vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_0_245_308 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7134_ _3189_ _3340_ _3341_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4346_ _0883_ _0961_ _0962_ _0963_ net167 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XFILLER_0_238_393 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7065_ _1224_ _3226_ _3277_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4277_ _0892_ _0837_ _0894_ _0895_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_226_566 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_185_86 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5275__A2 _1456_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6016_ _2357_ _2405_ _2406_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_214_728 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_198_407 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_2_534 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_118_91 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_179_632 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_179_643 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_222_761 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_68_107 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6224__A1 core_0.execute.alu_mul_div.div_cur\[7\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_38_964 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_83_1509 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_178_142 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_179_665 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xclkbuf_3_3_0_i_clk clknet_0_i_clk clknet_3_3_0_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_7967_ _0144_ clknet_leaf_45_i_clk core_0.execute.mem_stage_pc\[2\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__6775__A2 _3041_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_221_282 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_49_343 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4786__A1 _1290_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_159_2425 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6918_ _2988_ _3130_ _3144_ _0344_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_166_348 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7898_ _0089_ clknet_leaf_69_i_clk core_0.decode.i_imm_pass\[7\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_49_387 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_65_836 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_9_440 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_76_173 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_119_242 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_147_551 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_92_633 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_135_702 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_65_858 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6849_ _2994_ _3087_ _3104_ _0315_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_147_562 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6527__A2 _2190_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_181_318 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__3918__I _0553_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_9_473 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_92_677 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_839 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_91_176 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4002__A3 _0527_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_17_262 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_220_37 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_33_766 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_32_243 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_552 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_32_265 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_405 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_690 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_94_1638 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_103_632 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_32_276 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_32_287 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_130_451 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_20_449 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_103_687 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_130_473 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5073__C _1461_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4710__A1 net40 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_183_2710 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_217_555 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_217_566 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_205_706 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_245_12 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4069__A3 _0526_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_204_205 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_245_56 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_4_6__f_i_clk clknet_3_3_0_i_clk clknet_4_6__leaf_i_clk vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__6215__A1 _2591_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_276 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_169_131 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_213_772 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87_438 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_169_142 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_169_153 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_200_411 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6913__B _3139_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_197_484 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4777__A1 core_0.fetch.prev_request_pc\[6\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4777__B2 net173 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_28_505 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_184_123 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_95_460 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_103_1745 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_28_527 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_28_549 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_644 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_172_307 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_55_346 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7715__A1 core_0.decode.i_imm_pass\[2\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_18 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4529__A1 _1037_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_125_201 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_817 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_125_212 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_71_839 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_83_699 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_126_757 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_711 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_130_26 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_181_863 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8194__CLK clknet_leaf_129_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_130_37 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xrebuffer3 _1641_ net223 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_130_59 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_140_215 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_180_384 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_58_1213 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_11_416 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_210_81 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4659__I _1216_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7494__A3 _2579_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4200_ _0725_ _0817_ _0818_ _0819_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_139_46 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5180_ _0776_ _1626_ _1627_ _1628_ _1629_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai211_4
XTAP_TAPCELL_ROW_114_1885 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_225_3216 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_4131_ core_0.execute.prev_pc_high\[5\] _0748_ _0749_ _0750_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__5257__A2 _1693_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5501__I0 net99 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4062_ _0567_ core_0.execute.rf.reg_outputs\[4\]\[3\] net229 _0686_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_223_525 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6095__B core_0.dec_mem_access vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_143_2226 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_147_Right_147 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__4608__B _0813_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_211_709 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_207_2993 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_69_1342 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_188_440 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7821_ _3769_ _3767_ _3878_ _0513_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_204_794 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6757__A2 _3042_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_203_282 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_35_934 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4768__B2 net169 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4964_ _1301_ _1418_ _0116_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_7752_ core_0.dec_jump_cond_code\[3\] _1062_ _3829_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_58_162 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_171_66 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6703_ _3020_ _3021_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XTAP_TAPCELL_ROW_236_3345 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_47_858 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3915_ _0534_ _0542_ _0544_ core_0.execute.rf.reg_outputs\[5\]\[15\] _0551_ vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_0_129_562 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_163_307 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_190_104 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4895_ core_0.execute.alu_mul_div.cbit\[0\] core_0.execute.alu_mul_div.cbit\[1\]
+ _1362_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__6509__A2 _1455_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7683_ _1128_ _3778_ _3779_ _3782_ _3783_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and4_1
XANTENNA__7706__A1 core_0.dec_mem_we vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_191_638 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_156_370 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6634_ _2930_ core_0.ew_data\[7\] _2976_ _2977_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_4
XFILLER_0_46_379 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_15_691 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_62_839 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_27_571 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_13_91 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7182__A2 _3373_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_144_543 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_190_159 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_27_582 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_172_863 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_154_2355 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5193__A1 _1603_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_116_267 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6565_ _2923_ _0212_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_154_2366 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_15_766 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_132_749 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8304_ _0480_ clknet_leaf_76_i_clk net189 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_4
X_5516_ core_0.de_jmp_pred core_0.decode.i_jmp_pred_pass _1946_ _1947_ vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__4940__A1 core_0.execute.sreg_long_ptr_en vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6496_ _1996_ _2085_ _2874_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_131_248 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4940__B2 _1391_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_73_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5447_ core_0.execute.alu_mul_div.div_cur\[11\] _1812_ _1841_ _1885_ vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_8235_ _0411_ clknet_leaf_43_i_clk core_0.execute.sreg_irq_pc.o_d\[7\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_100_613 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_140_793 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_58_Left_305 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_196_63 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5378_ core_0.execute.alu_mul_div.div_cur\[2\] _1811_ _1825_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_8166_ _0342_ clknet_leaf_88_i_clk net103 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_4
XANTENNA_input45_I i_req_data[16] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_227_842 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4329_ _0946_ _0947_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
X_7117_ _1225_ _3276_ _3325_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_8097_ _0273_ clknet_leaf_113_i_clk core_0.execute.rf.reg_outputs\[4\]\[4\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_242_801 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_226_352 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5248__A2 _1696_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7048_ _1222_ _3260_ _3261_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__6996__A2 _2436_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_114_Right_114 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_165_2495 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_242_856 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_241_333 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8067__CLK clknet_leaf_111_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_416 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_167_602 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6733__B _3031_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6748__A2 _3042_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output201_I net201 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_166_101 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_38_803 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_139_326 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4759__A1 core_0.decode.i_flush vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_67_Left_314 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_210_764 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_96_279 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5956__B1 _2265_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5956__C2 net105 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_194_465 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_166_156 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_167_679 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_92_430 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_42_1014 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_37_346 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_132 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_713 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_107_212 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_677 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_135_532 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_231_69 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_839 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5184__A1 core_0.execute.rf.reg_outputs\[5\]\[4\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_107_267 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5184__B2 core_0.execute.rf.reg_outputs\[7\]\[4\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_52_349 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_45_390 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_80_669 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_122_215 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6920__A2 _3130_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_162_384 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7283__C _1736_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_100_18 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_116_790 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_122_237 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4931__A1 _0722_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_76_Left_323 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_103_473 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_257 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6684__A1 _2977_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5487__A2 _1568_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_53_1143 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_229_190 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_53_1154 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_233_801 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_217_352 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5239__A2 _1451_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6436__A1 _1137_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_189_259 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_220_3157 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_85_Left_332 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_87_224 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_88_769 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6739__A2 _2934_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4942__I net204 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_87_279 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_200_241 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_158_657 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_185_454 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_29_836 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_200_263 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_123_i_clk clknet_4_1__leaf_i_clk clknet_leaf_123_i_clk vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__5411__A2 _1812_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_173_605 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_205_92 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_29_858 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_28_335 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_28_346 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_655 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_172_104 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_173_627 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_64_1283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_138_370 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_34 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_71_603 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_45 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4680_ _0721_ _0727_ _1168_ _1235_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_0_44_839 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_70_102 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_485 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_187 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_636 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_496 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6372__B1 _2577_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_12_661 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_113_204 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_114_727 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_126_587 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_40_992 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_116_1903 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6911__A2 _3135_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6350_ _2090_ _2728_ _2731_ _2732_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_113_226 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_180_181 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_94_Left_341 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_231_3286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_5301_ core_0.execute.alu_mul_div.div_cur\[15\] _1711_ _1749_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_EDGE_ROW_216_Right_216 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_11_224 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6281_ _2356_ _2664_ _2665_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_59_54 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_246 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5478__A2 _1592_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_8020_ _0197_ clknet_leaf_30_i_clk net124 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5232_ _1642_ _1680_ _1480_ _1681_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__6675__A1 _2956_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_227_105 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_121_292 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6818__B _3083_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5163_ net100 net219 _1612_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_224_801 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6427__A1 _1458_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4114_ core_0.execute.prev_pc_high\[3\] _0733_ _0734_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_208_363 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_75_64 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5094_ net94 _1492_ _1543_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__6978__A2 _3193_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_224_856 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4045_ _0664_ _0669_ _0670_ _0671_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_2
XANTENNA__5650__A2 _1567_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_78_224 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_182_43 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_195_207 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_79_769 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_204_591 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_148_101 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_182_76 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7804_ _0776_ _1134_ _3867_ _1279_ _0507_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_5996_ _1433_ _2386_ _0798_ _2387_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_47_622 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_96_i_clk_I clknet_4_6__leaf_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_148_145 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_176_465 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7735_ net181 core_0.decode.i_imm_pass\[12\] _1946_ _3819_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_176_476 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4947_ core_0.execute.sreg_priv_control.o_d\[5\] _1394_ _1406_ _1391_ _1407_ vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_24_90 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_163_104 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_176_487 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_346 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_148_189 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5884__S _2190_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7666_ _1414_ _3766_ _3769_ _3767_ _3770_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_4878_ core_0.decode.i_imm_pass\[14\] _1341_ _1353_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_62_625 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7155__A2 _1809_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_74_485 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7384__B _3545_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6617_ core_0.execute.rf.reg_outputs\[7\]\[4\] _2962_ _1978_ _2963_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_132_502 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_117_587 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_132_513 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7597_ core_0.execute.pc_high_out\[5\] core_0.execute.pc_high_out\[4\] _3695_ _3715_
+ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__6902__A2 _3135_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4508__A4 _1084_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_61_157 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_172_693 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_132_535 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4913__A1 _1375_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_104_237 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_160_855 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6548_ net131 _1985_ _2915_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_42_360 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_171_192 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_91_1608 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6479_ core_0.execute.alu_mul_div.div_res\[14\] _1114_ _1432_ _2858_ vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XANTENNA__5469__A2 _1711_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_8218_ _0394_ clknet_leaf_35_i_clk net75 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_4
XFILLER_0_219_628 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_112_281 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_167_2513 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_100_443 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4141__A2 _0544_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_246_469 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8149_ _0325_ clknet_leaf_107_i_clk core_0.execute.rf.reg_outputs\[1\]\[8\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_10_290 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6418__A1 _1088_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6969__A2 _3181_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7091__A1 core_0.execute.alu_mul_div.mul_res\[10\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_199_535 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_241_130 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_214_344 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_97_500 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_226_69 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_214_377 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_97_522 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_241_174 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_40_i_clk clknet_4_11__leaf_i_clk clknet_leaf_40_i_clk vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__5858__I net185 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_195_730 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4762__I _1283_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_195_741 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_69_279 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6182__C _1432_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_195_774 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_194_251 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_139_156 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_178_2653 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_210_594 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_194_262 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_38_644 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_155_627 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_100_1715 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_167_498 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_65_463 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_93_772 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_55_i_clk clknet_4_14__leaf_i_clk clknet_leaf_55_i_clk vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__3955__A2 _0535_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_26_839 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_80_411 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_182_457 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_136_863 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5157__A1 _0770_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5593__I _1491_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7697__A3 _1041_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_163_682 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_20_37 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_162_170 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4904__A1 _1369_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_80_477 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_150_321 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_40_319 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_33_360 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_60_190 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_150_387 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6657__A1 _2941_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8232__CLK clknet_leaf_43_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_209_3019 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_189_2782 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5542__B _1964_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_111_1844 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4132__A2 _0748_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7313__I _3398_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_218_661 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6409__A1 net75 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6409__B2 _2537_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5880__A2 _2270_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7082__A1 core_0.execute.alu_mul_div.mul_res\[10\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_221_804 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_66_1301 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_204_2963 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_118_i_clk_I clknet_4_6__leaf_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_216_80 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_76_706 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_17_720 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4672__I core_0.execute.alu_mul_div.cbit\[1\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_220_358 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_88_577 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_0_36 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5850_ core_0.dec_sreg_load core_0.dec_sreg_jal_over _2243_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_69_780 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7385__A2 _3543_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_791 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_158_465 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4801_ _1305_ _1306_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XANTENNA__4199__A2 net49 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_201_594 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_158_476 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_185_273 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_61_66 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5781_ _1988_ _2180_ _2181_ _2182_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XTAP_TAPCELL_ROW_122_1973 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_131_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_233_3304 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_229_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_29_666 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7520_ _0626_ _3640_ _3655_ _0435_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_139_690 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4732_ core_0.fetch.out_buffer_data_instr\[20\] net50 _1246_ _1267_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_84_783 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7137__A2 _1941_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_71_422 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_282 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_138_2169 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_161_619 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_28_198 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7451_ core_0.execute.mem_stage_pc\[12\] _3606_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_4663_ _1219_ net210 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_154_671 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_160_107 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_114_524 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_4_733 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_126_384 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5699__A2 _1553_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6402_ core_0.execute.alu_mul_div.div_cur\[12\] _2279_ _2782_ _2783_ vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_4
XANTENNA__6896__A1 _2946_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_151_2325 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_3_221 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_488 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_142_855 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_153_192 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4594_ core_0.ew_data\[3\] core_0.ew_data\[11\] _1150_ _1162_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_7382_ _3547_ _3548_ _3549_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_52_680 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_77_1441 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_101_72 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_101_207 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6333_ core_0.execute.alu_mul_div.div_cur\[10\] _1117_ _2713_ _2715_ _2716_ vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XANTENNA__5008__I core_0.decode.oc_alu_mode\[4\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6648__A1 _2941_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_12_588 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6264_ _1433_ _2648_ _0798_ _2649_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_177_43 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_86_41 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8003_ _0180_ clknet_leaf_54_i_clk core_0.ew_data\[2\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_2
X_5215_ _1658_ _1663_ _1664_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5452__B _1817_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6195_ core_0.execute.pc_high_buff_out\[7\] _2249_ _2534_ net14 _2581_ vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_TAPCELL_ROW_244_3444 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_209_672 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_209_683 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5146_ _1556_ _1557_ _1595_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_TAPCELL_ROW_149_2298 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_36_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_208_193 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7073__A1 _1367_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_224_664 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5077_ _1467_ net181 _1526_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_2
XTAP_TAPCELL_ROW_162_2454 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_79_522 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6820__A1 core_0.execute.rf.reg_outputs\[2\]\[1\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_211_314 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4028_ _0532_ _0540_ _0543_ core_0.execute.rf.reg_outputs\[5\]\[6\] _0655_ vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_4
XTAP_TAPCELL_ROW_88_1570 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_196_527 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_79_566 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_189_590 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_79_577 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_192_700 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5387__A1 _1374_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_136_104 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_137_627 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5979_ _1578_ _1532_ _1558_ _2370_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_75_772 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3937__A2 _0542_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7718_ _2246_ _0514_ _3810_ _0478_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_47_474 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_783 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_164_457 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7128__A2 _3328_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_47_496 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_35_636 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_118_863 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5139__A1 core_0.execute.rf.reg_outputs\[7\]\[8\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_23_789 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5627__B _2013_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6336__B1 _2534_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7649_ _1217_ _3757_ _0462_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_117_373 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_191_298 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_105_524 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_117_384 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_34_168 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6887__A1 _2994_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_173_2583 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_173_2594 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_105_579 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_842 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_132_387 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6639__B2 net35 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_30_363 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_246_200 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output76_I net76 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_219_436 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_246_244 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4114__A2 _0733_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5311__A1 core_0.execute.alu_mul_div.div_cur\[7\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4757__I _0726_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_50_1113 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_246_288 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5862__A2 _2249_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_199_310 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4693__S _1241_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_89_308 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_199_332 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_199_343 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_215_697 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_214_163 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5614__A2 _2014_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6811__A1 _2994_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7289__B net75 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_202_325 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_230_645 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_202_336 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_58_706 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_97_352 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_230_667 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_58_717 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_216 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7367__A2 _3495_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_48_1086 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_168_785 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4425__I0 core_0.fetch.prev_request_pc\[0\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6921__B _3139_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_452 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_155_446 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_61_1242 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_65_260 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3928__A2 _0521_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_183_777 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_422 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_65_282 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_142_107 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_108_362 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_41_606 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_80_241 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_215_3089 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6878__A1 _2986_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_53_477 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_80_263 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_124_855 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_41_628 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5550__A1 _0996_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_330 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_238_734 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6368__B _2279_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5272__B net211 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5302__A1 core_0.execute.alu_mul_div.div_cur\[15\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_72_1371 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_5000_ net88 _1446_ _1449_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_2
XTAP_TAPCELL_ROW_72_1382 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_56_66 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7055__A1 _2648_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_56_77 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_179_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_205_130 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_89_842 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6951_ _1088_ core_0.execute.alu_mul_div.comp _3164_ _3171_ _3172_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_4
XANTENNA__8128__CLK clknet_leaf_94_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_163_34 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_49_706 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_88_341 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_221_656 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_88_352 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_163_56 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5902_ _2293_ _2294_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XANTENNA__5081__A3 _1528_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6882_ _2990_ _3108_ _3123_ _0329_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__7358__A2 _2888_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_29_430 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5833_ net136 _2209_ _2229_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6831__B _3083_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_9_836 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_118_104 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_201_391 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_146_435 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8278__CLK clknet_leaf_26_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_9_858 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_57_772 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_158_295 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_22_Left_269 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_173_232 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5764_ _1754_ _2035_ _2164_ _2165_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_16_102 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5447__B _1841_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7503_ core_0.execute.sreg_scratch.o_d\[3\] _3641_ _3516_ _3645_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_72_753 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6318__B1 _1576_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4715_ core_0.fetch.out_buffer_data_instr\[13\] _1257_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_5695_ _2094_ _2095_ _1554_ _2096_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_173_298 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_20_748 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_71_263 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7434_ _3547_ _3591_ _3592_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4646_ core_0.dec_jump_cond_code\[4\] _1204_ _1205_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_31_116 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7530__A2 _3641_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_31_138 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_842 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4344__A2 _0883_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5541__A1 _1013_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4577_ _1153_ net147 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_188_53 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_4_585 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_12_330 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_102_527 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_7365_ _3528_ _3533_ _3495_ _3534_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_114_387 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_188_64 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_661 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_141_184 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_229_723 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6316_ _2698_ _2060_ _1121_ _2699_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_228_211 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_683 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7296_ _3469_ _3472_ _1395_ _0394_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__7294__A1 _2783_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_31_Left_278 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_110_571 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6247_ _2010_ _2013_ _2149_ _2632_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_0_216_428 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6178_ _2295_ _2547_ _2564_ _2565_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_0_243_269 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5129_ _1482_ _1568_ _1577_ _1531_ _1578_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_0_212_601 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_197_836 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_197_858 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_28_848 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_79_352 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_output114_I net114 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_211_144 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_200_807 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_211_155 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4280__A1 core_0.fetch.prev_request_pc\[13\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_94_311 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_184_508 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4280__B2 core_0.fetch.prev_request_pc\[14\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_196_379 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_184_519 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_40_Left_287 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_0_495 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_137_413 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_175_2612 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_48_772 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_164_221 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_82_539 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_63_720 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_94_399 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_109_159 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_180_703 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_282 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_422 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_800 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_811 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_124_107 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_164_276 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5780__A1 _1107_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_62_241 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_90_594 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_105_343 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7521__A2 _3646_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_127 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_105_365 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_120_302 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_121_836 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_132_162 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_121_858 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_31_694 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_30_182 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7285__A1 net74 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_219_244 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_186_2741 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_207_406 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_219_277 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_207_417 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5835__A2 _2226_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4638__A3 net191 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_234_247 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_234_258 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7588__A2 _3672_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5599__A1 _1676_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_188_836 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_187_313 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_202_133 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_58_503 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_201_2922 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_230_464 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_202_166 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_187_368 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_311 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_97_171 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_202_177 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_106_1787 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_217_3118 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_197_2881 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_39_761 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6012__A2 core_0.execute.sreg_irq_pc.o_d\[3\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_772 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_128_457 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_183_541 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4023__A1 core_0.execute.rf.reg_outputs\[7\]\[6\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_128_468 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_38_293 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5267__B _1705_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_143_416 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4574__A2 net157 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_6_839 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4171__B _0789_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5982__S _1558_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_54_775 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_115_129 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_135_2128 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_143_449 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_170_235 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_263 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_786 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_181 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4500_ _0514_ _1078_ _1090_ _1091_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_0_41_414 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5480_ _1909_ _1576_ _1912_ _1913_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_124_641 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_14_639 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4431_ _0733_ net111 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA_1 _1357_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4326__A2 net49 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_458 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_111_302 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5523__A1 core_0.decode.i_flush vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_111_313 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_74_1400 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_4362_ net75 _0977_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_2
X_7150_ _1980_ _0807_ _0366_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_158_34 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_158_45 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6101_ net12 _2260_ _2264_ core_0.execute.sreg_irq_pc.o_d\[5\] _2489_ vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_TAPCELL_ROW_228_3247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_7081_ _2053_ _3178_ _3289_ _3291_ _3292_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_4293_ _0909_ _0835_ _0910_ _0911_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_67_76 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_226_737 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_238_597 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_67_98 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6032_ _2002_ _2422_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_241_3403 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_226_748 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_225_258 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_146_2268 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7579__A2 _3675_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_83_53 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xrebuffer13 net232 net235 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlya_2
XFILLER_0_179_836 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7983_ _0160_ clknet_leaf_28_i_clk core_0.execute.prev_pc_high\[2\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_174_99 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_178_335 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_179_858 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_221_453 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6934_ _1223_ _1369_ _3153_ _3155_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_1
XTAP_TAPCELL_ROW_25_807 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_25_818 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_9_600 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_88_193 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_49_558 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6865_ core_0.execute.rf.reg_outputs\[1\]\[4\] _3114_ _3112_ _3115_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_92_804 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_239_3376 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_64_506 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_193_349 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6003__A2 _2209_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7200__A1 _1431_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5816_ _1655_ _1656_ _1657_ _2214_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_2
XANTENNA__4014__A1 _0533_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_147_766 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6796_ core_0.execute.rf.reg_outputs\[3\]\[7\] _3070_ _3072_ _3075_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_29_271 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_162_703 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_29_282 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_17_422 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_9_699 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_106_107 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4565__A2 _0947_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5747_ _1998_ _2146_ _2147_ _2148_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA__5762__A1 _1754_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_106_129 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_162_747 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_157_2397 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_60_734 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5678_ _2074_ _2075_ _2079_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__7503__A2 _3641_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_170_2553 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_7417_ _3563_ net84 _3553_ _3577_ _3578_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_0_115_685 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_130_611 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5514__A1 _1419_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_32_469 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_115_696 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4629_ core_0.execute.alu_flag_reg.o_d\[4\] _1186_ _1187_ core_0.dec_jump_cond_code\[1\]
+ core_0.dec_jump_cond_code\[2\] _1188_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_0_103_858 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_13_672 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7348_ _1719_ _2888_ _3518_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__7267__A1 _2690_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_12_193 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_130_699 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7279_ _2716_ _3393_ _3457_ _3458_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__4100__I _0720_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5817__A2 _1444_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_218_37 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_244_545 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_216_247 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_5_576 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6490__A2 _2859_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_231_206 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_231_228 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_225_792 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_197_611 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_181_2682 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4256__B _0813_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_212_453 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_240_773 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_234_69 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_240_795 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_200_626 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_200_648 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7567__B core_0.execute.pc_high_out\[2\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_67_344 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_184_338 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_208 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_45_1056 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_137_232 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7286__C _1735_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4005__A1 _0517_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_82_314 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_94_174 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_137_243 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_165_552 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_325 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_82_358 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4556__A2 _1092_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_153_758 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_51_712 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_263 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_211 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_663 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_212_3059 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_133_460 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4308__A2 _0843_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5505__A1 _1367_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50_244 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_161_791 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_128_Right_128 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_121_688 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_130_2069 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7258__A1 net86 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_56_1185 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
Xoutput82 net82 dbg_pc[4] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
Xoutput93 net93 dbg_r0[14] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_128_37 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_207_225 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4867__I0 _0844_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6481__A2 _2579_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7321__I core_0.execute.alu_flag_reg.o_d\[0\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_108_1805 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_222_228 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_223_3188 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7430__A1 _0637_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6233__A2 _1386_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_53_56 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_144_69 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4980_ _1419_ _1429_ _0121_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_230_272 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_176_839 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3931_ _0532_ _0565_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_19_709 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5992__A1 _1676_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_86_664 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_187_198 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_86_675 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_175_349 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_129_755 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6650_ core_0.execute.rf.reg_outputs\[7\]\[11\] _2962_ _2984_ _2989_ vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_128_243 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5601_ _2001_ _1599_ _2002_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_156_585 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_80_1470 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_211_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6581_ _2932_ _0219_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_160_79 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6941__B1 _1761_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_128_298 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_26_263 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_6_658 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8320_ _0496_ clknet_leaf_86_i_clk core_0.dec_rf_ie\[0\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5532_ net80 _1959_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_30_876 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_119_1945 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_81_380 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_131_419 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_41_244 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8251_ _0427_ clknet_leaf_15_i_clk core_0.execute.sreg_scratch.o_d\[1\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5463_ core_0.execute.alu_mul_div.div_cur\[14\] _1898_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_0_41_266 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_78_53 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7202_ _3385_ _3389_ _0383_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_151_290 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4414_ _0883_ _1018_ _1019_ _0963_ net170 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_4
X_8182_ _0358_ clknet_leaf_125_i_clk core_0.execute.alu_mul_div.mul_res\[8\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_1_352 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5394_ _1233_ _1832_ _1837_ _1838_ _1839_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XANTENNA__7249__A1 _3409_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_100_839 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7133_ _3149_ _3338_ _3339_ net214 _3209_ _3340_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai32_1
X_4345_ _0877_ _0963_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_10_675 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4276_ core_0.fetch.prev_request_pc\[11\] _0854_ _0894_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7064_ _3247_ _3275_ _1229_ _3276_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_214_707 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_105_Left_352 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
X_6015_ _1380_ _2400_ _2404_ _2405_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_241_515 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4483__A1 _1068_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_2_535 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_241_548 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6224__A2 _1117_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_38_965 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_222_784 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4235__A1 _0824_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7966_ _0143_ clknet_leaf_45_i_clk core_0.execute.mem_stage_pc\[1\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_139_508 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_167_839 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_179_699 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6917_ net90 _3135_ _3139_ _3144_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_159_2415 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_159_2426 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_7897_ _0088_ clknet_leaf_70_i_clk core_0.decode.i_imm_pass\[6\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_178_198 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_77_675 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_92_601 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_9_430 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6848_ core_0.execute.rf.reg_outputs\[2\]\[14\] _3085_ _3098_ _3104_ vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_18_720 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_135_714 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_114_Left_361 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_80_807 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_92_667 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5735__A1 _2090_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_17_241 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6779_ _3063_ _3065_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_119_298 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_135_747 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_135_769 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4002__A4 core_0.execute.rf.reg_outputs\[6\]\[8\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_60_531 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_72_391 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_134_279 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output181_I net181 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_115_471 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_255 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3934__I _0567_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_94_1639 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_60_586 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_597 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6160__A1 _2294_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_102_165 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_103_699 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4710__A2 _1253_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_217_523 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_123_Left_370 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_183_2711 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_229_394 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_245_865 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_232_559 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_169_110 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_197_430 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7412__A1 net227 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_200_423 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_68_642 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_184_102 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4777__A2 _1285_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_197_496 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5974__A1 _1596_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_200_445 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_67_152 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_103_1746 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_166_861 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_194_2840 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7715__A2 _1064_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_165_371 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5726__A1 _1124_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_165_393 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_181_842 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_317 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_177 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_153_544 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_70_328 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_723 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_36_594 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_180_352 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_113_419 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xrebuffer4 net223 net224 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_180_374 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_58_1203 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_153_599 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_58_1214 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_11_406 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_51_575 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_586 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_11_428 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_51_597 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6151__A1 net84 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6151__B2 _2537_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_48_34 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_114_1875 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_139_58 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_114_1886 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_4130_ core_0.execute.prev_pc_high\[4\] _0743_ _0749_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_225_3217 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_48_89 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_236_865 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_219_80 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4061_ _0533_ _0524_ _0526_ core_0.execute.rf.reg_outputs\[6\]\[3\] _0685_ vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_4
XANTENNA__5257__A3 _1525_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7651__A1 _1132_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_223_537 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_64_33 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_143_2227 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_223_559 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_161_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_69_1343 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_78_406 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_207_2994 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_64_77 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7403__A1 core_0.execute.sreg_irq_pc.o_d\[3\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_210_209 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7820_ core_0.dec_pc_inc _1032_ _3831_ _1216_ _3878_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai211_1
XTAP_TAPCELL_ROW_35_935 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_7751_ _3663_ _3828_ _0493_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_176_636 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4768__A2 _1285_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4963_ core_0.execute.sreg_priv_control.o_d\[10\] _1394_ _1417_ _1391_ _1418_ vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_59_664 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_86_461 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_86_472 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6702_ core_0.ew_reg_ie\[5\] _2934_ _3020_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_0_191_606 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3914_ _0539_ core_0.execute.rf.reg_outputs\[3\]\[15\] _0549_ _0550_ vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_2
XTAP_TAPCELL_ROW_236_3346 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_7682_ _1037_ _1082_ _3780_ _3781_ _3782_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_171_78 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4894_ _1321_ _1360_ _1361_ _0103_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_191_628 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_129_574 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__7706__A2 _1053_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_62_807 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6633_ _2929_ _2974_ _2975_ _2976_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_0_104_72 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_550 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_156_382 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_172_831 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3991__A3 net231 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_15_692 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_73_166 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6390__A1 _2287_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_89_30 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6564_ core_0.dec_rf_ie\[2\] core_0.ew_reg_ie\[2\] _1985_ _2923_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_154_2356 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_171_352 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_380 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6390__B2 _1690_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_144_577 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_531 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_54_391 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_8303_ _0479_ clknet_leaf_76_i_clk net188 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_4
XFILLER_0_14_244 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_89_63 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5515_ _1063_ _1946_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_171_396 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6495_ _2872_ _2180_ _2873_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__4940__A2 _1394_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_14_266 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8234_ _0410_ clknet_leaf_34_i_clk core_0.execute.sreg_irq_pc.o_d\[6\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_42_597 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_737 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6142__A1 core_0.ew_data\[5\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5446_ core_0.execute.alu_mul_div.div_cur\[10\] _1814_ _1817_ _1883_ _1884_ vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_66_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_2_683 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6693__A2 _3006_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_8165_ _0341_ clknet_leaf_89_i_clk net102 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_4
X_5377_ _1748_ _1813_ _1824_ _0123_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_1
XANTENNA_clkbuf_leaf_92_i_clk_I clknet_4_6__leaf_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7116_ _1364_ _3322_ _3323_ _1367_ _3324_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai211_2
X_4328_ _0934_ _0942_ _0945_ _0946_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_4
X_8096_ _0272_ clknet_leaf_94_i_clk core_0.execute.rf.reg_outputs\[4\]\[3\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_input38_I i_req_data[0] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_129_80 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7642__A1 _0745_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6445__A2 _2279_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_242_813 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7047_ _1224_ _1909_ core_0.execute.alu_mul_div.cbit\[1\] _3260_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_2
X_4259_ core_0.fetch.pc_flush_override _0876_ _0877_ _0878_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_165_2496 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_198_249 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_179_430 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_201_209 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_69_428 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4208__A1 _0723_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_210_732 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_96_247 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7949_ _0127_ clknet_leaf_3_i_clk core_0.execute.alu_mul_div.div_cur\[5\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_2
XANTENNA__4759__A2 _1279_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3929__I _0563_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5956__B2 core_0.execute.alu_flag_reg.o_d\[2\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_65_623 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_64_111 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_42_1015 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_166_179 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_65_667 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_107_202 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_147_382 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_282 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_107_224 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_163_842 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_52_317 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_64_177 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_135_566 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5184__A2 _1604_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_135_577 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6381__A1 _2242_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_107_279 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4931__A2 _0731_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7136__I core_0.execute.alu_mul_div.mul_res\[15\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6133__A1 _2295_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_60_383 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_131_772 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_20_247 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_103_485 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6684__A2 _2999_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_130_293 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_53_1144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_218_865 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7633__A1 _3732_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_18_37 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6436__A2 _1702_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_233_813 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_129_2060 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_244_161 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8011__CLK clknet_leaf_53_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4447__A1 _1038_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_232_312 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_189_227 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4998__A2 _1444_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_220_3147 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_88_737 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_220_3158 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_198_772 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_197_271 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_197_282 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_185_422 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__8161__CLK clknet_leaf_88_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5947__A1 _2335_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_158_647 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_56_623 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_185_466 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_138_360 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_44_807 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_28_358 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_64_1284 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7755__B _1032_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_144 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_126_522 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_464 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_138_382 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_615 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_153_341 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_154_864 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_12_651 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_12_662 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_55_199 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_153_352 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_71_659 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_40_993 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_116_1904 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7879__CLK clknet_leaf_83_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_180_171 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_231_3287 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_180_Right_180 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_3_458 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_59_22 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5300_ _1747_ _1748_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA__6124__A1 _1061_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_114_i_clk_I clknet_4_4__leaf_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6280_ _2624_ _2661_ _2662_ _2664_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_1
XANTENNA__6124__B2 _1109_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_219_Left_466 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_59_66 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7490__B _1284_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_88 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5231_ _1601_ _1679_ _1680_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6675__A2 _2999_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_209_821 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4686__A1 net49 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5162_ _0776_ _1607_ _1609_ _1610_ _1611_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai211_4
XFILLER_0_208_331 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_166_34 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_209_865 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_224_813 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7624__A1 core_0.execute.pc_high_buff_out\[1\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4113_ core_0.execute.pc_high_out\[3\] _0732_ _0733_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_4
X_5093_ _1531_ _1541_ _1542_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4438__A1 _0721_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_236_695 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_76 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_75_87 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4044_ net99 _0578_ _0670_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_79_704 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclone9 _0547_ net231 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dlya_2
XFILLER_0_189_772 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_182_55 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_228_Left_475 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_78_247 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7803_ core_0.decode.i_instr_l\[13\] _3788_ _3866_ core_0.decode.i_instr_l\[10\]
+ _1133_ _3867_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_0_149_625 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_149_636 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4354__B _0970_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_188_282 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5938__A1 _2281_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_176_422 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5995_ core_0.execute.alu_mul_div.mul_res\[2\] _2386_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_0_93_206 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_39_i_clk_I clknet_4_11__leaf_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6060__B1 _2257_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_93_228 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_59_483 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7734_ _3818_ _0486_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4946_ _1195_ net205 _1406_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_19_325 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_122 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_117_500 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_157_680 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7665_ _1066_ _1069_ _3769_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_4877_ _0830_ _1321_ _1352_ _0095_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_145_842 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_163_138 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_317 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_46_177 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_6_241 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6616_ _2935_ _2962_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XANTENNA__6363__A1 _2411_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_172_661 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7596_ _3663_ _3714_ _0452_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_6547_ _2914_ _0203_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XPHY_EDGE_ROW_237_Left_484 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_132_569 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6478_ _1088_ _2854_ _2856_ _2332_ _2857_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai211_4
XFILLER_0_113_772 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_91_1609 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_8217_ _0393_ clknet_leaf_36_i_clk net74 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_4
XFILLER_0_30_567 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5429_ _1232_ _1868_ _1869_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_30_589 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_167_2514 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_246_426 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8148_ _0324_ clknet_leaf_116_i_clk core_0.execute.rf.reg_outputs\[1\]\[7\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_246_459 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7615__A1 _3729_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6418__A2 _2797_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_227_684 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8079_ _0255_ clknet_leaf_117_i_clk core_0.execute.rf.reg_outputs\[5\]\[2\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_226_161 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_226_37 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__7091__A2 _3285_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_241_142 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_246_Left_493 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_69_203 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_230_849 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5929__A1 _1819_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_167_422 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_179_282 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_210_551 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_38_601 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6051__B1 _2440_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_194_230 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_84_217 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_178_2643 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_178_2654 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_182_403 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_100_1716 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_37_133 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_108_500 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_38_667 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_37_144 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_26_807 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_182_425 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_191_2810 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_154_127 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_615 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3955__A3 _0536_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_92_261 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_25_317 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5157__A2 _0773_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_111_18 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_135_352 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_151_812 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_18_391 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_52_136 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_599 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_150_300 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4904__A2 _1221_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6106__A1 _1378_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_61_692 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_104_761 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_21_556 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6919__B _3139_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4117__B1 _0736_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6657__A2 _2992_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_103_282 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_209_117 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_189_2783 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_111_1845 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_206_802 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7606__A1 core_0.execute.pc_high_out\[6\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6409__A2 _2531_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_224_109 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_217_150 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_245_481 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_233_621 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_245_492 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_233_632 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7082__A2 _3177_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_136_37 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_232_131 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_205_345 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5093__A1 _1531_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_66_1302 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_177_208 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_204_2964 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_88_545 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4840__A1 core_0.decode.i_instr_l\[14\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4691__I1 net63 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_17_721 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_76_729 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_40_i_clk_I clknet_4_11__leaf_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_201_562 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_61_34 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_75_228 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4800_ _1169_ _1305_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_185_252 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6593__A1 _2936_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5780_ _1107_ _1989_ _2181_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_118_308 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_122_1974 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_158_488 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_61_78 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_233_3305 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_4731_ _0855_ _1238_ _1266_ _0035_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_127_842 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_56_475 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_124_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_28_177 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_317 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7450_ _3581_ _3605_ _0415_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_43_114 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6345__A1 _2576_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4662_ _1209_ core_0.execute.sreg_priv_control.o_d\[0\] _0810_ _1219_ vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_0_44_659 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_126_363 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_71_456 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_153_160 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_158 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6401_ _2279_ _2780_ _2781_ _2782_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_2
XANTENNA__6896__A2 _3129_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_141_322 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7381_ core_0.execute.mem_stage_pc\[0\] _3548_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_151_2326 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_4593_ _1161_ net140 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__8057__CLK clknet_leaf_99_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_372 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_12_512 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_77_1431 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_77_1442 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6332_ _2714_ _1114_ _1117_ _2715_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_3_277 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_545 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_180 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_865 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6829__B _3083_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6648__A2 _2986_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6263_ core_0.execute.alu_mul_div.mul_res\[8\] _2648_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__inv_3
XFILLER_0_122_591 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8002_ _0179_ clknet_leaf_48_i_clk core_0.ew_data\[1\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_2
X_5214_ _1659_ _1660_ _1661_ _1662_ _1663_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_0_86_53 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6194_ core_0.execute.sreg_priv_control.o_d\[7\] _1386_ _2579_ core_0.execute.sreg_scratch.o_d\[7\]
+ _2580_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__5320__A2 _1557_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_244_3445 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_243_407 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_215_109 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5145_ _1482_ _1585_ _1593_ _1531_ _1594_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai211_2
XTAP_TAPCELL_ROW_149_2299 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_223_131 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5076_ _1521_ _1522_ _1523_ _1524_ _1525_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_4
XTAP_TAPCELL_ROW_162_2455 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_29_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4027_ _0516_ core_0.execute.rf.reg_outputs\[3\]\[6\] net231 _0654_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_2
XANTENNA__6820__A2 _3087_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_168_208 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_88_1571 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_211_337 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_149_422 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_94_515 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_177_742 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_217 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_176_241 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_177_764 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_149_466 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_192_712 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5978_ _1559_ _1555_ _2300_ _2369_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_94_559 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_176_263 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7781__B1 _3827_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_192_734 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_192_745 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_75_762 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7717_ core_0.decode.i_imm_pass\[3\] _1064_ _3810_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__7395__B _3546_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_81_209 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4929_ _1392_ _1390_ _1393_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_0_191_233 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3937__A3 _0544_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_47_486 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_75_795 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_7648_ core_0.execute.pc_high_buff_out\[7\] _3732_ _3756_ _3757_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__5627__C _2014_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_117_352 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6336__B2 net2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7533__B1 _1398_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_90_776 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_132_311 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_173_2584 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6887__A2 _3108_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7579_ net203 _3675_ _3699_ _3700_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__4898__A1 _1364_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4103__I core_0.fetch.out_buffer_valid vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_120_506 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_132_399 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6639__A2 core_0.ew_data\[8\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3942__I net92 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_30_375 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_101_753 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_246_234 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5311__A2 _1758_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4259__B _0877_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_50_1114 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_227_492 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_215_632 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_126_2030 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_214_131 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5075__A1 net93 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_242_451 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_215_687 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_199_366 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6811__A2 _3065_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_203_838 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_18 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_159_208 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_98_865 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_15_38 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_57_206 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_729 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_97_375 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_48_1087 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5378__A2 _1811_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_167_263 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4425__I1 _0851_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_431 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7772__B1 _3833_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_127_116 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_109_842 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_61_1243 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_93_570 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_65_272 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_509 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_341 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6327__A1 _2090_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_26_648 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5537__C _1950_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_182_277 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_445 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6878__A2 _3108_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_53_489 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4889__A1 _1357_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_123_344 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5550__A2 _1956_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_111_528 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_150_163 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_865 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_21_342 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5553__B _1964_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_237_212 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7917__CLK clknet_4_3__leaf_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5302__A2 _1711_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_56_34 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_72_1372 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_56_45 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_205_142 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5066__A1 _1466_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4683__I _1236_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6802__A2 _3070_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6950_ _3166_ _3169_ _3170_ _1225_ _1223_ _3171_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai221_4
XFILLER_0_220_101 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_221_646 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5901_ net223 _2112_ _2293_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_2
XANTENNA__5081__A4 _1529_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_159_731 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_241_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_88_364 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6881_ core_0.execute.rf.reg_outputs\[1\]\[12\] _3114_ _3112_ _3123_ vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_163_68 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_88_375 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_48_228 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_76_548 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5832_ _2226_ _2227_ _2228_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_220_189 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_3_0_0_i_clk_I clknet_0_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_146_403 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_159_786 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_8_325 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_173_222 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_17_604 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5763_ _1756_ _1592_ _2164_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_17_615 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_118_149 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_486 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_134_609 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_581 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7502_ _3514_ _3640_ _3644_ _0428_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_56_283 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4714_ _1255_ _1237_ _1256_ _0028_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_56_294 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6318__A1 _2286_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5694_ _1123_ _1620_ _2091_ _2092_ _2095_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai211_2
XANTENNA__6318__B2 _1455_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_20_749 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_114_311 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7433_ core_0.execute.mem_stage_pc\[9\] _3591_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__6869__A2 _3114_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_4_520 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_253 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4645_ _1195_ _1203_ _1204_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_25_670 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_130_804 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_142_664 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_102_506 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7364_ _2384_ _2434_ _3532_ _3533_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor3_1
X_4576_ core_0.ew_data\[2\] net157 _1153_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__5541__A2 _1956_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_4_597 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_342 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_188_76 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6315_ _2045_ _2050_ _2698_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_7295_ _3409_ _3471_ _3472_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_188_98 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_40_695 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7294__A2 _3393_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6246_ _1121_ _2630_ _2631_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6177_ _2549_ _2551_ _2563_ _2564_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_244_749 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_54_i_clk clknet_4_11__leaf_i_clk clknet_leaf_54_i_clk vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_209_492 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5128_ _1482_ _1576_ _1577_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_input20_I i_mem_ack vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_224_440 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5057__A1 _0619_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6294__B core_0.decode.oc_alu_mode\[7\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_137_80 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_224_473 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5059_ _1466_ _0608_ _0613_ _0614_ _1508_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_0_79_331 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4804__A1 _0816_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_28_849 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_39_206 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4280__A2 _0830_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_69_i_clk clknet_4_15__leaf_i_clk clknet_leaf_69_i_clk vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__6006__B1 _2250_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_0_496 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_175_2613 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_165_745 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6309__A1 core_0.ew_data\[9\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_109_Right_109 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_118_661 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_192_586 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_180_737 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_117_171 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_35_478 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_629 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_121_804 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_50_448 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_160_461 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_120_314 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_132_174 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6580__I1 core_0.ew_mem_width vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_8_i_clk_I clknet_4_3__leaf_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7809__A1 _1038_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_30_150 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_186_2742 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4638__A4 net190 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5048__A1 _0789_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_26_37 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_188_815 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_187_303 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5599__A2 _1641_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_202_123 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_86_802 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_201_2923 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_97_150 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_230_498 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6548__A1 net131 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_106_1788 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_217_3119 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_197_2871 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_197_2882 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_168_594 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_38_261 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4023__A2 _0529_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5220__A1 _0771_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_155_244 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_6_807 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_26_423 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_155_266 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_672 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_115_108 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_170_203 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_183_586 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_26_445 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5771__A2 _1568_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_135_2129 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_14_607 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_562 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_108_171 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_54_798 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_170_247 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_297 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_112_804 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4430_ _0735_ net110 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_13_139 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7482__C _1950_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_2 net101 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_651 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_74_1401 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_4361_ _0972_ _0966_ _0976_ _0963_ net165 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XFILLER_0_21_150 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1_556 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_238_521 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6100_ core_0.execute.sreg_priv_control.o_d\[5\] _1385_ _2257_ core_0.execute.pc_high_out\[5\]
+ _2448_ _2488_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_0_1_578 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_228_3248 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_7080_ _3149_ _3290_ _3291_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_4292_ core_0.fetch.prev_request_pc\[3\] _0857_ _0910_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_191_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_226_727 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_225_204 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6031_ _2009_ _2421_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_67_88 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_241_3404 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_146_2269 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_174_34 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5039__A1 _0789_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_169_Left_416 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
X_7982_ _0159_ clknet_leaf_28_i_clk core_0.execute.prev_pc_high\[1\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__6787__A1 _2956_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_83_76 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_178_314 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4346__C _0963_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_83_87 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_89_651 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6933_ core_0.execute.alu_mul_div.cbit\[3\] core_0.execute.alu_mul_div.cbit\[2\]
+ _3152_ _3153_ _3154_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor4_4
XTAP_TAPCELL_ROW_85_1530 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_107_72 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_194_807 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6842__B _3098_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_89_684 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_25_808 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_88_172 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6864_ _3106_ _3114_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_119_403 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_239_3377 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_193_339 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_146_211 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_147_734 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_36_209 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_111 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5815_ _2211_ _2212_ _2213_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__7200__A2 _0709_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6795_ _2972_ _3064_ _3074_ _0291_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__4014__A2 _0523_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5211__A1 _0782_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_146_244 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_91_337 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_91_348 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5746_ _1997_ _2147_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_45_754 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_8_177 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_106_119 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_162_737 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_91 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_96_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_174_597 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_45_776 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_146_299 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_157_2398 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_72_562 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_161_247 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_EDGE_ROW_178_Left_425 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
X_5677_ _2062_ _2066_ _2071_ _2077_ _2078_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XFILLER_0_142_450 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_161_269 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7416_ _3547_ _3576_ _3577_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_130_601 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_170_2554 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_4628_ _1176_ core_0.execute.alu_flag_reg.o_d\[0\] core_0.execute.alu_flag_reg.o_d\[1\]
+ _1187_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XANTENNA__5514__A2 _1945_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_114_174 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_130_623 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6562__I1 core_0.ew_reg_ie\[1\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_96_1670 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_102_325 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input68_I i_req_data[8] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7347_ _3510_ _3515_ _3517_ _0400_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_13_684 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4559_ _1049_ _1139_ _1140_ _1141_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_130_667 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8000__D _0177_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7267__A2 _3391_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7278_ _1400_ core_0.execute.sreg_irq_pc.o_d\[10\] _1417_ _1430_ _3457_ vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_6229_ core_0.ew_data\[7\] _2486_ _2615_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_110_391 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_218_49 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7019__A2 _3181_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_187_Left_434 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_5_577 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_99_415 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_181_2683 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_234_37 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_86_109 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6242__A3 _1721_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_150 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_169_347 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6752__B _3045_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5450__A1 _1374_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_197_678 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_95_632 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_184_317 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_196_177 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_137_200 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_138_734 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5368__B core_0.execute.alu_mul_div.comp vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_87_i_clk_I clknet_4_12__leaf_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_138_745 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_177_380 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_45_1057 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_55_529 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_389 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_83_838 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_193_862 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4005__A2 _0535_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5202__A1 net95 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_137_266 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_196_Left_443 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_125_428 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_180_523 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6950__B2 _1225_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_51_702 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_63_562 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_152_247 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_223 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_121_601 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_51_768 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6702__A1 core_0.ew_reg_ie\[5\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_133_472 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_174 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_106_697 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_105_185 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4498__I _1063_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50_278 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_31_470 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7258__A2 net85 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5269__A1 core_0.decode.oc_alu_mode\[12\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_120_199 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xoutput72 net72 dbg_pc[0] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XTAP_TAPCELL_ROW_56_1186 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
Xoutput83 net83 dbg_pc[5] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
Xoutput94 net94 dbg_r0[15] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_235_546 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_128_49 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_108_1806 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4492__A2 _1084_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_199_2900 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_188_612 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_223_3189 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_231_741 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_144_37 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__7430__A2 _3544_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_203_454 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_230_251 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_86_610 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_98_470 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6662__B _2984_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_176_807 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_203_476 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_312 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_68 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_187_166 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3930_ core_0.execute.rf.reg_outputs\[2\]\[13\] _0564_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_230_284 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_141_2199 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5992__A2 _1456_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_85_142 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_378 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_86_687 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_175 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_129_767 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7194__A1 net79 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5600_ _1676_ _2001_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_128_255 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_348 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_116_406 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_80_1471 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6580_ core_0.dec_mem_width core_0.ew_mem_width _2201_ _2932_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__6941__A1 _1231_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_143_214 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_144_737 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_171_523 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_551 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6941__B2 _1926_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_54_562 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5531_ _1024_ _1956_ _1958_ _0143_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__7493__B _1395_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_5_136 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_119_1935 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_204_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_119_1946 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_41_212 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_30_877 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_124_450 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8250_ _0426_ clknet_leaf_23_i_clk core_0.execute.sreg_scratch.o_d\[0\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5462_ _1798_ _1817_ _1897_ _1748_ _0135_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_124_472 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7497__A2 _3641_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6544__I1 _2652_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_200_Left_447 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_111_100 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7741__I0 net184 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7201_ _1414_ core_0.execute.sreg_irq_pc.o_d\[1\] _3387_ _3388_ _1736_ _3389_ vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_4413_ net81 _0883_ _1019_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_111_122 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_8181_ _0357_ clknet_leaf_126_i_clk core_0.execute.alu_mul_div.mul_res\[7\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_2_865 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_100_807 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5393_ _1809_ _1838_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_112_667 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7132_ _3336_ _3331_ _3337_ _3339_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_4344_ net78 _0883_ _0962_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_7063_ _1909_ _1592_ _3274_ _3275_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_4275_ _0892_ _0837_ _0844_ _0890_ _0893_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__7512__I _0722_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_226_557 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6014_ _1380_ core_0.execute.sreg_irq_pc.o_d\[3\] _2404_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_185_66 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4357__B _0945_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_185_99 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_213_218 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_118_82 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_2_536 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_206_292 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_178_111 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_178_122 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_221_240 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_11_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_38_966 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_7965_ _0142_ clknet_leaf_13_i_clk core_0.execute.mem_stage_pc\[0\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__4235__A2 net57 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_109_i_clk_I clknet_4_5__leaf_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5432__A1 _1747_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_77_632 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_167_829 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_178_155 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_334 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_166_306 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_76_120 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6916_ _2986_ _3130_ _3143_ _0343_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_159_2416 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_194_637 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_193_114 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_49_356 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7896_ _0087_ clknet_leaf_72_i_clk core_0.decode.i_imm_pass\[5\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_76_153 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_194_Right_194 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_147_542 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6847_ _2992_ _3087_ _3103_ _0314_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__7185__A1 _1748_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_64_326 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_92_635 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_18_732 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5196__B1 _1436_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_107_417 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6932__A1 _1362_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5196__C2 _1443_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6778_ _3063_ _3064_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_91_167 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_134_225 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_562 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_17_253 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_190_865 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5729_ _1549_ _2091_ _2130_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_17_264 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_134_247 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_17_286 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_72_381 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_115_483 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5499__A1 _1908_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_102_111 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output174_I net174 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_103_656 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_142_291 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_492 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4171__A1 core_0.ew_reg_ie\[4\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_245_800 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6747__B _3045_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6448__B1 _2577_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_183_2712 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_244_321 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_205_708 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_99_212 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_244_387 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_232_527 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5671__A1 _1528_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_213_730 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_99_267 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87_418 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7412__A2 _3544_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_158_807 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5423__A1 core_0.execute.alu_mul_div.div_cur\[7\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_157_306 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_240_593 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_142 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_157_339 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_95_462 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_103_1747 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7176__A1 _1223_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_161_Right_161 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_194_2841 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5726__A2 _1541_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_83_679 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6923__A1 net93 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_126_737 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_138_597 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_181_832 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_126_759 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_153_556 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_181_865 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_23_212 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xrebuffer5 _0879_ net225 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_3_618 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_58_1204 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_140_228 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7723__I0 net190 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_23_267 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_239_126 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6151__A2 _2531_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4021__I net216 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_121_475 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_114_1876 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5561__B _1964_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6439__B1 _2516_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_225_3207 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_225_3218 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_208_524 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7100__A1 _1230_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_236_855 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4060_ _0567_ core_0.execute.rf.reg_outputs\[3\]\[3\] net226 _0684_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_0_223_505 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_143_2228 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_207_2995 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_69_1344 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7403__A2 _3543_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_204_774 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_89 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_110_i_clk_I clknet_4_5__leaf_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5414__A1 core_0.execute.alu_mul_div.div_cur\[7\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_154_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_59_632 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_82_1500 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_4962_ _1381_ _0615_ _1417_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_35_936 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_7750_ core_0.dec_jump_cond_code\[2\] _3766_ _1070_ _3827_ _3828_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_148_317 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5965__A2 core_0.dec_sreg_jal_over vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_86_451 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_176_648 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_33 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3913_ _0548_ _0549_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_8
XANTENNA__3976__A1 _0565_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_74_613 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6701_ _2996_ _3000_ _3019_ _0252_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_175_136 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7681_ _1066_ _1056_ _1048_ _1046_ _3781_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XANTENNA__7167__A1 _3357_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_73_101 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4893_ core_0.decode.i_jmp_pred_pass _1305_ _1361_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_157_862 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_236_3347 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_74_635 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6632_ net34 _1149_ _2975_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5178__B1 _1434_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6914__A1 _2983_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_15_693 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_15_702 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_13_82 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_172_843 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_73_178 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_116_247 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6563_ _2922_ _0211_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_172_865 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_154_2357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_8302_ _0478_ clknet_leaf_12_i_clk net187 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_4
XFILLER_0_144_589 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5514_ _1419_ _1945_ _0139_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_14_234 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_70_863 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6494_ _1988_ _1989_ _2872_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_131_228 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_42_565 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8233_ _0409_ clknet_leaf_42_i_clk core_0.execute.sreg_irq_pc.o_d\[5\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_14_278 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_120_83 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5445_ _1881_ _1882_ _1838_ _1883_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__6142__A2 _2486_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4153__A1 _0768_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_246_608 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_35_i_clk_I clknet_4_11__leaf_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_196_43 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8164_ _0340_ clknet_leaf_88_i_clk net101 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_4
X_5376_ core_0.execute.alu_mul_div.div_cur\[0\] _1814_ _1817_ _1823_ _1824_ vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_59_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_1_194 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7115_ _1364_ _3295_ _3323_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4327_ _0877_ _0944_ _0871_ _0941_ _0945_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or4_4
X_8095_ _0271_ clknet_leaf_110_i_clk core_0.execute.rf.reg_outputs\[4\]\[2\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_7046_ _3243_ _3252_ _3258_ _3259_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XANTENNA__7642__A2 _3729_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4258_ core_0.fetch.pc_reset_override _0877_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XANTENNA__5653__A1 _1789_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_226_387 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_214_527 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_199_729 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_165_2497 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_4189_ core_0.execute.alu_mul_div.comp _0804_ _0807_ _0808_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__nor3_4
XANTENNA__5405__A1 _1747_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_194_401 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_222_593 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_120 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_167_626 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7948_ _0126_ clknet_leaf_3_i_clk core_0.execute.alu_mul_div.div_cur\[4\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5956__A2 _2264_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4759__A3 _0813_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3967__A1 _0517_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7879_ _0070_ clknet_leaf_83_i_clk core_0.decode.i_instr_l\[4\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_2
XANTENNA__4106__I _0725_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_42_1016 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_64_134 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_64_145 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_92_454 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6905__A1 _2967_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_181_128 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_65_679 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_135_534 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_147_394 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_190_640 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6381__A2 _0604_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output99_I net99 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_598 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6133__A2 _2501_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5192__I0 net186 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4144__B2 core_0.ew_reg_ie\[1\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_236_107 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_0_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_53_1145 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_217_332 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7950__CLK clknet_leaf_4_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_245_674 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_129_2061 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_245_696 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_230_Right_230 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__5644__A1 _2026_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4447__A2 _1039_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_233_858 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_220_3148 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_16_Right_16 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_87_226 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8306__CLK clknet_leaf_76_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_37 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_87_237 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_201_722 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_198_784 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4217__S _0723_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_197_261 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_157_103 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_205_50 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_197_294 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_201_766 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_613 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_68_473 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_7_209 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_64_1285 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7755__C _1084_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_56_679 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_172_139 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_70_104 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_71_627 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_329 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_638 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6372__A2 _1386_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_12_652 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_71_649 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_113_206 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4383__A1 _0844_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_40_994 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_25_Right_25 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_52_863 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_116_1905 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_231_3288 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6124__A2 _1693_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_51_384 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_226 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_122_773 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5230_ _1643_ _1654_ _1624_ _1678_ _1679_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__4135__A1 _0731_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4686__A2 _1238_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5883__A1 _2242_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_227_129 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5161_ core_0.execute.rf.reg_outputs\[4\]\[6\] _1436_ _1437_ core_0.execute.rf.reg_outputs\[2\]\[6\]
+ _1610_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_0_209_855 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4112_ net105 _0732_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XANTENNA__7624__A2 _3732_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_166_57 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5092_ net214 _1541_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__inv_2
XFILLER_0_224_836 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5635__A1 _1754_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4438__A2 _1032_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_208_387 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_223_324 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4043_ _0665_ _0666_ _0667_ _0668_ _0669_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and4_1
XPHY_EDGE_ROW_34_Right_34 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_75_99 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_223_346 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_78_204 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_142_Left_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_182_34 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_79_749 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_195_209 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_91_43 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_149_615 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7802_ _3837_ _3859_ _3863_ _3865_ _3866_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_4
X_5994_ _2281_ _2384_ _2385_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_91_76 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6060__A1 core_0.execute.pc_high_buff_out\[4\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_451 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_115_50 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_176_434 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3949__A1 _0534_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_115_72 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4945_ _1301_ _1405_ _0110_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_7733_ net180 core_0.decode.i_imm_pass\[11\] _1946_ _3818_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_86_270 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6850__B _3098_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_74_421 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_136_309 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_74_432 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_176_489 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_46_134 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4876_ core_0.decode.i_imm_pass\[13\] _1341_ _1352_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_46_145 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_74_454 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7664_ _3663_ _3768_ _0466_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_62_605 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_465 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_34_307 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_74_487 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_117_545 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6615_ _2930_ core_0.ew_data\[4\] _2960_ _2961_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_4
XFILLER_0_34_329 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_638 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7595_ core_0.execute.pc_high_out\[5\] _3673_ _3713_ _3714_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__oai21_1
XPHY_EDGE_ROW_43_Right_43 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__7560__A1 core_0.execute.pc_high_out\[1\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6363__A2 _2642_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_144_364 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_61_148 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6546_ net130 _2690_ _2906_ _2914_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__5185__C net219 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_151_Left_398 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_6_297 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7681__B _1048_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_30_513 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7312__A1 _1395_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6477_ _1433_ _2855_ _2856_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_113_762 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4126__A1 core_0.execute.pc_high_out\[6\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_112_261 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8216_ _0392_ clknet_leaf_35_i_clk net73 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_4
X_5428_ _1867_ _1785_ _1868_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA_input50_I i_req_data[20] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_218_107 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_140_592 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_167_2515 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_218_129 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8147_ _0323_ clknet_leaf_116_i_clk core_0.execute.rf.reg_outputs\[1\]\[6\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5359_ _1751_ _1805_ _1806_ _1807_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_8078_ _0254_ clknet_leaf_117_i_clk core_0.execute.rf.reg_outputs\[5\]\[1\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_2
XPHY_EDGE_ROW_52_Right_52 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_199_504 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5626__A1 _2010_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_226_173 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_214_313 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7029_ _3237_ _3241_ _3242_ _3243_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA_output137_I net137 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_199_559 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_242_677 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_186_209 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_97_546 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_195_710 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_241_198 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_195_721 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_69_259 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_167_412 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_85_719 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5929__A2 _1665_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_139_125 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_167_434 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6051__A1 _2403_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_242_37 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6051__B2 _2360_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_195_765 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_178_2644 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6760__B _3045_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_37_123 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_194_275 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_657 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_100_1717 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_155_629 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_93_752 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_191_2800 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_148_681 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_61_Right_61 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_147_180 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_154_139 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_627 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5376__B _1817_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_52_104 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_136_865 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_135_342 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_457 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_863 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_150_312 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_479 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_33_384 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_60_170 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_103_272 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_237_416 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_29_26 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_189_2784 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5865__A1 _1382_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_70_Right_70 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_111_1846 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7606__A2 core_0.execute.pc_high_out\[5\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_205_302 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6935__B _1230_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_205_313 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_205_324 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5093__A2 _1541_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_205_368 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_221_828 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_66_1303 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_204_2965 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4840__A2 _1307_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_17_711 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_186_721 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_17_722 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_88_568 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_216_93 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_185_220 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_152_37 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_56_410 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7846__CLK clknet_leaf_67_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_29_646 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6593__A2 _2940_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7790__A1 _0536_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_122_1975 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_173_415 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4730_ net48 _1253_ _1266_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_233_3306 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_29_668 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_145_128 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_173_448 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_56_487 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_126_331 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_4661_ _1218_ _0014_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_44_649 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_126 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_142_802 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_154_662 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7542__A1 _3663_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_117_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_4_713 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6400_ core_0.execute.alu_mul_div.div_res\[12\] _1114_ _2781_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7380_ net37 _3547_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
X_4592_ core_0.ew_data\[2\] core_0.ew_data\[10\] _1150_ _1161_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_3_212 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_151_2327 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_181_492 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_52_671 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_114_559 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_153_194 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_77_1432 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6331_ core_0.execute.alu_mul_div.div_res\[10\] _2714_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_0_12_524 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_384 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_101_209 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_40_855 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_12_557 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4108__A1 net37 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5733__C _2133_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6262_ _2281_ _2646_ _2647_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5213_ core_0.execute.rf.reg_outputs\[1\]\[3\] _1615_ _1483_ _1662_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_8001_ _0178_ clknet_leaf_49_i_clk core_0.ew_data\[0\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_228_438 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_177_67 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6193_ _2254_ _2579_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XTAP_TAPCELL_ROW_244_3435 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7721__S _1946_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_244_3446 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_5144_ _1481_ _1592_ _1593_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_243_419 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5075_ net93 _0521_ _0557_ _0562_ _1461_ _1524_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai221_4
XANTENNA__6281__A1 _2356_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_193_66 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5084__A2 _1438_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_162_2456 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_4026_ _0532_ _0523_ _0526_ core_0.execute.rf.reg_outputs\[6\]\[6\] _0653_ vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_4
XTAP_TAPCELL_ROW_88_1572 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_223_187 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_79_546 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_211_349 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_189_592 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_79_579 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_94_527 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_149_456 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5977_ _1457_ _2366_ _2367_ _2368_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_149_489 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_192_724 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_176_275 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_191_212 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_47_454 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7716_ _1196_ _0514_ _3809_ _0477_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4928_ core_0.execute.prev_sys _0730_ _1392_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or2_2
XFILLER_0_136_139 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_191_245 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_145_640 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_118_865 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7647_ net216 _3733_ _3731_ _3755_ _3756_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__6336__A2 _2579_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_191_278 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_562 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_62_435 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4859_ core_0.decode.i_imm_pass\[5\] _1341_ _1343_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_117_364 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7533__B2 core_0.execute.sreg_irq_flags.o_d\[0\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_144_161 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_145_695 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_16_863 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_173_2585 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_7578_ _3675_ _3698_ _3699_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_105_559 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4898__A2 _1221_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_15_384 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6529_ net116 _1985_ _2905_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_120_518 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4320__S _0725_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_30_365 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5847__A1 _2202_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_30_387 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_208_3010 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_246_268 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_50_1115 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_227_482 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_126_2020 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_242_430 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_215_666 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6272__A1 _2576_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5075__A2 _0521_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_215_699 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_202_327 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_98_855 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_199_389 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4822__A2 core_0.fetch.submitable vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_97_365 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_4_i_clk_I clknet_4_2__leaf_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7586__B _3675_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_410 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_183_702 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_195_562 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_38_421 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_48_1088 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_168_798 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4586__A1 core_0.ew_data\[7\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_443 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_454 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_26_605 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4050__A3 net231 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_61_1244 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_183_768 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_413 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_170_407 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7524__A1 _0604_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_81_744 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_124_802 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_766 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_137_2160 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4338__A1 core_0.fetch.prev_request_pc\[13\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_22_780 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_80_265 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_151_632 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_163_492 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_21_310 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7605__I core_0.execute.pc_high_out\[7\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_855 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_21_321 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_151_698 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_398 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_238_769 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_72_1373 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4510__A1 _1098_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_56_68 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_206_655 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_205_132 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5066__A2 net190 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_221_603 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4813__A2 core_0.fetch.submitable vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_72_34 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5900_ _1458_ _2283_ _2291_ _2292_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_221_669 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6880_ _2988_ _3108_ _3122_ _0328_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_159_743 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6015__A1 _1380_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_72_67 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_88_387 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_186_551 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5831_ _2221_ _2220_ _2219_ _2227_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_201_360 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_234_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_201_371 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_119_618 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_146_415 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_158_275 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_118_117 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5762_ _1754_ _2035_ _2163_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_173_212 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_251 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4041__A3 _0548_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_17_627 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_104 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7501_ core_0.execute.sreg_scratch.o_d\[2\] _3641_ _3516_ _3644_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4713_ net41 _1253_ _1256_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_clkbuf_3_4_0_i_clk_I clknet_0_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_44_435 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_17_649 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5693_ _2091_ _2092_ _2093_ _2094_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_2
XANTENNA__6318__A2 _1789_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6949__S0 _1915_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_161_418 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_173_278 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_457 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7432_ _3581_ _3590_ _0412_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_4644_ core_0.dec_sreg_store _1202_ _1203_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_112_73 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_543 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8174__CLK clknet_leaf_129_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_141_142 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4575_ _1152_ net146 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_12_310 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7363_ _3529_ _3530_ _3531_ _3532_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_141_153 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_141_175 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6314_ _2058_ _2695_ _2696_ _2697_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_7294_ _2783_ _3393_ _3470_ _2791_ _3471_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_0_228_213 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_12_387 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_228_224 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6245_ _2628_ _2042_ _2630_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_229_769 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_243_205 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6176_ _2553_ _2554_ _2558_ _2562_ _2563_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_0_41_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5127_ net89 _1492_ _1571_ _1575_ _1576_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai22_4
XANTENNA_clone2_I _0671_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_619 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_98_107 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_224_452 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_2_Right_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__5057__A2 _0624_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6254__A1 _1592_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5058_ _1503_ _1504_ _1505_ _1506_ _1507_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and4_2
XFILLER_0_98_129 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input13_I i_core_int_sreg[6] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_224_485 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_224_496 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4804__A2 _1306_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4009_ _0637_ net208 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_211_135 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_67_505 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6006__A1 core_0.execute.sreg_long_ptr_en vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_376 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_149_231 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_95_858 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_165_702 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_177_562 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_0_497 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_153_80 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_165_713 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_48_752 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_94_357 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_175_2614 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_109_128 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_164_234 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_785 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_413 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_180_705 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_47_284 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_180_716 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6309__A2 _2486_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_35_435 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_62_221 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_124_109 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_63_766 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_133_621 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_619 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_265 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_63_788 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_574 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_145_492 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_214_3080 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_50_438 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_160_451 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_105_367 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_15_181 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7809__A2 _1094_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output81_I net81 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_219_235 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_186_2743 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_101_562 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_83_i_clk_I clknet_4_12__leaf_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6493__A1 _2576_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_101_584 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_219_279 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_228_780 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_234_249 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_227_290 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_117_18 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_215_441 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_117_29 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_199_142 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_242_260 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6796__A2 _3070_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_201_2924 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_202_157 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_58_527 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_98_696 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_97_184 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6548__A2 _1985_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_42_37 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_106_1789 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_197_2872 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_128_415 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4225__S _0824_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_155_212 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5548__C _1950_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_128_448 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_26_402 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_711 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5220__A2 _0773_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_213_72 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__8197__CLK clknet_leaf_129_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_155_278 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_329 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_170_215 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_276 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_151_473 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_74_1402 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_4360_ _0970_ _0973_ _0975_ _0976_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_0_22_663 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_803 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_37 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_67_34 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_158_47 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4291_ core_0.fetch.prev_request_pc\[4\] _0909_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XTAP_TAPCELL_ROW_228_3249 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6484__A1 net77 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6030_ _1456_ _2420_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__inv_1
XANTENNA__6484__B2 _2537_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_219_780 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_input5_I i_core_int_sreg[13] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_241_3405 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_184_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_225_238 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7028__A3 _1939_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_146_2259 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6236__A1 _1379_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_175_Right_175 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
X_7981_ _0158_ clknet_leaf_28_i_clk core_0.execute.prev_pc_high\[0\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__6787__A2 _3064_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_233_282 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6932_ _1362_ _1451_ _3153_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_2
XTAP_TAPCELL_ROW_85_1531 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_89_674 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_25_809 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_16_82 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_77_836 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_89_696 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_193_307 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_538 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_190_34 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6863_ _2956_ _3107_ _3113_ _0320_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_77_858 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_147_702 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_159_562 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_119_415 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_239_3378 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_190_67 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_9_624 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_119_426 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_190_78 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5814_ _2205_ _2206_ _2183_ _2196_ _2212_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_0_147_746 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6794_ core_0.execute.rf.reg_outputs\[3\]\[6\] _3070_ _3072_ _3074_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_29_251 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_92_839 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_45_711 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4014__A3 _0526_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5211__A2 _0768_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_121_i_clk clknet_4_3__leaf_i_clk clknet_leaf_121_i_clk vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_45_722 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_582 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_8_156 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_123_72 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_45_744 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5745_ _2002_ _2144_ _2145_ _2146_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_0_44_221 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_32_81 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_167 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_162_727 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_45_766 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_44_254 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_157_2399 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_115_632 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_127_492 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4970__A1 core_0.execute.sreg_priv_control.o_d\[12\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
X_5676_ _2076_ _2077_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__4970__B2 _1390_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_44_287 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_89_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7415_ core_0.execute.mem_stage_pc\[6\] _3576_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__4869__I _0837_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_4_340 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_115_665 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_449 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4627_ core_0.dec_jump_cond_code\[1\] _1176_ _1186_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_2
XTAP_TAPCELL_ROW_170_2555 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_130_613 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_142_473 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6711__A2 _3022_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_96_1660 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5193__C net223 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_105_i_clk_I clknet_4_5__leaf_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4722__A1 net44 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_229_500 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4558_ _1041_ _1066_ _1048_ _1140_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_4
X_7346_ core_0.execute.alu_flag_reg.o_d\[2\] _3510_ _3516_ _3517_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_40_482 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_12_173 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7277_ net73 _3398_ _3399_ _3455_ _3456_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_4489_ _1041_ _1056_ _1082_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_244_503 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_110_381 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6228_ _2242_ _2612_ _2613_ _2614_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_6159_ _2293_ _2381_ _2546_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_244_569 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_209_290 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_5_567 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6227__A1 _2242_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_5_578 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_225_772 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_EDGE_ROW_142_Right_142 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_225_794 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_224_282 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_181_2684 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_224_293 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4789__A1 core_0.fetch.prev_request_pc\[12\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_212_444 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4789__B2 net164 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_196_123 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_169_337 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_240_775 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_79_162 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_95_611 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_67_357 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_55_508 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_137_212 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_45_1047 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_55_519 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5368__C _0801_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_45_1058 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4005__A3 _0527_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5202__A2 _1446_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_137_278 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_192_384 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_35_243 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_552 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_777 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4961__A1 _1301_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_90_371 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_133_440 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_142 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6702__A2 _2934_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_133_484 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4713__A1 net41 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_208_706 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6466__A1 _1059_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput73 net73 dbg_pc[10] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XTAP_TAPCELL_ROW_56_1187 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
Xoutput84 net84 dbg_pc[6] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
Xoutput95 net95 dbg_r0[1] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_207_216 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_207_227 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_235_558 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_222_208 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_108_1807 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_203_422 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_199_2901 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6769__A2 _3049_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_53_14 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_230_241 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5559__B _1964_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_203_488 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_858 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_129_702 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_224_82 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_74_839 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7194__A2 _1739_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_184_863 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_582 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_160_37 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_39_593 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_221 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_80_1472 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_27_766 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6941__A2 _1758_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4952__A1 _1400_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5530_ core_0.execute.mem_stage_pc\[1\] _1957_ _1217_ _1958_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xclkbuf_leaf_53_i_clk clknet_4_14__leaf_i_clk clknet_leaf_53_i_clk vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_TAPCELL_ROW_30_867 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_26_276 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_119_1936 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_171_557 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_30_878 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_81_382 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5294__B _1735_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_4_11__f_i_clk clknet_3_5_0_i_clk clknet_4_11__leaf_i_clk vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_5461_ core_0.execute.alu_mul_div.div_cur\[12\] _1838_ _1816_ _1896_ _1897_ vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_112_613 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7741__I1 core_0.decode.i_imm_pass\[15\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_152_793 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4412_ _1017_ _0857_ _0959_ _1018_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_7200_ _1431_ _0709_ _1414_ _3388_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_8180_ _0356_ clknet_leaf_126_i_clk core_0.execute.alu_mul_div.mul_res\[6\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_2_855 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5392_ _1233_ _1836_ _1837_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XPHY_EDGE_ROW_244_Right_244 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_112_657 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_239_842 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_EDGE_ROW_99_Right_99 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_112_679 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4343_ _0947_ _0958_ _0960_ _0961_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_2
Xclkbuf_leaf_68_i_clk clknet_4_15__leaf_i_clk clknet_leaf_68_i_clk vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_7131_ _3336_ _3331_ _3337_ _3338_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_0_111_178 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7062_ _1909_ _1585_ _3274_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_4274_ core_0.fetch.prev_request_pc\[10\] _0892_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_0_226_547 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6013_ _2271_ _2342_ _2354_ _2402_ _2403_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or4_1
XFILLER_0_241_506 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4357__C _0830_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6209__A1 _1600_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_213_208 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_207_761 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_207_772 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_241_539 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_2_537 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_27_81 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_234_591 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_222_753 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_19_Left_266 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
X_7964_ _0014_ clknet_leaf_28_i_clk net107 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_38_967 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6915_ net89 _3135_ _3139_ _3143_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_77_644 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_31_i_clk_I clknet_4_10__leaf_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_77_655 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7709__A1 _1085_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_159_2417 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_7895_ _0086_ clknet_leaf_72_i_clk core_0.decode.i_imm_pass\[4\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_147_510 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_178_189 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6144__I _2268_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_187_690 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_119_212 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6846_ core_0.execute.rf.reg_outputs\[2\]\[13\] _3092_ _3098_ _3103_ vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_77_699 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_119_245 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7684__B _1094_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_64_349 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_147_576 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_221 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6777_ core_0.ew_reg_ie\[3\] _2934_ _3063_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_2
X_3989_ _0616_ _0594_ _0617_ _0618_ _0619_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai211_4
XANTENNA__6932__A2 _1451_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_162_524 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4943__A1 _1400_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5728_ _2123_ _2125_ _2128_ _2129_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__5916__C _1624_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4599__I _1164_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6145__B1 _2264_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_28_Left_275 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_72_393 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5659_ _2058_ _2059_ _2060_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XTAP_TAPCELL_ROW_211_3050 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5499__A2 _1931_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_4_170 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_192 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_211_Right_211 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_103_668 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_4_1__f_i_clk_I clknet_3_0_0_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7329_ core_0.dec_sreg_store _2265_ _3502_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_0_217_525 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_183_2713 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_99_202 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5671__A2 _1529_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_37_Left_284 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_169_123 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5959__B1 _2260_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6620__A1 net32 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5423__A2 _1814_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_158_819 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_157_318 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_184_104 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_169_189 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_200_469 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_103_1748 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_56_839 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_138_543 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7176__A2 _1809_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_83_625 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_194_2842 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_83_636 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_95_496 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5187__A1 _0776_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_193_671 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_165_362 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_180_321 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_181_844 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_46_Left_293 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_36_563 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_319 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_130_18 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_180_332 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_91_691 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xrebuffer6 _0519_ net228 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_51_533 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_63_393 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_2_107 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_58_1205 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_140_218 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_180_387 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_2_118 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6687__A1 core_0.execute.rf.reg_outputs\[6\]\[9\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8235__CLK clknet_leaf_43_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_23_279 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_239_138 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_121_487 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6439__A1 _1059_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_114_1877 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_225_3208 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6439__B2 _2815_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_235_311 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_235_344 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_143_2229 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_207_2996 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_69_1345 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_78_419 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_204_786 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_188_454 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_59_622 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6611__A1 _2936_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5414__A2 _1758_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_82_1501 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_176_616 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_231_594 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4961_ _1301_ _1416_ _0115_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_35_937 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_147_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_19_508 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6700_ core_0.execute.rf.reg_outputs\[6\]\[15\] _2998_ _3016_ _3019_ vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3912_ _0547_ _0548_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_86_463 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7680_ _1113_ _1116_ _3780_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_47_839 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4892_ _1280_ core_0.fetch.out_buffer_data_pred _1359_ _1360_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_236_3348 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_58_187 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_156_340 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_175_159 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6631_ net27 _1148_ _2974_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_190_107 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_46_349 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5178__B2 core_0.execute.rf.reg_outputs\[6\]\[5\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_73_135 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_72 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6914__A2 _3129_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_156_384 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_27_552 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_15_694 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_rebuffer3_I _1641_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_144_535 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_156_395 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4925__A1 _0810_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6562_ core_0.dec_rf_ie\[1\] core_0.ew_reg_ie\[1\] _1985_ _2922_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_171_332 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_6_457 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_89_32 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_154_2358 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_42_522 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_89_43 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8301_ _0477_ clknet_leaf_12_i_clk net186 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_4
X_5513_ _0754_ _0756_ _1172_ _1945_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_0_171_376 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6493_ _2576_ _2870_ _2871_ _0192_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__6678__A1 _2961_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_112_421 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8232_ _0408_ clknet_leaf_43_i_clk core_0.execute.sreg_irq_pc.o_d\[4\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5444_ _1233_ _1872_ _1882_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_140_741 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_93_1630 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_112_454 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6848__B _3098_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_2_663 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_100_605 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_2_685 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4153__A2 _0769_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_8163_ _0339_ clknet_leaf_89_i_clk net100 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_4
XFILLER_0_1_162 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5375_ _1375_ _1818_ _1821_ _1822_ _1823_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_112_487 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5244__S _1460_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7114_ _1227_ _1501_ _3321_ _3322_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA__5471__C _1822_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4326_ _0725_ net49 _0943_ _0944_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_238_171 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8094_ _0270_ clknet_leaf_109_i_clk core_0.execute.rf.reg_outputs\[4\]\[1\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5102__A1 _1467_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7045_ _2587_ _3250_ _3258_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_4257_ core_0.fetch.dbg_out _0876_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__5043__I _1446_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_242_815 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_199_719 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5653__A2 _2053_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7679__B _1078_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_165_2487 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_241_325 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4700__I1 net67 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4188_ _0805_ net20 _0806_ _0807_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_4
XTAP_TAPCELL_ROW_165_2498 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_207_580 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_241_347 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_241_358 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_97_728 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_222_550 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6602__A1 _2929_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_210_734 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_96_249 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7947_ _0125_ clknet_leaf_5_i_clk core_0.execute.alu_mul_div.div_cur\[3\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_210_745 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_166_115 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_210_756 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_210_778 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_49_165 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_194_457 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_38_839 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_37_316 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7878_ _0069_ clknet_leaf_47_i_clk core_0.decode.i_instr_l\[3\] vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_4
XFILLER_0_77_496 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5169__A1 _0776_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_42_1017 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_6829_ core_0.execute.rf.reg_outputs\[2\]\[5\] _3092_ _3083_ _3094_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_65_658 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6905__A2 _3129_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_135_524 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_161_80 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_162_310 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8258__CLK clknet_leaf_36_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_64_179 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_190_652 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_45_360 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_33_500 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_61_842 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_162_365 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_116_771 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_122_207 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_150_527 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_162_387 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_103_410 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6758__B _3045_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5341__A1 _1508_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4144__A2 _0520_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5192__I1 net202 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_218_823 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5381__C _1822_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_53_1146 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_245_642 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_217_344 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_233_815 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5644__A2 _2034_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6841__A1 _2986_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4447__A3 _1041_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_129_2062 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_233_837 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_232_314 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_205_528 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_189_218 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5888__I core_0.execute.alu_mul_div.i_mul vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3910__B _0520_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_125_18 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_220_3149 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_87_216 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7397__A2 _3542_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_158_605 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_201_734 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_185_413 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_200_233 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_68_452 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_205_62 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3958__A2 _0578_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4080__A1 _0567_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7149__A2 _3177_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6940__C _1230_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_83_411 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_96_794 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_422 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_95_282 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XPHY_EDGE_ROW_54_Left_301 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__5837__B _2231_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_64_1275 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_172_107 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_64_1286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_126_513 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_50_37 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_126_524 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_138_384 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_126_535 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_138_395 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_126_557 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_12_653 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_24_522 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_114_719 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_221_72 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_36_382 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4383__A2 _0947_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_40_995 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_116_1906 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_12_706 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_180_184 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_231_3289 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_12_728 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_59_24 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_11_216 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_121_251 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4135__A2 _0753_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7343__I net202 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6387__C _2626_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5160_ core_0.execute.rf.reg_outputs\[1\]\[6\] _1608_ _1434_ core_0.execute.rf.reg_outputs\[6\]\[6\]
+ _1609_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XPHY_EDGE_ROW_63_Left_310 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__5883__A2 _0720_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_209_834 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7085__A1 _1909_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4111_ core_0.execute.prev_sys _0730_ _0731_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_0_75_34 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5091_ net93 _1492_ _1535_ _1539_ _1540_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai22_2
XFILLER_0_236_664 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_75_56 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4042_ core_0.execute.rf.reg_outputs\[7\]\[5\] _0529_ _0668_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6832__A1 _2972_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7499__B _3516_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_223_336 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_223_369 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_91_33 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_188_251 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7801_ _3796_ _3864_ _3865_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_78_249 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5399__A1 core_0.execute.alu_mul_div.div_cur\[5\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_430 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_182_68 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_441 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5993_ _2380_ _2383_ _2384_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_176_413 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_188_284 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_87_761 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7719__S _1946_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6060__A2 _2249_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3949__A2 _0542_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_87_772 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7732_ _3817_ _0485_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_19_305 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_176_457 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4944_ core_0.execute.sreg_priv_control.o_d\[4\] _1394_ _1404_ _1391_ _1405_ vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_164_608 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_327 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_59_496 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_176_479 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_163_107 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7663_ core_0.dec_sys _3766_ _1074_ _3767_ _3768_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_4875_ _0823_ _1321_ _1351_ _0094_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_46_157 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6899__A1 net97 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6614_ _2929_ _2958_ _2959_ _2960_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_0_46_168 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5466__C _1809_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_117_557 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7594_ _3675_ _3711_ _3712_ _3672_ _3713_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_7_766 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_61_116 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7560__A2 core_0.execute.pc_high_out\[0\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_160_803 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_579 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_842 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_131_72 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5571__A1 _1980_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6545_ _2913_ _0202_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_144_387 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_42_352 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_42_363 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7681__C _1046_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6476_ core_0.execute.alu_mul_div.mul_res\[14\] _2855_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__inv_2
XFILLER_0_71_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_112_240 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8215_ _0391_ clknet_leaf_36_i_clk net87 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_2
X_5427_ _1782_ _1784_ _1757_ _1867_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_100_435 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_772 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_167_2516 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_8146_ _0322_ clknet_leaf_115_i_clk core_0.execute.rf.reg_outputs\[1\]\[5\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_100_457 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5358_ core_0.execute.alu_mul_div.div_cur\[14\] _1713_ _1806_ vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA_input43_I i_req_data[14] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3885__A1 _0517_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_10_282 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7076__A1 core_0.execute.alu_mul_div.mul_res\[9\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
X_4309_ _0925_ _0887_ _0893_ _0926_ _0927_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_8077_ _0253_ clknet_leaf_92_i_clk core_0.execute.rf.reg_outputs\[5\]\[0\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_242_601 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5702__S _2102_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5289_ _1193_ _1738_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__inv_1
XANTENNA__6823__A1 _2951_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7028_ _1371_ core_0.execute.alu_mul_div.mul_res\[6\] _1939_ _3242_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_242_645 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_230_807 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_241_144 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4318__S _0725_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_97_558 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_194_210 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_178_2645 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_242_49 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_194_243 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4062__A1 _0567_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_139_148 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_194_254 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_65_422 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_77_282 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_100_1707 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_210_597 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_100_1718 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_154_107 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_182_416 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_194_287 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_191_2801 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_108_524 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_182_449 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_477 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_136_855 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_92_274 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_18_382 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5562__A1 _0964_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_162_162 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_33_352 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_151_858 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_150_357 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_150_368 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_clkbuf_leaf_0_i_clk_I clknet_4_0__leaf_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4117__A2 _0735_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5314__A1 core_0.execute.alu_mul_div.div_cur\[6\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_104_796 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_189_2785 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5865__A2 _1196_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_111_1847 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7067__A1 _1372_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_218_664 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_206_804 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6814__A1 _2996_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_232_111 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_232_155 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_232_177 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_204_2955 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_66_1304 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_216_72 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_204_2966 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_198_571 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_17_712 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_186_733 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_772 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_75_208 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4053__A1 net98 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_158_457 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_28_102 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_271 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7790__A2 _1134_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_61_58 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_122_1976 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_78_i_clk_I clknet_4_13__leaf_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_185_276 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_69 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_139_671 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_230 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_233_3307 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_84_775 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_84_786 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_166_490 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_232_82 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_28_179 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4660_ _1217_ _1214_ _1218_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_71_436 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_842 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_71_458 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_114_527 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_126_387 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4600__I0 core_0.ew_data\[6\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4591_ _1160_ net154 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_24_341 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_151_2328 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_153_184 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_24_352 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6330_ _1088_ _2711_ _2712_ _2332_ _2713_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai211_4
XFILLER_0_141_346 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_77_1433 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_51_182 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4697__I _1236_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_3_279 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6261_ _2626_ _2627_ _2645_ _2646_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_0_12_569 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_110_733 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8000_ _0177_ clknet_leaf_18_i_clk core_0.ew_submit vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_2
X_5212_ _0771_ core_0.execute.rf.reg_outputs\[4\]\[3\] _0778_ _1661_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_6192_ core_0.execute.pc_high_out\[7\] _2257_ _2577_ core_0.execute.sreg_irq_pc.o_d\[7\]
+ _2578_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_20_580 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_244_3436 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_208_130 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5143_ _1591_ _1592_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_209_664 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_209_675 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_224_612 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6805__A1 _2988_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_208_174 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5074_ _1467_ net183 _1523_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_236_494 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_223_133 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_224_667 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4025_ _0649_ _0594_ _0650_ _0651_ _0652_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai211_4
XTAP_TAPCELL_ROW_162_2457 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_223_155 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4292__A1 core_0.fetch.prev_request_pc\[3\] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_211_317 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_196_519 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_88_1573 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_79_569 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_220_862 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4044__A1 net99 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5976_ _1121_ _2007_ _2367_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_75_720 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_47_422 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_59_282 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_118_800 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7781__A2 _1133_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7715_ core_0.decode.i_imm_pass\[2\] _1064_ _3809_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_136_107 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_4927_ _1390_ _1391_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_192_758 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_90_701 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_263 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_118_855 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7646_ net115 _3729_ _3755_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_74_274 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_191_257 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7940__CLK clknet_leaf_43_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4858_ _0906_ _1306_ _1342_ _0086_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_90_745 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7533__A2 net18 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7577_ core_0.execute.pc_high_buff_out\[3\] _3682_ _3697_ _3698_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_27_190 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_62_469 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_144_173 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4789_ core_0.fetch.prev_request_pc\[12\] net225 _0880_ net164 _1299_ vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_0_160_633 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_173_2586 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_15_352 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_133_858 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6528_ _1729_ _2190_ _2904_ _0194_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_42_160 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_396 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7297__A1 _2825_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6459_ _2576_ _2837_ _2838_ _0191_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_30_355 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_189_Right_189 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__4400__I net83 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_2_290 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_399 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_208_3011 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_11_591 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8129_ _0305_ clknet_leaf_112_i_clk core_0.execute.rf.reg_outputs\[2\]\[4\] vccd1
+ vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_50_1116 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_227_494 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_126_2021 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_202_317 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_230_659 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6771__B _3057_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_168_722 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_506 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7221__A1 _1414_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_211_862 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_195_530 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_195_541 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7221__B2 _1431_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_97_399 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_48_1089 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7772__A2 _3766_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_219_3140 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_210_383 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4586__A2 net157 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_195_596 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5783__A1 _1711_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_155_438 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_65_252 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_155_449 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_26_617 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_61_1245 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_65_274 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_81_734 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_680 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_354 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7524__A2 _3641_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_182_279 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_191_780 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_137_2161 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_163_471 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_22_781 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_108_387 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7094__S _3189_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_801 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_123_335 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4889__A3 net20 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_119 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_34_683 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_156_Right_156 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_238_737 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5838__A2 _2231_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_72_1374 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_56_58 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_206_634 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_148_2290 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7460__A1 _0580_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_233_486 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_178_519 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_205_199 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6681__B _3004_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_202_851 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_48_208 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7212__A1 _1172_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6015__A2 _2400_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5830_ _1626_ _2225_ _2226_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_88_399 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_69_591 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_159_799 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_56_230 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5761_ _2036_ _2040_ _2162_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5774__A1 _2168_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_227_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7500_ _0709_ _3640_ _3643_ _0427_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_4712_ core_0.fetch.out_buffer_data_instr\[12\] _1255_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_173_246 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5692_ _1714_ _1592_ _2093_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_56_285 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_72_734 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7515__A2 _3646_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_112_41 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6949__S1 _1364_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7431_ core_0.execute.sreg_irq_pc.o_d\[8\] _3543_ _3589_ _3590_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_115_836 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_127_696 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4643_ _1196_ _1198_ _1201_ _1202_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_0_21_72 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_72_789 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_31_108 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_115_858 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7362_ _1724_ _2328_ _3531_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_97_10 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4574_ core_0.ew_data\[1\] net157 _1152_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_188_34 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_25_694 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7279__A1 _2716_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6313_ _2058_ _2695_ _1457_ _2696_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_130_839 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_40_653 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7293_ _1430_ _1422_ _3470_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_97_76 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5829__A2 _1615_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_697 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_0_750 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6244_ _2628_ _2042_ _2629_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_2
XPHY_EDGE_ROW_123_Right_123 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_228_247 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_244_707 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6348__S _2123_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4501__A2 _1091_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_244_729 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6175_ _1480_ _2559_ _2561_ _1684_ _2562_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_4
X_5126_ _1572_ _1573_ _1574_ _1575_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_0_224_420 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6254__A2 _1455_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6147__I _2260_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_197_806 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5057_ _0619_ _0624_ _0625_ _1460_ _1506_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai31_2
XFILLER_0_137_93 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4008_ _0630_ _0635_ _0636_ _0637_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_0_196_327 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7203__A1 _1430_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6006__A2 _1385_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4017__A1 _0567_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_0_498 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_137_405 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_220_692 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_153_92 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_175_2615 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_94_369 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_137_438 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5959_ core_0.execute.sreg_scratch.o_d\[2\] _2254_ _2260_ net9 _2350_ vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_35_403 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_165_769 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_118_641 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7506__A2 _3646_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_164_268 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_164_279 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_180_728 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5935__B _2326_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_7629_ _3732_ _3741_ _3742_ _0457_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA_output197_I net197 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_62_255 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_661 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_214_3081 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_22_119 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_90_597 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_160_463 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_133_699 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_31_664 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_686 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_174 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_132_2091 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_219_225 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_26_i_clk_I clknet_4_10__leaf_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output74_I net74 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_219_247 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_186_2744 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7690__A1 _1084_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_199_121 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_215_453 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7442__A1 _0615_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4256__A1 _0726_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_188_828 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_187_316 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_86_804 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_4_9__f_i_clk clknet_3_4_0_i_clk clknet_4_9__leaf_i_clk vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_TAPCELL_ROW_201_2925 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_27_840 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_97_163 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4008__A1 _0630_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_106_1779 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_97_196 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_195_360 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_197_2873 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_38_241 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_66_572 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_225_Right_225 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_38_285 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_143_408 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_745 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5508__A1 _1223_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6556__I0 net120 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_14_609 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_255 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7616__I _3731_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_123_110 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_163_290 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_299 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_22_631 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_112_839 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_74_1403 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6308__I0 _0626_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4731__A2 _1238_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_111_349 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4290_ core_0.fetch.prev_request_pc\[4\] _0906_ _0907_ core_0.fetch.prev_request_pc\[5\]
+ _0908_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_158_37 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_21_185 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6484__A2 _2531_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7681__A1 _1066_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_241_3406 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_225_228 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_219_792 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_206_420 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_177_2 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_83_34 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7980_ _0157_ clknet_leaf_43_i_clk core_0.execute.mem_stage_pc\[15\] vccd1 vccd1
+ vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_233_261 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5800__S _2190_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_83_67 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6931_ core_0.execute.alu_mul_div.mul_res\[0\] _3152_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_233_294 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4798__A2 _1241_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_16_61 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_85_1532 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_49_506 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_76_314 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6862_ core_0.execute.rf.reg_outputs\[1\]\[3\] _3108_ _3112_ _3113_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_88_174 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_221_489 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_92_807 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5813_ _2195_ _2203_ _2207_ _2211_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_0_174_511 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_239_3379 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_8_102 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6793_ _2967_ _3064_ _3073_ _0290_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_147_758 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7727__S _1946_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4014__A4 core_0.execute.rf.reg_outputs\[6\]\[7\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5211__A3 _0776_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5744_ _2000_ _2145_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_174_577 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_146_279 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_155_780 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5675_ _2074_ _2075_ _2076_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_161_238 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4970__A2 _1393_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_44_266 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_842 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_115_644 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_199_66 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7414_ _3543_ _3574_ _3575_ _0409_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__6172__A1 _1559_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_4626_ _1173_ _1179_ _1180_ _1181_ _1184_ _1185_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XTAP_TAPCELL_ROW_170_2556 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_96_1661 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_7345_ _0722_ _3516_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_40_450 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_13_664 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4557_ _1065_ _1043_ _1139_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_4
XANTENNA__4722__A2 _1253_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_130_647 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7276_ _3453_ _3454_ _3455_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_40_494 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4488_ _1037_ _1080_ _1081_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_12_196 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5490__B _1651_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_217_718 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6227_ _2242_ net216 _2613_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__7672__A1 _1431_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_0_580 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4486__A1 _1078_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6158_ _2099_ _2106_ _2123_ _2545_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_5_568 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6227__A2 net216 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7424__A1 _0648_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_5109_ _1556_ _1557_ _1558_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_4
XANTENNA__4238__A1 _0824_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_6089_ core_0.execute.alu_mul_div.i_mul core_0.execute.alu_mul_div.mul_res\[4\] _2478_
+ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_240_721 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_181_2685 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5986__A1 _2300_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4834__B _1170_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output112_I net112 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_67_336 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_184_319 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_193_842 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_45_1048 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_82_306 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_165_533 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_317 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_216_3110 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4005__A4 core_0.execute.rf.reg_outputs\[2\]\[8\] vccd1 vccd1 vssd1 vssd1
+ gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_94_177 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_137_246 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_520 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4410__A1 _1013_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_745 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_91_862 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_134_2120 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_145_290 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_63_597 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_383 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6163__A1 _2022_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_51_748 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_50_247 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_121_625 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5910__A1 _1531_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_121_636 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4713__A2 _1253_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_101_371 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput74 net74 dbg_pc[11] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XTAP_TAPCELL_ROW_56_1188 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_101_382 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7663__B2 _3767_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput85 net85 dbg_pc[7] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xoutput96 net96 dbg_r0[2] vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA__8014__CLK clknet_leaf_53_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4477__A1 _1066_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_108_1808 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_231_710 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_208_73 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_243_570 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_231_721 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_199_2902 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_188_636 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_231_754 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5977__A1 _1457_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8164__CLK clknet_leaf_88_i_clk vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_187_135 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_230_253 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_58_314 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_58_325 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_230_286 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7718__A2 _0514_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_175_319 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_74_807 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_168_371 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_46_509 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5729__A1 _1549_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_168_393 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_129_769 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_183_330 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_183_352 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_80_1473 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_143_227 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4952__A2 net216 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_119_1937 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_30_868 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_54_586 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5460_ _1822_ _1895_ _1896_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_2_801 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4411_ core_0.fetch.prev_request_pc\[3\] _0949_ _1017_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__5901__A1 net223 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_78_34 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_78_45 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5391_ _1763_ _1775_ _1836_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_7130_ _2855_ _1941_ _3337_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_4342_ _0827_ _0959_ _0960_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_78_89 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_10_667 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7061_ _3259_ _3269_ _3267_ _3273_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_4273_ _0889_ _0843_ _0844_ _0890_ _0891_ vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_0_10_678 vccd1 vccd1 vssd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6012_ _1378_ core_0.execute.sreg_irq_pc.o_d\[3\] _2401_ _2402_ vccd1 vccd1 vssd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
.ends

