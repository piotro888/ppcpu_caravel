VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO logo
  CLASS BLOCK ;
  FOREIGN logo ;
  ORIGIN 0.000 0.000 ;
  SIZE 740.000 BY 80.000 ;
  OBS
      LAYER Metal5 ;
        RECT -10.000 -10.000 750.000 90.000 ;
  END
END logo
END LIBRARY
